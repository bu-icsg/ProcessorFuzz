`define toAscii(x) { x / 8'ha + 8'h30, x % 8'ha + 8'h30 }

module RocketTile(
  input         cov_store,
  input         clock,
  input         reset,
  output        auto_broadcast_out_0_valid,
  output [39:0] auto_broadcast_out_0_iaddr,
  output [31:0] auto_broadcast_out_0_insn,
  output [2:0]  auto_broadcast_out_0_priv,
  output        auto_broadcast_out_0_exception,
  output        auto_broadcast_out_0_interrupt,
  output [63:0] auto_broadcast_out_0_cause,
  output [39:0] auto_broadcast_out_0_tval,
  output        auto_wfi_out_0,
  output        auto_cease_out_0,
  output        auto_halt_out_0,
  input         auto_int_in_xing_in_2_sync_0,
  input         auto_int_in_xing_in_1_sync_0,
  input         auto_int_in_xing_in_0_sync_0,
  input         auto_int_in_xing_in_0_sync_1,
  input         auto_intsink_in_sync_0,
  output        auto_trace_core_source_out_group_0_iretire,
  output [31:0] auto_trace_core_source_out_group_0_iaddr,
  output [3:0]  auto_trace_core_source_out_group_0_itype,
  output        auto_trace_core_source_out_group_0_ilastsize,
  output [3:0]  auto_trace_core_source_out_priv,
  output [31:0] auto_trace_core_source_out_tval,
  output [31:0] auto_trace_core_source_out_cause,
  input         auto_nmi_in_rnmi,
  input  [31:0] auto_nmi_in_rnmi_interrupt_vector,
  input  [31:0] auto_nmi_in_rnmi_exception_vector,
  input         auto_nmi_in_unmi,
  input  [31:0] auto_nmi_in_unmi_interrupt_vector,
  input  [31:0] auto_nmi_in_unmi_exception_vector,
  input  [31:0] auto_reset_vector_in,
  input         auto_hartid_in,
  input         auto_tl_master_xing_out_a_ready,
  output        auto_tl_master_xing_out_a_valid,
  output [2:0]  auto_tl_master_xing_out_a_bits_opcode,
  output [2:0]  auto_tl_master_xing_out_a_bits_param,
  output [3:0]  auto_tl_master_xing_out_a_bits_size,
  output [1:0]  auto_tl_master_xing_out_a_bits_source,
  output [31:0] auto_tl_master_xing_out_a_bits_address,
  output [7:0]  auto_tl_master_xing_out_a_bits_mask,
  output [63:0] auto_tl_master_xing_out_a_bits_data,
  output        auto_tl_master_xing_out_a_bits_corrupt,
  output        auto_tl_master_xing_out_b_ready,
  input         auto_tl_master_xing_out_b_valid,
  input  [2:0]  auto_tl_master_xing_out_b_bits_opcode,
  input  [1:0]  auto_tl_master_xing_out_b_bits_param,
  input  [3:0]  auto_tl_master_xing_out_b_bits_size,
  input  [1:0]  auto_tl_master_xing_out_b_bits_source,
  input  [31:0] auto_tl_master_xing_out_b_bits_address,
  input  [7:0]  auto_tl_master_xing_out_b_bits_mask,
  input  [63:0] auto_tl_master_xing_out_b_bits_data,
  input         auto_tl_master_xing_out_b_bits_corrupt,
  input         auto_tl_master_xing_out_c_ready,
  output        auto_tl_master_xing_out_c_valid,
  output [2:0]  auto_tl_master_xing_out_c_bits_opcode,
  output [2:0]  auto_tl_master_xing_out_c_bits_param,
  output [3:0]  auto_tl_master_xing_out_c_bits_size,
  output [1:0]  auto_tl_master_xing_out_c_bits_source,
  output [31:0] auto_tl_master_xing_out_c_bits_address,
  output [63:0] auto_tl_master_xing_out_c_bits_data,
  output        auto_tl_master_xing_out_c_bits_corrupt,
  output        auto_tl_master_xing_out_d_ready,
  input         auto_tl_master_xing_out_d_valid,
  input  [2:0]  auto_tl_master_xing_out_d_bits_opcode,
  input  [1:0]  auto_tl_master_xing_out_d_bits_param,
  input  [3:0]  auto_tl_master_xing_out_d_bits_size,
  input  [1:0]  auto_tl_master_xing_out_d_bits_source,
  input  [1:0]  auto_tl_master_xing_out_d_bits_sink,
  input         auto_tl_master_xing_out_d_bits_denied,
  input  [63:0] auto_tl_master_xing_out_d_bits_data,
  input         auto_tl_master_xing_out_d_bits_corrupt,
  input         auto_tl_master_xing_out_e_ready,
  output        auto_tl_master_xing_out_e_valid,
  output [1:0]  auto_tl_master_xing_out_e_bits_sink,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset,
  input         tlMasterXbar_halt,
  input         intXbar_halt,
  input         fpuOpt_halt,
  input         dcacheArb_halt,
  input         frontend_halt,
  input         dcache_halt,
  input         broadcast_3_halt,
  input         core_halt,
  input         broadcast_halt,
  input         broadcast_1_halt,
  input         ptw_halt,
  input         eos, // chath: added an end of simulation flag
  input         cov_sr,
  output reg    eos_hs, // eos handshake
  output reg [39:0] cmt_instr
);

  reg debug_print;
  string trace_dir;
  string test_dir;
  reg trace_en;
  integer fd;
  integer iteration;
  string iter;
  wire [63:0] mstatus_wire;

  initial begin
    test_dir = "/projectnb2/risc-v/chath/difuzzrtl/Fuzzer/17output/tests/";
    iteration = 0;
    if (!$value$plusargs("DEBUG=%d", debug_print)) begin
      debug_print = 0;
      //clock_count = 0;
    end
    if (!$value$plusargs("TRACE=%s", trace_dir)) begin
      trace_en = 0;
      trace_dir = "rtl_";
      fd = 0;
    end else begin 
      trace_en = 1;
      fd = 0; 
    end
  end


`ifndef SYNTHESIS
//integer x;
  always@(posedge eos) begin //chath: closing the file using the end of sim flag
    if (trace_en) begin
      if (fd!=32'd0) begin
	//for (int x = 0; x < 10 ; x++)begin
        $fflush(fd);
        $display("FLUSH CALLED");
 	$fclose(fd);
        eos_hs = 1'b1;
      end
    end
  end
  
  always@(negedge metaReset) begin
    if (trace_en) begin
      if (fd!=32'd0) begin
        $fflush(fd);
        $fclose(fd);
        $display("FLUSH CALLED");
      end
      eos_hs = 1'b0;
      iter.itoa(iteration);
      $display("TRACE enabled - %s", {trace_dir, "rtl_", iter,".log"});
      fd = $fopen({trace_dir, "rtl_", iter,".log"},"w");
      $fwrite(fd, "HartID mode PC INSTR WDATA COV\n");
      //sf = $fopen({test_dir,".input_0_",iter,".symbols_sub"}, "r");
      //init_queue(sf, sym_addrs_q);
      iteration = iteration + 1;
    end
  end

  assign mstatus_wire = {core.csr.io_status_sd, core.csr.io_status_zero2, core.csr.read_mstatus_hi_lo, core.csr.read_mstatus_lo};


  always @(posedge clock) begin
    cmt_instr = core.csr_io_trace_0_iaddr;
  end
  
  always @(posedge clock) begin
    if (trace_en) begin

      if (core.coreMonitorBundle_valid & ~core.reset) begin
        $fwrite(fd, "%d %d 0x%x ", core.io_hartid, core.csr_io_status_prv, core.csr_io_trace_0_iaddr);
        $fwrite(fd,"0x%x 0x%x", core.csr_io_trace_0_insn, core.coreMonitorBundle_wrenx ? core.rf_wdata : ( (core._GEN_262 || core.wb_ctrl_wfd) ? 64'hdeadbeef : 64'h0)); // @[core.scala 1258:17]
	$fwrite(fd," %x", mstatus_wire);
	$fwrite(fd," %x", core.csr.reg_mcause[7:0]);
	$fwrite(fd," %x", core.csr.reg_scause[7:0]);
	$fwrite(fd," %x", core.csr.reg_medeleg);
	$fwrite(fd," %x", core.csr.reg_mcounteren);
	$fwrite(fd," %x", core.csr.reg_scounteren);
	$fwrite(fd," %x", core.csr.reg_dcsr);
	$fwrite(fd," %d\n", io_covSum);
      end
      else if (core.csr_io_trace_0_exception) begin
        $fwrite(fd, "%d %d 0x%x ", core.io_hartid, core.csr_io_status_prv, core.csr_io_trace_0_iaddr);
        $fwrite(fd,"0x%x 0x%x", core.csr_io_trace_0_insn, core.coreMonitorBundle_wrenx ? core.rf_wdata : 64'h0);
	$fwrite(fd," %x", mstatus_wire);
	$fwrite(fd," %x", core.csr.reg_mcause[7:0]);
	$fwrite(fd," %x", core.csr.reg_scause[7:0]);
	$fwrite(fd," %x", core.csr.reg_medeleg);
	$fwrite(fd," %x", core.csr.reg_mcounteren);
	$fwrite(fd," %x", core.csr.reg_scounteren);
	$fwrite(fd," %x", core.csr.reg_dcsr);
	$fwrite(fd," %d EXCEPTION\n", io_covSum); 
      end
      if (core._T_159 & ~core.reset) begin
          $fwrite(fd, "DELAYED r%0d=%x\n",core.rf_waddr,core.rf_wdata);
      end
      if ( fpuOpt.frfWriteBundle_1_wrenf & ~core.reset ) begin
          $fwrite(fd, "DELAYED f%0d=%x %x\n",fpuOpt.waddr,fpuOpt._T_40, core.csr.reg_fflags);
      end
      if ( fpuOpt.load_wb & ~core.reset) begin
          $fwrite(fd, "DELAYED f%0d=%x %x\n",fpuOpt.load_wb_tag,fpuOpt.load_wb_data, core.csr.reg_fflags);
      end
    end
  end

`endif

`ifdef COV_SR
  integer i;
  //integer fd;
  reg cov_restore;
  integer c;
  reg [7:0] proc_num;
  reg [8*100:1] out;
  initial begin
    if ($value$plusargs("OUT=%s", out)) begin
      $display("Output directory: %0s\n", out);
    end
    if ($value$plusargs("COV_RESTORE=%b", cov_restore)) begin
      $display("Restoring coverage...");
    end
    proc_num = 8'd0;
    if (cov_restore) begin
      //$display("COV RESTORE");
      fd = $fopen({out, "/covmap/ptw.PTW_cov.dat"}, "r");
      if (fd == 0)
        $display("No saved %s, starting from zero", "ptw.PTW_cov");
      else begin
        for (i=0; i<1048576; i=i+1) begin
          c = $fgetc(fd);
          ptw.PTW_cov[i] = c[0];
        end
        $fclose(fd);
      end
      fd = $fopen({out, "/covmap/dcacheArb.HellaCacheArbiter_cov.dat"}, "r");
      if (fd == 0)
        $display("No saved %s, starting from zero", "dcacheArb.HellaCacheArbiter_cov");
      else begin
        for (i=0; i<2; i=i+1) begin
          c = $fgetc(fd);
          dcacheArb.HellaCacheArbiter_cov[i] = c[0];
        end
        $fclose(fd);
      end
      fd = $fopen({out, "/covmap/tlMasterXbar.TLXbar_7_cov.dat"}, "r");
      if (fd == 0)
        $display("No saved %s, starting from zero", "tlMasterXbar.TLXbar_7_cov");
      else begin
        for (i=0; i<8; i=i+1) begin
          c = $fgetc(fd);
          tlMasterXbar.TLXbar_7_cov[i] = c[0];
        end
        $fclose(fd);
      end
      fd = $fopen({out, "/covmap/dcache.DCache_cov.dat"}, "r");
      if (fd == 0)
        $display("No saved %s, starting from zero", "dcache.DCache_cov");
      else begin
        for (i=0; i<1048576; i=i+1) begin
          c = $fgetc(fd);
          dcache.DCache_cov[i] = c[0];
        end
        $fclose(fd);
      end
      fd = $fopen({out, "/covmap/dcache.pma_checker.TLB_cov.dat"}, "r");
      if (fd == 0)
        $display("No saved %s, starting from zero", "dcache.pma_checker.TLB_cov");
      else begin
        for (i=0; i<1048576; i=i+1) begin
          c = $fgetc(fd);
          dcache.pma_checker.TLB_cov[i] = c[0];
        end
        $fclose(fd);
      end
      fd = $fopen({out, "/covmap/dcache.tlb.TLB_cov.dat"}, "r");
      if (fd == 0)
        $display("No saved %s, starting from zero", "dcache.tlb.TLB_cov");
      else begin
        for (i=0; i<1048576; i=i+1) begin
          c = $fgetc(fd);
          dcache.tlb.TLB_cov[i] = c[0];
        end
        $fclose(fd);
      end
      fd = $fopen({out, "/covmap/core.Rocket_cov.dat"}, "r");
      if (fd == 0)
        $display("No saved %s, starting from zero", "core.Rocket_cov");
      else begin
        for (i=0; i<1048576; i=i+1) begin
          c = $fgetc(fd);
          core.Rocket_cov[i] = c[0];
        end
        $fclose(fd);
      end
      fd = $fopen({out, "/covmap/core.csr.CSRFile_cov.dat"}, "r");
      if (fd == 0)
        $display("No saved %s, starting from zero", "core.csr.CSRFile_cov");
      else begin
        for (i=0; i<1048576; i=i+1) begin
          c = $fgetc(fd);
          core.csr.CSRFile_cov[i] = c[0];
        end
        $fclose(fd);
      end
      fd = $fopen({out, "/covmap/core.div.MulDiv_cov.dat"}, "r");
      if (fd == 0)
        $display("No saved %s, starting from zero", "core.div.MulDiv_cov");
      else begin
        for (i=0; i<1048576; i=i+1) begin
          c = $fgetc(fd);
          core.div.MulDiv_cov[i] = c[0];
        end
        $fclose(fd);
      end
      fd = $fopen({out, "/covmap/core.ibuf.IBuf_cov.dat"}, "r");
      if (fd == 0)
        $display("No saved %s, starting from zero", "core.ibuf.IBuf_cov");
      else begin
        for (i=0; i<4; i=i+1) begin
          c = $fgetc(fd);
          core.ibuf.IBuf_cov[i] = c[0];
        end
        $fclose(fd);
      end
      fd = $fopen({out, "/covmap/fpuOpt.FPU_cov.dat"}, "r");
      if (fd == 0)
        $display("No saved %s, starting from zero", "fpuOpt.FPU_cov");
      else begin
        for (i=0; i<1048576; i=i+1) begin
          c = $fgetc(fd);
          fpuOpt.FPU_cov[i] = c[0];
        end
        $fclose(fd);
      end
      fd = $fopen({out, "/covmap/fpuOpt.divSqrt_1.divSqrtRecFNToRaw.divSqrtRawFN_.DivSqrtRawFN_small_1_cov.dat"}, "r");
      if (fd == 0)
        $display("No saved %s, starting from zero", "fpuOpt.divSqrt_1.divSqrtRecFNToRaw.divSqrtRawFN_.DivSqrtRawFN_small_1_cov");
      else begin
        for (i=0; i<32; i=i+1) begin
          c = $fgetc(fd);
          fpuOpt.divSqrt_1.divSqrtRecFNToRaw.divSqrtRawFN_.DivSqrtRawFN_small_1_cov[i] = c[0];
        end
        $fclose(fd);
      end
      fd = $fopen({out, "/covmap/fpuOpt.ifpu.IntToFP_cov.dat"}, "r");
      if (fd == 0)
        $display("No saved %s, starting from zero", "fpuOpt.ifpu.IntToFP_cov");
      else begin
        for (i=0; i<16; i=i+1) begin
          c = $fgetc(fd);
          fpuOpt.ifpu.IntToFP_cov[i] = c[0];
        end
        $fclose(fd);
      end
      fd = $fopen({out, "/covmap/fpuOpt.divSqrt.divSqrtRecFNToRaw.divSqrtRawFN_.DivSqrtRawFN_small_cov.dat"}, "r");
      if (fd == 0)
        $display("No saved %s, starting from zero", "fpuOpt.divSqrt.divSqrtRecFNToRaw.divSqrtRawFN_.DivSqrtRawFN_small_cov");
      else begin
        for (i=0; i<32; i=i+1) begin
          c = $fgetc(fd);
          fpuOpt.divSqrt.divSqrtRecFNToRaw.divSqrtRawFN_.DivSqrtRawFN_small_cov[i] = c[0];
        end
        $fclose(fd);
      end
      fd = $fopen({out, "/covmap/fpuOpt.fpmu.FPToFP_cov.dat"}, "r");
      if (fd == 0)
        $display("No saved %s, starting from zero", "fpuOpt.fpmu.FPToFP_cov");
      else begin
        for (i=0; i<64; i=i+1) begin
          c = $fgetc(fd);
          fpuOpt.fpmu.FPToFP_cov[i] = c[0];
        end
        $fclose(fd);
      end
      fd = $fopen({out, "/covmap/fpuOpt.dfma.fma.MulAddRecFNPipe_1_cov.dat"}, "r");
      if (fd == 0)
        $display("No saved %s, starting from zero", "fpuOpt.dfma.fma.MulAddRecFNPipe_1_cov");
      else begin
        for (i=0; i<2; i=i+1) begin
          c = $fgetc(fd);
          fpuOpt.dfma.fma.MulAddRecFNPipe_1_cov[i] = c[0];
        end
        $fclose(fd);
      end
      fd = $fopen({out, "/covmap/fpuOpt.fpiu.FPToInt_cov.dat"}, "r");
      if (fd == 0)
        $display("No saved %s, starting from zero", "fpuOpt.fpiu.FPToInt_cov");
      else begin
        for (i=0; i<16; i=i+1) begin
          c = $fgetc(fd);
          fpuOpt.fpiu.FPToInt_cov[i] = c[0];
        end
        $fclose(fd);
      end
      fd = $fopen({out, "/covmap/fpuOpt.sfma.fma.MulAddRecFNPipe_cov.dat"}, "r");
      if (fd == 0)
        $display("No saved %s, starting from zero", "fpuOpt.sfma.fma.MulAddRecFNPipe_cov");
      else begin
        for (i=0; i<2; i=i+1) begin
          c = $fgetc(fd);
          fpuOpt.sfma.fma.MulAddRecFNPipe_cov[i] = c[0];
        end
        $fclose(fd);
      end
      fd = $fopen({out, "/covmap/frontend.Frontend_cov.dat"}, "r");
      if (fd == 0)
        $display("No saved %s, starting from zero", "frontend.Frontend_cov");
      else begin
        for (i=0; i<64; i=i+1) begin
          c = $fgetc(fd);
          frontend.Frontend_cov[i] = c[0];
        end
        $fclose(fd);
      end
      fd = $fopen({out, "/covmap/frontend.icache.ICache_cov.dat"}, "r");
      if (fd == 0)
        $display("No saved %s, starting from zero", "frontend.icache.ICache_cov");
      else begin
        for (i=0; i<64; i=i+1) begin
          c = $fgetc(fd);
          frontend.icache.ICache_cov[i] = c[0];
        end
        $fclose(fd);
      end
      fd = $fopen({out, "/covmap/frontend.fq.ShiftQueue_cov.dat"}, "r");
      if (fd == 0)
        $display("No saved %s, starting from zero", "frontend.fq.ShiftQueue_cov");
      else begin
        for (i=0; i<2; i=i+1) begin
          c = $fgetc(fd);
          frontend.fq.ShiftQueue_cov[i] = c[0];
        end
        $fclose(fd);
      end
      fd = $fopen({out, "/covmap/frontend.tlb.TLB_1_cov.dat"}, "r");
      if (fd == 0)
        $display("No saved %s, starting from zero", "frontend.tlb.TLB_1_cov");
      else begin
        for (i=0; i<1048576; i=i+1) begin
          c = $fgetc(fd);
          frontend.tlb.TLB_1_cov[i] = c[0];
        end
        $fclose(fd);
      end
      fd = $fopen({out, "/covmap/frontend.btb.BTB_cov.dat"}, "r");
      if (fd == 0)
        $display("No saved %s, starting from zero", "frontend.btb.BTB_cov");
      else begin
        for (i=0; i<1048576; i=i+1) begin
          c = $fgetc(fd);
          frontend.btb.BTB_cov[i] = c[0];
        end
        $fclose(fd);
      end
    end

  end

  always @(posedge cov_sr) begin
    if (cov_store) begin
      fd = $fopen({out, "/covmap/ptw.PTW_cov.dat"}, "w");
      for (i=0; i<1048576; i=i+1)
        $fwrite(fd, "%0b", ptw.PTW_cov[i]);
      $fclose(fd);
      fd = $fopen({out, "/covmap/dcacheArb.HellaCacheArbiter_cov.dat"}, "w");
      for (i=0; i<2; i=i+1)
        $fwrite(fd, "%0b", dcacheArb.HellaCacheArbiter_cov[i]);
      $fclose(fd);
      fd = $fopen({out, "/covmap/tlMasterXbar.TLXbar_7_cov.dat"}, "w");
      for (i=0; i<8; i=i+1)
        $fwrite(fd, "%0b", tlMasterXbar.TLXbar_7_cov[i]);
      $fclose(fd);
      fd = $fopen({out, "/covmap/dcache.DCache_cov.dat"}, "w");
      for (i=0; i<1048576; i=i+1)
        $fwrite(fd, "%0b", dcache.DCache_cov[i]);
      $fclose(fd);
      fd = $fopen({out, "/covmap/dcache.pma_checker.TLB_cov.dat"}, "w");
      for (i=0; i<1048576; i=i+1)
        $fwrite(fd, "%0b", dcache.pma_checker.TLB_cov[i]);
      $fclose(fd);
      fd = $fopen({out, "/covmap/dcache.tlb.TLB_cov.dat"}, "w");
      for (i=0; i<1048576; i=i+1)
        $fwrite(fd, "%0b", dcache.tlb.TLB_cov[i]);
      $fclose(fd);
      fd = $fopen({out, "/covmap/core.Rocket_cov.dat"}, "w");
      for (i=0; i<1048576; i=i+1)
        $fwrite(fd, "%0b", core.Rocket_cov[i]);
      $fclose(fd);
      fd = $fopen({out, "/covmap/core.csr.CSRFile_cov.dat"}, "w");
      for (i=0; i<1048576; i=i+1)
        $fwrite(fd, "%0b", core.csr.CSRFile_cov[i]);
      $fclose(fd);
      fd = $fopen({out, "/covmap/core.div.MulDiv_cov.dat"}, "w");
      for (i=0; i<1048576; i=i+1)
        $fwrite(fd, "%0b", core.div.MulDiv_cov[i]);
      $fclose(fd);
      fd = $fopen({out, "/covmap/core.ibuf.IBuf_cov.dat"}, "w");
      for (i=0; i<4; i=i+1)
        $fwrite(fd, "%0b", core.ibuf.IBuf_cov[i]);
      $fclose(fd);
      fd = $fopen({out, "/covmap/fpuOpt.FPU_cov.dat"}, "w");
      for (i=0; i<1048576; i=i+1)
        $fwrite(fd, "%0b", fpuOpt.FPU_cov[i]);
      $fclose(fd);
      fd = $fopen({out, "/covmap/fpuOpt.divSqrt_1.divSqrtRecFNToRaw.divSqrtRawFN_.DivSqrtRawFN_small_1_cov.dat"}, "w");
      for (i=0; i<32; i=i+1)
        $fwrite(fd, "%0b", fpuOpt.divSqrt_1.divSqrtRecFNToRaw.divSqrtRawFN_.DivSqrtRawFN_small_1_cov[i]);
      $fclose(fd);
      fd = $fopen({out, "/covmap/fpuOpt.ifpu.IntToFP_cov.dat"}, "w");
      for (i=0; i<16; i=i+1)
        $fwrite(fd, "%0b", fpuOpt.ifpu.IntToFP_cov[i]);
      $fclose(fd);
      fd = $fopen({out, "/covmap/fpuOpt.divSqrt.divSqrtRecFNToRaw.divSqrtRawFN_.DivSqrtRawFN_small_cov.dat"}, "w");
      for (i=0; i<32; i=i+1)
        $fwrite(fd, "%0b", fpuOpt.divSqrt.divSqrtRecFNToRaw.divSqrtRawFN_.DivSqrtRawFN_small_cov[i]);
      $fclose(fd);
      fd = $fopen({out, "/covmap/fpuOpt.fpmu.FPToFP_cov.dat"}, "w");
      for (i=0; i<64; i=i+1)
        $fwrite(fd, "%0b", fpuOpt.fpmu.FPToFP_cov[i]);
      $fclose(fd);
      fd = $fopen({out, "/covmap/fpuOpt.dfma.fma.MulAddRecFNPipe_1_cov.dat"}, "w");
      for (i=0; i<2; i=i+1)
        $fwrite(fd, "%0b", fpuOpt.dfma.fma.MulAddRecFNPipe_1_cov[i]);
      $fclose(fd);
      fd = $fopen({out, "/covmap/fpuOpt.fpiu.FPToInt_cov.dat"}, "w");
      for (i=0; i<16; i=i+1)
        $fwrite(fd, "%0b", fpuOpt.fpiu.FPToInt_cov[i]);
      $fclose(fd);
      fd = $fopen({out, "/covmap/fpuOpt.sfma.fma.MulAddRecFNPipe_cov.dat"}, "w");
      for (i=0; i<2; i=i+1)
        $fwrite(fd, "%0b", fpuOpt.sfma.fma.MulAddRecFNPipe_cov[i]);
      $fclose(fd);
      fd = $fopen({out, "/covmap/frontend.Frontend_cov.dat"}, "w");
      for (i=0; i<64; i=i+1)
        $fwrite(fd, "%0b", frontend.Frontend_cov[i]);
      $fclose(fd);
      fd = $fopen({out, "/covmap/frontend.icache.ICache_cov.dat"}, "w");
      for (i=0; i<64; i=i+1)
        $fwrite(fd, "%0b", frontend.icache.ICache_cov[i]);
      $fclose(fd);
      fd = $fopen({out, "/covmap/frontend.fq.ShiftQueue_cov.dat"}, "w");
      for (i=0; i<2; i=i+1)
        $fwrite(fd, "%0b", frontend.fq.ShiftQueue_cov[i]);
      $fclose(fd);
      fd = $fopen({out, "/covmap/frontend.tlb.TLB_1_cov.dat"}, "w");
      for (i=0; i<1048576; i=i+1)
        $fwrite(fd, "%0b", frontend.tlb.TLB_1_cov[i]);
      $fclose(fd);
      fd = $fopen({out, "/covmap/frontend.btb.BTB_cov.dat"}, "w");
      for (i=0; i<1048576; i=i+1)
        $fwrite(fd, "%0b", frontend.btb.BTB_cov[i]);
      $fclose(fd);
    end
  end
`endif


  wire  tlMasterXbar_clock; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_reset; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_in_1_a_ready; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_in_1_a_valid; // @[BaseTile.scala 195:42]
  wire [31:0] tlMasterXbar_auto_in_1_a_bits_address; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_in_1_d_valid; // @[BaseTile.scala 195:42]
  wire [2:0] tlMasterXbar_auto_in_1_d_bits_opcode; // @[BaseTile.scala 195:42]
  wire [3:0] tlMasterXbar_auto_in_1_d_bits_size; // @[BaseTile.scala 195:42]
  wire [63:0] tlMasterXbar_auto_in_1_d_bits_data; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_in_1_d_bits_corrupt; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_in_0_a_ready; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_in_0_a_valid; // @[BaseTile.scala 195:42]
  wire [2:0] tlMasterXbar_auto_in_0_a_bits_opcode; // @[BaseTile.scala 195:42]
  wire [2:0] tlMasterXbar_auto_in_0_a_bits_param; // @[BaseTile.scala 195:42]
  wire [3:0] tlMasterXbar_auto_in_0_a_bits_size; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_in_0_a_bits_source; // @[BaseTile.scala 195:42]
  wire [31:0] tlMasterXbar_auto_in_0_a_bits_address; // @[BaseTile.scala 195:42]
  wire [7:0] tlMasterXbar_auto_in_0_a_bits_mask; // @[BaseTile.scala 195:42]
  wire [63:0] tlMasterXbar_auto_in_0_a_bits_data; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_in_0_b_ready; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_in_0_b_valid; // @[BaseTile.scala 195:42]
  wire [1:0] tlMasterXbar_auto_in_0_b_bits_param; // @[BaseTile.scala 195:42]
  wire [3:0] tlMasterXbar_auto_in_0_b_bits_size; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_in_0_b_bits_source; // @[BaseTile.scala 195:42]
  wire [31:0] tlMasterXbar_auto_in_0_b_bits_address; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_in_0_c_ready; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_in_0_c_valid; // @[BaseTile.scala 195:42]
  wire [2:0] tlMasterXbar_auto_in_0_c_bits_opcode; // @[BaseTile.scala 195:42]
  wire [2:0] tlMasterXbar_auto_in_0_c_bits_param; // @[BaseTile.scala 195:42]
  wire [3:0] tlMasterXbar_auto_in_0_c_bits_size; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_in_0_c_bits_source; // @[BaseTile.scala 195:42]
  wire [31:0] tlMasterXbar_auto_in_0_c_bits_address; // @[BaseTile.scala 195:42]
  wire [63:0] tlMasterXbar_auto_in_0_c_bits_data; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_in_0_d_ready; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_in_0_d_valid; // @[BaseTile.scala 195:42]
  wire [2:0] tlMasterXbar_auto_in_0_d_bits_opcode; // @[BaseTile.scala 195:42]
  wire [1:0] tlMasterXbar_auto_in_0_d_bits_param; // @[BaseTile.scala 195:42]
  wire [3:0] tlMasterXbar_auto_in_0_d_bits_size; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_in_0_d_bits_source; // @[BaseTile.scala 195:42]
  wire [1:0] tlMasterXbar_auto_in_0_d_bits_sink; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_in_0_d_bits_denied; // @[BaseTile.scala 195:42]
  wire [63:0] tlMasterXbar_auto_in_0_d_bits_data; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_in_0_e_ready; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_in_0_e_valid; // @[BaseTile.scala 195:42]
  wire [1:0] tlMasterXbar_auto_in_0_e_bits_sink; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_out_a_ready; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_out_a_valid; // @[BaseTile.scala 195:42]
  wire [2:0] tlMasterXbar_auto_out_a_bits_opcode; // @[BaseTile.scala 195:42]
  wire [2:0] tlMasterXbar_auto_out_a_bits_param; // @[BaseTile.scala 195:42]
  wire [3:0] tlMasterXbar_auto_out_a_bits_size; // @[BaseTile.scala 195:42]
  wire [1:0] tlMasterXbar_auto_out_a_bits_source; // @[BaseTile.scala 195:42]
  wire [31:0] tlMasterXbar_auto_out_a_bits_address; // @[BaseTile.scala 195:42]
  wire [7:0] tlMasterXbar_auto_out_a_bits_mask; // @[BaseTile.scala 195:42]
  wire [63:0] tlMasterXbar_auto_out_a_bits_data; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_out_b_ready; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_out_b_valid; // @[BaseTile.scala 195:42]
  wire [2:0] tlMasterXbar_auto_out_b_bits_opcode; // @[BaseTile.scala 195:42]
  wire [1:0] tlMasterXbar_auto_out_b_bits_param; // @[BaseTile.scala 195:42]
  wire [3:0] tlMasterXbar_auto_out_b_bits_size; // @[BaseTile.scala 195:42]
  wire [1:0] tlMasterXbar_auto_out_b_bits_source; // @[BaseTile.scala 195:42]
  wire [31:0] tlMasterXbar_auto_out_b_bits_address; // @[BaseTile.scala 195:42]
  wire [7:0] tlMasterXbar_auto_out_b_bits_mask; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_out_b_bits_corrupt; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_out_c_ready; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_out_c_valid; // @[BaseTile.scala 195:42]
  wire [2:0] tlMasterXbar_auto_out_c_bits_opcode; // @[BaseTile.scala 195:42]
  wire [2:0] tlMasterXbar_auto_out_c_bits_param; // @[BaseTile.scala 195:42]
  wire [3:0] tlMasterXbar_auto_out_c_bits_size; // @[BaseTile.scala 195:42]
  wire [1:0] tlMasterXbar_auto_out_c_bits_source; // @[BaseTile.scala 195:42]
  wire [31:0] tlMasterXbar_auto_out_c_bits_address; // @[BaseTile.scala 195:42]
  wire [63:0] tlMasterXbar_auto_out_c_bits_data; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_out_d_ready; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_out_d_valid; // @[BaseTile.scala 195:42]
  wire [2:0] tlMasterXbar_auto_out_d_bits_opcode; // @[BaseTile.scala 195:42]
  wire [1:0] tlMasterXbar_auto_out_d_bits_param; // @[BaseTile.scala 195:42]
  wire [3:0] tlMasterXbar_auto_out_d_bits_size; // @[BaseTile.scala 195:42]
  wire [1:0] tlMasterXbar_auto_out_d_bits_source; // @[BaseTile.scala 195:42]
  wire [1:0] tlMasterXbar_auto_out_d_bits_sink; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_out_d_bits_denied; // @[BaseTile.scala 195:42]
  wire [63:0] tlMasterXbar_auto_out_d_bits_data; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_out_d_bits_corrupt; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_out_e_ready; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_auto_out_e_valid; // @[BaseTile.scala 195:42]
  wire [1:0] tlMasterXbar_auto_out_e_bits_sink; // @[BaseTile.scala 195:42]
  wire [29:0] tlMasterXbar_io_covSum; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_metaAssert; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_metaReset; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_monitor_halt; // @[BaseTile.scala 195:42]
  wire  tlMasterXbar_monitor_1_halt; // @[BaseTile.scala 195:42]
  wire  intXbar_auto_int_in_3_0; // @[BaseTile.scala 197:37]
  wire  intXbar_auto_int_in_2_0; // @[BaseTile.scala 197:37]
  wire  intXbar_auto_int_in_1_0; // @[BaseTile.scala 197:37]
  wire  intXbar_auto_int_in_1_1; // @[BaseTile.scala 197:37]
  wire  intXbar_auto_int_in_0_0; // @[BaseTile.scala 197:37]
  wire  intXbar_auto_int_out_0; // @[BaseTile.scala 197:37]
  wire  intXbar_auto_int_out_1; // @[BaseTile.scala 197:37]
  wire  intXbar_auto_int_out_2; // @[BaseTile.scala 197:37]
  wire  intXbar_auto_int_out_3; // @[BaseTile.scala 197:37]
  wire  intXbar_auto_int_out_4; // @[BaseTile.scala 197:37]
  wire [29:0] intXbar_io_covSum; // @[BaseTile.scala 197:37]
  wire  intXbar_metaAssert; // @[BaseTile.scala 197:37]
  wire  broadcast_auto_in; // @[BundleBridge.scala 196:31]
  wire  broadcast_auto_out; // @[BundleBridge.scala 196:31]
  wire [29:0] broadcast_io_covSum; // @[BundleBridge.scala 196:31]
  wire  broadcast_metaAssert; // @[BundleBridge.scala 196:31]
  wire [31:0] broadcast_1_auto_in; // @[BundleBridge.scala 196:31]
  wire [31:0] broadcast_1_auto_out_1; // @[BundleBridge.scala 196:31]
  wire [29:0] broadcast_1_io_covSum; // @[BundleBridge.scala 196:31]
  wire  broadcast_1_metaAssert; // @[BundleBridge.scala 196:31]
  wire  broadcast_3_auto_in_0_valid; // @[BundleBridge.scala 196:31]
  wire [39:0] broadcast_3_auto_in_0_iaddr; // @[BundleBridge.scala 196:31]
  wire [31:0] broadcast_3_auto_in_0_insn; // @[BundleBridge.scala 196:31]
  wire [2:0] broadcast_3_auto_in_0_priv; // @[BundleBridge.scala 196:31]
  wire  broadcast_3_auto_in_0_exception; // @[BundleBridge.scala 196:31]
  wire  broadcast_3_auto_in_0_interrupt; // @[BundleBridge.scala 196:31]
  wire [63:0] broadcast_3_auto_in_0_cause; // @[BundleBridge.scala 196:31]
  wire [39:0] broadcast_3_auto_in_0_tval; // @[BundleBridge.scala 196:31]
  wire  broadcast_3_auto_out_0_valid; // @[BundleBridge.scala 196:31]
  wire [39:0] broadcast_3_auto_out_0_iaddr; // @[BundleBridge.scala 196:31]
  wire [31:0] broadcast_3_auto_out_0_insn; // @[BundleBridge.scala 196:31]
  wire [2:0] broadcast_3_auto_out_0_priv; // @[BundleBridge.scala 196:31]
  wire  broadcast_3_auto_out_0_exception; // @[BundleBridge.scala 196:31]
  wire  broadcast_3_auto_out_0_interrupt; // @[BundleBridge.scala 196:31]
  wire [63:0] broadcast_3_auto_out_0_cause; // @[BundleBridge.scala 196:31]
  wire [39:0] broadcast_3_auto_out_0_tval; // @[BundleBridge.scala 196:31]
  wire [29:0] broadcast_3_io_covSum; // @[BundleBridge.scala 196:31]
  wire  broadcast_3_metaAssert; // @[BundleBridge.scala 196:31]
  wire  dcache_gated_clock; // @[HellaCache.scala 265:43]
  wire  dcache_reset; // @[HellaCache.scala 265:43]
  wire  dcache_auto_out_a_ready; // @[HellaCache.scala 265:43]
  wire  dcache_auto_out_a_valid; // @[HellaCache.scala 265:43]
  wire [2:0] dcache_auto_out_a_bits_opcode; // @[HellaCache.scala 265:43]
  wire [2:0] dcache_auto_out_a_bits_param; // @[HellaCache.scala 265:43]
  wire [3:0] dcache_auto_out_a_bits_size; // @[HellaCache.scala 265:43]
  wire  dcache_auto_out_a_bits_source; // @[HellaCache.scala 265:43]
  wire [31:0] dcache_auto_out_a_bits_address; // @[HellaCache.scala 265:43]
  wire [7:0] dcache_auto_out_a_bits_mask; // @[HellaCache.scala 265:43]
  wire [63:0] dcache_auto_out_a_bits_data; // @[HellaCache.scala 265:43]
  wire  dcache_auto_out_b_ready; // @[HellaCache.scala 265:43]
  wire  dcache_auto_out_b_valid; // @[HellaCache.scala 265:43]
  wire [1:0] dcache_auto_out_b_bits_param; // @[HellaCache.scala 265:43]
  wire [3:0] dcache_auto_out_b_bits_size; // @[HellaCache.scala 265:43]
  wire  dcache_auto_out_b_bits_source; // @[HellaCache.scala 265:43]
  wire [31:0] dcache_auto_out_b_bits_address; // @[HellaCache.scala 265:43]
  wire  dcache_auto_out_c_ready; // @[HellaCache.scala 265:43]
  wire  dcache_auto_out_c_valid; // @[HellaCache.scala 265:43]
  wire [2:0] dcache_auto_out_c_bits_opcode; // @[HellaCache.scala 265:43]
  wire [2:0] dcache_auto_out_c_bits_param; // @[HellaCache.scala 265:43]
  wire [3:0] dcache_auto_out_c_bits_size; // @[HellaCache.scala 265:43]
  wire  dcache_auto_out_c_bits_source; // @[HellaCache.scala 265:43]
  wire [31:0] dcache_auto_out_c_bits_address; // @[HellaCache.scala 265:43]
  wire [63:0] dcache_auto_out_c_bits_data; // @[HellaCache.scala 265:43]
  wire  dcache_auto_out_d_ready; // @[HellaCache.scala 265:43]
  wire  dcache_auto_out_d_valid; // @[HellaCache.scala 265:43]
  wire [2:0] dcache_auto_out_d_bits_opcode; // @[HellaCache.scala 265:43]
  wire [1:0] dcache_auto_out_d_bits_param; // @[HellaCache.scala 265:43]
  wire [3:0] dcache_auto_out_d_bits_size; // @[HellaCache.scala 265:43]
  wire  dcache_auto_out_d_bits_source; // @[HellaCache.scala 265:43]
  wire [1:0] dcache_auto_out_d_bits_sink; // @[HellaCache.scala 265:43]
  wire  dcache_auto_out_d_bits_denied; // @[HellaCache.scala 265:43]
  wire [63:0] dcache_auto_out_d_bits_data; // @[HellaCache.scala 265:43]
  wire  dcache_auto_out_e_ready; // @[HellaCache.scala 265:43]
  wire  dcache_auto_out_e_valid; // @[HellaCache.scala 265:43]
  wire [1:0] dcache_auto_out_e_bits_sink; // @[HellaCache.scala 265:43]
  wire  dcache_io_cpu_req_ready; // @[HellaCache.scala 265:43]
  wire  dcache_io_cpu_req_valid; // @[HellaCache.scala 265:43]
  wire [39:0] dcache_io_cpu_req_bits_addr; // @[HellaCache.scala 265:43]
  wire [6:0] dcache_io_cpu_req_bits_tag; // @[HellaCache.scala 265:43]
  wire [4:0] dcache_io_cpu_req_bits_cmd; // @[HellaCache.scala 265:43]
  wire [1:0] dcache_io_cpu_req_bits_size; // @[HellaCache.scala 265:43]
  wire  dcache_io_cpu_req_bits_signed; // @[HellaCache.scala 265:43]
  wire  dcache_io_cpu_req_bits_phys; // @[HellaCache.scala 265:43]
  wire  dcache_io_cpu_s1_kill; // @[HellaCache.scala 265:43]
  wire [63:0] dcache_io_cpu_s1_data_data; // @[HellaCache.scala 265:43]
  wire  dcache_io_cpu_s2_nack; // @[HellaCache.scala 265:43]
  wire  dcache_io_cpu_resp_valid; // @[HellaCache.scala 265:43]
  wire [6:0] dcache_io_cpu_resp_bits_tag; // @[HellaCache.scala 265:43]
  wire [1:0] dcache_io_cpu_resp_bits_size; // @[HellaCache.scala 265:43]
  wire [63:0] dcache_io_cpu_resp_bits_data; // @[HellaCache.scala 265:43]
  wire  dcache_io_cpu_resp_bits_replay; // @[HellaCache.scala 265:43]
  wire  dcache_io_cpu_resp_bits_has_data; // @[HellaCache.scala 265:43]
  wire [63:0] dcache_io_cpu_resp_bits_data_word_bypass; // @[HellaCache.scala 265:43]
  wire  dcache_io_cpu_replay_next; // @[HellaCache.scala 265:43]
  wire  dcache_io_cpu_s2_xcpt_ma_ld; // @[HellaCache.scala 265:43]
  wire  dcache_io_cpu_s2_xcpt_ma_st; // @[HellaCache.scala 265:43]
  wire  dcache_io_cpu_s2_xcpt_pf_ld; // @[HellaCache.scala 265:43]
  wire  dcache_io_cpu_s2_xcpt_pf_st; // @[HellaCache.scala 265:43]
  wire  dcache_io_cpu_s2_xcpt_ae_ld; // @[HellaCache.scala 265:43]
  wire  dcache_io_cpu_s2_xcpt_ae_st; // @[HellaCache.scala 265:43]
  wire  dcache_io_cpu_ordered; // @[HellaCache.scala 265:43]
  wire  dcache_io_cpu_perf_release; // @[HellaCache.scala 265:43]
  wire  dcache_io_cpu_perf_grant; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_req_ready; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_req_valid; // @[HellaCache.scala 265:43]
  wire [26:0] dcache_io_ptw_req_bits_bits_addr; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_resp_valid; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_resp_bits_ae; // @[HellaCache.scala 265:43]
  wire [53:0] dcache_io_ptw_resp_bits_pte_ppn; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_resp_bits_pte_d; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_resp_bits_pte_a; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_resp_bits_pte_g; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_resp_bits_pte_u; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_resp_bits_pte_x; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_resp_bits_pte_w; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_resp_bits_pte_r; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_resp_bits_pte_v; // @[HellaCache.scala 265:43]
  wire [1:0] dcache_io_ptw_resp_bits_level; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_resp_bits_homogeneous; // @[HellaCache.scala 265:43]
  wire [3:0] dcache_io_ptw_ptbr_mode; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_status_debug; // @[HellaCache.scala 265:43]
  wire [1:0] dcache_io_ptw_status_dprv; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_status_mxr; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_status_sum; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_pmp_0_cfg_l; // @[HellaCache.scala 265:43]
  wire [1:0] dcache_io_ptw_pmp_0_cfg_a; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_pmp_0_cfg_x; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_pmp_0_cfg_w; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_pmp_0_cfg_r; // @[HellaCache.scala 265:43]
  wire [29:0] dcache_io_ptw_pmp_0_addr; // @[HellaCache.scala 265:43]
  wire [31:0] dcache_io_ptw_pmp_0_mask; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_pmp_1_cfg_l; // @[HellaCache.scala 265:43]
  wire [1:0] dcache_io_ptw_pmp_1_cfg_a; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_pmp_1_cfg_x; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_pmp_1_cfg_w; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_pmp_1_cfg_r; // @[HellaCache.scala 265:43]
  wire [29:0] dcache_io_ptw_pmp_1_addr; // @[HellaCache.scala 265:43]
  wire [31:0] dcache_io_ptw_pmp_1_mask; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_pmp_2_cfg_l; // @[HellaCache.scala 265:43]
  wire [1:0] dcache_io_ptw_pmp_2_cfg_a; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_pmp_2_cfg_x; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_pmp_2_cfg_w; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_pmp_2_cfg_r; // @[HellaCache.scala 265:43]
  wire [29:0] dcache_io_ptw_pmp_2_addr; // @[HellaCache.scala 265:43]
  wire [31:0] dcache_io_ptw_pmp_2_mask; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_pmp_3_cfg_l; // @[HellaCache.scala 265:43]
  wire [1:0] dcache_io_ptw_pmp_3_cfg_a; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_pmp_3_cfg_x; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_pmp_3_cfg_w; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_pmp_3_cfg_r; // @[HellaCache.scala 265:43]
  wire [29:0] dcache_io_ptw_pmp_3_addr; // @[HellaCache.scala 265:43]
  wire [31:0] dcache_io_ptw_pmp_3_mask; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_pmp_4_cfg_l; // @[HellaCache.scala 265:43]
  wire [1:0] dcache_io_ptw_pmp_4_cfg_a; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_pmp_4_cfg_x; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_pmp_4_cfg_w; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_pmp_4_cfg_r; // @[HellaCache.scala 265:43]
  wire [29:0] dcache_io_ptw_pmp_4_addr; // @[HellaCache.scala 265:43]
  wire [31:0] dcache_io_ptw_pmp_4_mask; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_pmp_5_cfg_l; // @[HellaCache.scala 265:43]
  wire [1:0] dcache_io_ptw_pmp_5_cfg_a; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_pmp_5_cfg_x; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_pmp_5_cfg_w; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_pmp_5_cfg_r; // @[HellaCache.scala 265:43]
  wire [29:0] dcache_io_ptw_pmp_5_addr; // @[HellaCache.scala 265:43]
  wire [31:0] dcache_io_ptw_pmp_5_mask; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_pmp_6_cfg_l; // @[HellaCache.scala 265:43]
  wire [1:0] dcache_io_ptw_pmp_6_cfg_a; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_pmp_6_cfg_x; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_pmp_6_cfg_w; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_pmp_6_cfg_r; // @[HellaCache.scala 265:43]
  wire [29:0] dcache_io_ptw_pmp_6_addr; // @[HellaCache.scala 265:43]
  wire [31:0] dcache_io_ptw_pmp_6_mask; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_pmp_7_cfg_l; // @[HellaCache.scala 265:43]
  wire [1:0] dcache_io_ptw_pmp_7_cfg_a; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_pmp_7_cfg_x; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_pmp_7_cfg_w; // @[HellaCache.scala 265:43]
  wire  dcache_io_ptw_pmp_7_cfg_r; // @[HellaCache.scala 265:43]
  wire [29:0] dcache_io_ptw_pmp_7_addr; // @[HellaCache.scala 265:43]
  wire [31:0] dcache_io_ptw_pmp_7_mask; // @[HellaCache.scala 265:43]
  wire [29:0] dcache_io_covSum; // @[HellaCache.scala 265:43]
  wire  dcache_metaAssert; // @[HellaCache.scala 265:43]
  wire  dcache_metaReset; // @[HellaCache.scala 265:43]
  wire  dcache_data_halt; // @[HellaCache.scala 265:43]
  wire  dcache_tlb_halt; // @[HellaCache.scala 265:43]
  wire  dcache_pma_checker_halt; // @[HellaCache.scala 265:43]
  wire  dcache_lfsr_prng_halt; // @[HellaCache.scala 265:43]
  wire  frontend_gated_clock; // @[Frontend.scala 350:28]
  wire  frontend_reset; // @[Frontend.scala 350:28]
  wire  frontend_auto_icache_master_out_a_ready; // @[Frontend.scala 350:28]
  wire  frontend_auto_icache_master_out_a_valid; // @[Frontend.scala 350:28]
  wire [31:0] frontend_auto_icache_master_out_a_bits_address; // @[Frontend.scala 350:28]
  wire  frontend_auto_icache_master_out_d_valid; // @[Frontend.scala 350:28]
  wire [2:0] frontend_auto_icache_master_out_d_bits_opcode; // @[Frontend.scala 350:28]
  wire [3:0] frontend_auto_icache_master_out_d_bits_size; // @[Frontend.scala 350:28]
  wire [63:0] frontend_auto_icache_master_out_d_bits_data; // @[Frontend.scala 350:28]
  wire  frontend_auto_icache_master_out_d_bits_corrupt; // @[Frontend.scala 350:28]
  wire [31:0] frontend_auto_reset_vector_sink_in; // @[Frontend.scala 350:28]
  wire  frontend_io_cpu_might_request; // @[Frontend.scala 350:28]
  wire  frontend_io_cpu_req_valid; // @[Frontend.scala 350:28]
  wire [39:0] frontend_io_cpu_req_bits_pc; // @[Frontend.scala 350:28]
  wire  frontend_io_cpu_req_bits_speculative; // @[Frontend.scala 350:28]
  wire  frontend_io_cpu_sfence_valid; // @[Frontend.scala 350:28]
  wire  frontend_io_cpu_sfence_bits_rs1; // @[Frontend.scala 350:28]
  wire  frontend_io_cpu_sfence_bits_rs2; // @[Frontend.scala 350:28]
  wire [38:0] frontend_io_cpu_sfence_bits_addr; // @[Frontend.scala 350:28]
  wire  frontend_io_cpu_resp_ready; // @[Frontend.scala 350:28]
  wire  frontend_io_cpu_resp_valid; // @[Frontend.scala 350:28]
  wire  frontend_io_cpu_resp_bits_btb_taken; // @[Frontend.scala 350:28]
  wire  frontend_io_cpu_resp_bits_btb_bridx; // @[Frontend.scala 350:28]
  wire [4:0] frontend_io_cpu_resp_bits_btb_entry; // @[Frontend.scala 350:28]
  wire [7:0] frontend_io_cpu_resp_bits_btb_bht_history; // @[Frontend.scala 350:28]
  wire [39:0] frontend_io_cpu_resp_bits_pc; // @[Frontend.scala 350:28]
  wire [31:0] frontend_io_cpu_resp_bits_data; // @[Frontend.scala 350:28]
  wire  frontend_io_cpu_resp_bits_xcpt_pf_inst; // @[Frontend.scala 350:28]
  wire  frontend_io_cpu_resp_bits_xcpt_ae_inst; // @[Frontend.scala 350:28]
  wire  frontend_io_cpu_resp_bits_replay; // @[Frontend.scala 350:28]
  wire  frontend_io_cpu_btb_update_valid; // @[Frontend.scala 350:28]
  wire [4:0] frontend_io_cpu_btb_update_bits_prediction_entry; // @[Frontend.scala 350:28]
  wire [38:0] frontend_io_cpu_btb_update_bits_pc; // @[Frontend.scala 350:28]
  wire  frontend_io_cpu_btb_update_bits_isValid; // @[Frontend.scala 350:28]
  wire [38:0] frontend_io_cpu_btb_update_bits_br_pc; // @[Frontend.scala 350:28]
  wire [1:0] frontend_io_cpu_btb_update_bits_cfiType; // @[Frontend.scala 350:28]
  wire  frontend_io_cpu_bht_update_valid; // @[Frontend.scala 350:28]
  wire [7:0] frontend_io_cpu_bht_update_bits_prediction_history; // @[Frontend.scala 350:28]
  wire [38:0] frontend_io_cpu_bht_update_bits_pc; // @[Frontend.scala 350:28]
  wire  frontend_io_cpu_bht_update_bits_branch; // @[Frontend.scala 350:28]
  wire  frontend_io_cpu_bht_update_bits_taken; // @[Frontend.scala 350:28]
  wire  frontend_io_cpu_bht_update_bits_mispredict; // @[Frontend.scala 350:28]
  wire  frontend_io_cpu_flush_icache; // @[Frontend.scala 350:28]
  wire [39:0] frontend_io_cpu_npc; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_req_ready; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_req_valid; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_req_bits_valid; // @[Frontend.scala 350:28]
  wire [26:0] frontend_io_ptw_req_bits_bits_addr; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_resp_valid; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_resp_bits_ae; // @[Frontend.scala 350:28]
  wire [53:0] frontend_io_ptw_resp_bits_pte_ppn; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_resp_bits_pte_d; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_resp_bits_pte_a; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_resp_bits_pte_g; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_resp_bits_pte_u; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_resp_bits_pte_x; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_resp_bits_pte_w; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_resp_bits_pte_r; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_resp_bits_pte_v; // @[Frontend.scala 350:28]
  wire [1:0] frontend_io_ptw_resp_bits_level; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_resp_bits_homogeneous; // @[Frontend.scala 350:28]
  wire [3:0] frontend_io_ptw_ptbr_mode; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_status_debug; // @[Frontend.scala 350:28]
  wire [1:0] frontend_io_ptw_status_prv; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_pmp_0_cfg_l; // @[Frontend.scala 350:28]
  wire [1:0] frontend_io_ptw_pmp_0_cfg_a; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_pmp_0_cfg_x; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_pmp_0_cfg_w; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_pmp_0_cfg_r; // @[Frontend.scala 350:28]
  wire [29:0] frontend_io_ptw_pmp_0_addr; // @[Frontend.scala 350:28]
  wire [31:0] frontend_io_ptw_pmp_0_mask; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_pmp_1_cfg_l; // @[Frontend.scala 350:28]
  wire [1:0] frontend_io_ptw_pmp_1_cfg_a; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_pmp_1_cfg_x; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_pmp_1_cfg_w; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_pmp_1_cfg_r; // @[Frontend.scala 350:28]
  wire [29:0] frontend_io_ptw_pmp_1_addr; // @[Frontend.scala 350:28]
  wire [31:0] frontend_io_ptw_pmp_1_mask; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_pmp_2_cfg_l; // @[Frontend.scala 350:28]
  wire [1:0] frontend_io_ptw_pmp_2_cfg_a; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_pmp_2_cfg_x; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_pmp_2_cfg_w; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_pmp_2_cfg_r; // @[Frontend.scala 350:28]
  wire [29:0] frontend_io_ptw_pmp_2_addr; // @[Frontend.scala 350:28]
  wire [31:0] frontend_io_ptw_pmp_2_mask; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_pmp_3_cfg_l; // @[Frontend.scala 350:28]
  wire [1:0] frontend_io_ptw_pmp_3_cfg_a; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_pmp_3_cfg_x; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_pmp_3_cfg_w; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_pmp_3_cfg_r; // @[Frontend.scala 350:28]
  wire [29:0] frontend_io_ptw_pmp_3_addr; // @[Frontend.scala 350:28]
  wire [31:0] frontend_io_ptw_pmp_3_mask; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_pmp_4_cfg_l; // @[Frontend.scala 350:28]
  wire [1:0] frontend_io_ptw_pmp_4_cfg_a; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_pmp_4_cfg_x; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_pmp_4_cfg_w; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_pmp_4_cfg_r; // @[Frontend.scala 350:28]
  wire [29:0] frontend_io_ptw_pmp_4_addr; // @[Frontend.scala 350:28]
  wire [31:0] frontend_io_ptw_pmp_4_mask; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_pmp_5_cfg_l; // @[Frontend.scala 350:28]
  wire [1:0] frontend_io_ptw_pmp_5_cfg_a; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_pmp_5_cfg_x; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_pmp_5_cfg_w; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_pmp_5_cfg_r; // @[Frontend.scala 350:28]
  wire [29:0] frontend_io_ptw_pmp_5_addr; // @[Frontend.scala 350:28]
  wire [31:0] frontend_io_ptw_pmp_5_mask; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_pmp_6_cfg_l; // @[Frontend.scala 350:28]
  wire [1:0] frontend_io_ptw_pmp_6_cfg_a; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_pmp_6_cfg_x; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_pmp_6_cfg_w; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_pmp_6_cfg_r; // @[Frontend.scala 350:28]
  wire [29:0] frontend_io_ptw_pmp_6_addr; // @[Frontend.scala 350:28]
  wire [31:0] frontend_io_ptw_pmp_6_mask; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_pmp_7_cfg_l; // @[Frontend.scala 350:28]
  wire [1:0] frontend_io_ptw_pmp_7_cfg_a; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_pmp_7_cfg_x; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_pmp_7_cfg_w; // @[Frontend.scala 350:28]
  wire  frontend_io_ptw_pmp_7_cfg_r; // @[Frontend.scala 350:28]
  wire [29:0] frontend_io_ptw_pmp_7_addr; // @[Frontend.scala 350:28]
  wire [31:0] frontend_io_ptw_pmp_7_mask; // @[Frontend.scala 350:28]
  wire [63:0] frontend_io_ptw_customCSRs_csrs_0_value; // @[Frontend.scala 350:28]
  wire [29:0] frontend_io_covSum; // @[Frontend.scala 350:28]
  wire  frontend_metaAssert; // @[Frontend.scala 350:28]
  wire  frontend_metaReset; // @[Frontend.scala 350:28]
  wire  frontend_icache_halt; // @[Frontend.scala 350:28]
  wire  frontend_fq_halt; // @[Frontend.scala 350:28]
  wire  frontend_tlb_halt; // @[Frontend.scala 350:28]
  wire  frontend_btb_halt; // @[Frontend.scala 350:28]
  wire  fpuOpt_clock; // @[RocketTile.scala 202:62]
  wire  fpuOpt_reset; // @[RocketTile.scala 202:62]
  wire [31:0] fpuOpt_io_inst; // @[RocketTile.scala 202:62]
  wire [63:0] fpuOpt_io_fromint_data; // @[RocketTile.scala 202:62]
  wire [2:0] fpuOpt_io_fcsr_rm; // @[RocketTile.scala 202:62]
  wire  fpuOpt_io_fcsr_flags_valid; // @[RocketTile.scala 202:62]
  wire [4:0] fpuOpt_io_fcsr_flags_bits; // @[RocketTile.scala 202:62]
  wire [63:0] fpuOpt_io_store_data; // @[RocketTile.scala 202:62]
  wire [63:0] fpuOpt_io_toint_data; // @[RocketTile.scala 202:62]
  wire  fpuOpt_io_dmem_resp_val; // @[RocketTile.scala 202:62]
  wire [2:0] fpuOpt_io_dmem_resp_type; // @[RocketTile.scala 202:62]
  wire [4:0] fpuOpt_io_dmem_resp_tag; // @[RocketTile.scala 202:62]
  wire [63:0] fpuOpt_io_dmem_resp_data; // @[RocketTile.scala 202:62]
  wire  fpuOpt_io_valid; // @[RocketTile.scala 202:62]
  wire  fpuOpt_io_fcsr_rdy; // @[RocketTile.scala 202:62]
  wire  fpuOpt_io_nack_mem; // @[RocketTile.scala 202:62]
  wire  fpuOpt_io_illegal_rm; // @[RocketTile.scala 202:62]
  wire  fpuOpt_io_killx; // @[RocketTile.scala 202:62]
  wire  fpuOpt_io_killm; // @[RocketTile.scala 202:62]
  wire  fpuOpt_io_dec_wen; // @[RocketTile.scala 202:62]
  wire  fpuOpt_io_dec_ren1; // @[RocketTile.scala 202:62]
  wire  fpuOpt_io_dec_ren2; // @[RocketTile.scala 202:62]
  wire  fpuOpt_io_dec_ren3; // @[RocketTile.scala 202:62]
  wire  fpuOpt_io_sboard_set; // @[RocketTile.scala 202:62]
  wire  fpuOpt_io_sboard_clr; // @[RocketTile.scala 202:62]
  wire [4:0] fpuOpt_io_sboard_clra; // @[RocketTile.scala 202:62]
  wire [29:0] fpuOpt_io_covSum; // @[RocketTile.scala 202:62]
  wire  fpuOpt_metaAssert; // @[RocketTile.scala 202:62]
  wire  fpuOpt_metaReset; // @[RocketTile.scala 202:62]
  wire  fpuOpt_fpiu_halt; // @[RocketTile.scala 202:62]
  wire  fpuOpt_ifpu_halt; // @[RocketTile.scala 202:62]
  wire  fpuOpt_sfma_halt; // @[RocketTile.scala 202:62]
  wire  fpuOpt_fpmu_halt; // @[RocketTile.scala 202:62]
  wire  fpuOpt_divSqrt_1_halt; // @[RocketTile.scala 202:62]
  wire  fpuOpt_dfma_halt; // @[RocketTile.scala 202:62]
  wire  fpuOpt_divSqrt_halt; // @[RocketTile.scala 202:62]
  wire  dcacheArb_clock; // @[HellaCache.scala 276:25]
  wire  dcacheArb_io_requestor_0_req_ready; // @[HellaCache.scala 276:25]
  wire  dcacheArb_io_requestor_0_req_valid; // @[HellaCache.scala 276:25]
  wire [39:0] dcacheArb_io_requestor_0_req_bits_addr; // @[HellaCache.scala 276:25]
  wire  dcacheArb_io_requestor_0_s1_kill; // @[HellaCache.scala 276:25]
  wire  dcacheArb_io_requestor_0_s2_nack; // @[HellaCache.scala 276:25]
  wire  dcacheArb_io_requestor_0_resp_valid; // @[HellaCache.scala 276:25]
  wire [63:0] dcacheArb_io_requestor_0_resp_bits_data; // @[HellaCache.scala 276:25]
  wire  dcacheArb_io_requestor_0_s2_xcpt_ae_ld; // @[HellaCache.scala 276:25]
  wire  dcacheArb_io_requestor_1_req_ready; // @[HellaCache.scala 276:25]
  wire  dcacheArb_io_requestor_1_req_valid; // @[HellaCache.scala 276:25]
  wire [39:0] dcacheArb_io_requestor_1_req_bits_addr; // @[HellaCache.scala 276:25]
  wire [6:0] dcacheArb_io_requestor_1_req_bits_tag; // @[HellaCache.scala 276:25]
  wire [4:0] dcacheArb_io_requestor_1_req_bits_cmd; // @[HellaCache.scala 276:25]
  wire [1:0] dcacheArb_io_requestor_1_req_bits_size; // @[HellaCache.scala 276:25]
  wire  dcacheArb_io_requestor_1_req_bits_signed; // @[HellaCache.scala 276:25]
  wire  dcacheArb_io_requestor_1_s1_kill; // @[HellaCache.scala 276:25]
  wire [63:0] dcacheArb_io_requestor_1_s1_data_data; // @[HellaCache.scala 276:25]
  wire  dcacheArb_io_requestor_1_s2_nack; // @[HellaCache.scala 276:25]
  wire  dcacheArb_io_requestor_1_resp_valid; // @[HellaCache.scala 276:25]
  wire [6:0] dcacheArb_io_requestor_1_resp_bits_tag; // @[HellaCache.scala 276:25]
  wire [1:0] dcacheArb_io_requestor_1_resp_bits_size; // @[HellaCache.scala 276:25]
  wire [63:0] dcacheArb_io_requestor_1_resp_bits_data; // @[HellaCache.scala 276:25]
  wire  dcacheArb_io_requestor_1_resp_bits_replay; // @[HellaCache.scala 276:25]
  wire  dcacheArb_io_requestor_1_resp_bits_has_data; // @[HellaCache.scala 276:25]
  wire [63:0] dcacheArb_io_requestor_1_resp_bits_data_word_bypass; // @[HellaCache.scala 276:25]
  wire  dcacheArb_io_requestor_1_replay_next; // @[HellaCache.scala 276:25]
  wire  dcacheArb_io_requestor_1_s2_xcpt_ma_ld; // @[HellaCache.scala 276:25]
  wire  dcacheArb_io_requestor_1_s2_xcpt_ma_st; // @[HellaCache.scala 276:25]
  wire  dcacheArb_io_requestor_1_s2_xcpt_pf_ld; // @[HellaCache.scala 276:25]
  wire  dcacheArb_io_requestor_1_s2_xcpt_pf_st; // @[HellaCache.scala 276:25]
  wire  dcacheArb_io_requestor_1_s2_xcpt_ae_ld; // @[HellaCache.scala 276:25]
  wire  dcacheArb_io_requestor_1_s2_xcpt_ae_st; // @[HellaCache.scala 276:25]
  wire  dcacheArb_io_requestor_1_ordered; // @[HellaCache.scala 276:25]
  wire  dcacheArb_io_requestor_1_perf_release; // @[HellaCache.scala 276:25]
  wire  dcacheArb_io_requestor_1_perf_grant; // @[HellaCache.scala 276:25]
  wire  dcacheArb_io_mem_req_ready; // @[HellaCache.scala 276:25]
  wire  dcacheArb_io_mem_req_valid; // @[HellaCache.scala 276:25]
  wire [39:0] dcacheArb_io_mem_req_bits_addr; // @[HellaCache.scala 276:25]
  wire [6:0] dcacheArb_io_mem_req_bits_tag; // @[HellaCache.scala 276:25]
  wire [4:0] dcacheArb_io_mem_req_bits_cmd; // @[HellaCache.scala 276:25]
  wire [1:0] dcacheArb_io_mem_req_bits_size; // @[HellaCache.scala 276:25]
  wire  dcacheArb_io_mem_req_bits_signed; // @[HellaCache.scala 276:25]
  wire  dcacheArb_io_mem_req_bits_phys; // @[HellaCache.scala 276:25]
  wire  dcacheArb_io_mem_s1_kill; // @[HellaCache.scala 276:25]
  wire [63:0] dcacheArb_io_mem_s1_data_data; // @[HellaCache.scala 276:25]
  wire  dcacheArb_io_mem_s2_nack; // @[HellaCache.scala 276:25]
  wire  dcacheArb_io_mem_resp_valid; // @[HellaCache.scala 276:25]
  wire [6:0] dcacheArb_io_mem_resp_bits_tag; // @[HellaCache.scala 276:25]
  wire [1:0] dcacheArb_io_mem_resp_bits_size; // @[HellaCache.scala 276:25]
  wire [63:0] dcacheArb_io_mem_resp_bits_data; // @[HellaCache.scala 276:25]
  wire  dcacheArb_io_mem_resp_bits_replay; // @[HellaCache.scala 276:25]
  wire  dcacheArb_io_mem_resp_bits_has_data; // @[HellaCache.scala 276:25]
  wire [63:0] dcacheArb_io_mem_resp_bits_data_word_bypass; // @[HellaCache.scala 276:25]
  wire  dcacheArb_io_mem_replay_next; // @[HellaCache.scala 276:25]
  wire  dcacheArb_io_mem_s2_xcpt_ma_ld; // @[HellaCache.scala 276:25]
  wire  dcacheArb_io_mem_s2_xcpt_ma_st; // @[HellaCache.scala 276:25]
  wire  dcacheArb_io_mem_s2_xcpt_pf_ld; // @[HellaCache.scala 276:25]
  wire  dcacheArb_io_mem_s2_xcpt_pf_st; // @[HellaCache.scala 276:25]
  wire  dcacheArb_io_mem_s2_xcpt_ae_ld; // @[HellaCache.scala 276:25]
  wire  dcacheArb_io_mem_s2_xcpt_ae_st; // @[HellaCache.scala 276:25]
  wire  dcacheArb_io_mem_ordered; // @[HellaCache.scala 276:25]
  wire  dcacheArb_io_mem_perf_release; // @[HellaCache.scala 276:25]
  wire  dcacheArb_io_mem_perf_grant; // @[HellaCache.scala 276:25]
  wire [29:0] dcacheArb_io_covSum; // @[HellaCache.scala 276:25]
  wire  dcacheArb_metaAssert; // @[HellaCache.scala 276:25]
  wire  dcacheArb_metaReset; // @[HellaCache.scala 276:25]
  wire  ptw_clock; // @[PTW.scala 439:19]
  wire  ptw_reset; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_req_ready; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_req_valid; // @[PTW.scala 439:19]
  wire [26:0] ptw_io_requestor_0_req_bits_bits_addr; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_resp_valid; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_resp_bits_ae; // @[PTW.scala 439:19]
  wire [53:0] ptw_io_requestor_0_resp_bits_pte_ppn; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_resp_bits_pte_d; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_resp_bits_pte_a; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_resp_bits_pte_g; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_resp_bits_pte_u; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_resp_bits_pte_x; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_resp_bits_pte_w; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_resp_bits_pte_r; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_resp_bits_pte_v; // @[PTW.scala 439:19]
  wire [1:0] ptw_io_requestor_0_resp_bits_level; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_resp_bits_homogeneous; // @[PTW.scala 439:19]
  wire [3:0] ptw_io_requestor_0_ptbr_mode; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_status_debug; // @[PTW.scala 439:19]
  wire [1:0] ptw_io_requestor_0_status_dprv; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_status_mxr; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_status_sum; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_pmp_0_cfg_l; // @[PTW.scala 439:19]
  wire [1:0] ptw_io_requestor_0_pmp_0_cfg_a; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_pmp_0_cfg_x; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_pmp_0_cfg_w; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_pmp_0_cfg_r; // @[PTW.scala 439:19]
  wire [29:0] ptw_io_requestor_0_pmp_0_addr; // @[PTW.scala 439:19]
  wire [31:0] ptw_io_requestor_0_pmp_0_mask; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_pmp_1_cfg_l; // @[PTW.scala 439:19]
  wire [1:0] ptw_io_requestor_0_pmp_1_cfg_a; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_pmp_1_cfg_x; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_pmp_1_cfg_w; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_pmp_1_cfg_r; // @[PTW.scala 439:19]
  wire [29:0] ptw_io_requestor_0_pmp_1_addr; // @[PTW.scala 439:19]
  wire [31:0] ptw_io_requestor_0_pmp_1_mask; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_pmp_2_cfg_l; // @[PTW.scala 439:19]
  wire [1:0] ptw_io_requestor_0_pmp_2_cfg_a; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_pmp_2_cfg_x; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_pmp_2_cfg_w; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_pmp_2_cfg_r; // @[PTW.scala 439:19]
  wire [29:0] ptw_io_requestor_0_pmp_2_addr; // @[PTW.scala 439:19]
  wire [31:0] ptw_io_requestor_0_pmp_2_mask; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_pmp_3_cfg_l; // @[PTW.scala 439:19]
  wire [1:0] ptw_io_requestor_0_pmp_3_cfg_a; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_pmp_3_cfg_x; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_pmp_3_cfg_w; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_pmp_3_cfg_r; // @[PTW.scala 439:19]
  wire [29:0] ptw_io_requestor_0_pmp_3_addr; // @[PTW.scala 439:19]
  wire [31:0] ptw_io_requestor_0_pmp_3_mask; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_pmp_4_cfg_l; // @[PTW.scala 439:19]
  wire [1:0] ptw_io_requestor_0_pmp_4_cfg_a; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_pmp_4_cfg_x; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_pmp_4_cfg_w; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_pmp_4_cfg_r; // @[PTW.scala 439:19]
  wire [29:0] ptw_io_requestor_0_pmp_4_addr; // @[PTW.scala 439:19]
  wire [31:0] ptw_io_requestor_0_pmp_4_mask; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_pmp_5_cfg_l; // @[PTW.scala 439:19]
  wire [1:0] ptw_io_requestor_0_pmp_5_cfg_a; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_pmp_5_cfg_x; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_pmp_5_cfg_w; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_pmp_5_cfg_r; // @[PTW.scala 439:19]
  wire [29:0] ptw_io_requestor_0_pmp_5_addr; // @[PTW.scala 439:19]
  wire [31:0] ptw_io_requestor_0_pmp_5_mask; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_pmp_6_cfg_l; // @[PTW.scala 439:19]
  wire [1:0] ptw_io_requestor_0_pmp_6_cfg_a; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_pmp_6_cfg_x; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_pmp_6_cfg_w; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_pmp_6_cfg_r; // @[PTW.scala 439:19]
  wire [29:0] ptw_io_requestor_0_pmp_6_addr; // @[PTW.scala 439:19]
  wire [31:0] ptw_io_requestor_0_pmp_6_mask; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_pmp_7_cfg_l; // @[PTW.scala 439:19]
  wire [1:0] ptw_io_requestor_0_pmp_7_cfg_a; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_pmp_7_cfg_x; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_pmp_7_cfg_w; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_0_pmp_7_cfg_r; // @[PTW.scala 439:19]
  wire [29:0] ptw_io_requestor_0_pmp_7_addr; // @[PTW.scala 439:19]
  wire [31:0] ptw_io_requestor_0_pmp_7_mask; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_req_ready; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_req_valid; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_req_bits_valid; // @[PTW.scala 439:19]
  wire [26:0] ptw_io_requestor_1_req_bits_bits_addr; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_resp_valid; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_resp_bits_ae; // @[PTW.scala 439:19]
  wire [53:0] ptw_io_requestor_1_resp_bits_pte_ppn; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_resp_bits_pte_d; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_resp_bits_pte_a; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_resp_bits_pte_g; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_resp_bits_pte_u; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_resp_bits_pte_x; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_resp_bits_pte_w; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_resp_bits_pte_r; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_resp_bits_pte_v; // @[PTW.scala 439:19]
  wire [1:0] ptw_io_requestor_1_resp_bits_level; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_resp_bits_homogeneous; // @[PTW.scala 439:19]
  wire [3:0] ptw_io_requestor_1_ptbr_mode; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_status_debug; // @[PTW.scala 439:19]
  wire [1:0] ptw_io_requestor_1_status_prv; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_pmp_0_cfg_l; // @[PTW.scala 439:19]
  wire [1:0] ptw_io_requestor_1_pmp_0_cfg_a; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_pmp_0_cfg_x; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_pmp_0_cfg_w; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_pmp_0_cfg_r; // @[PTW.scala 439:19]
  wire [29:0] ptw_io_requestor_1_pmp_0_addr; // @[PTW.scala 439:19]
  wire [31:0] ptw_io_requestor_1_pmp_0_mask; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_pmp_1_cfg_l; // @[PTW.scala 439:19]
  wire [1:0] ptw_io_requestor_1_pmp_1_cfg_a; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_pmp_1_cfg_x; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_pmp_1_cfg_w; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_pmp_1_cfg_r; // @[PTW.scala 439:19]
  wire [29:0] ptw_io_requestor_1_pmp_1_addr; // @[PTW.scala 439:19]
  wire [31:0] ptw_io_requestor_1_pmp_1_mask; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_pmp_2_cfg_l; // @[PTW.scala 439:19]
  wire [1:0] ptw_io_requestor_1_pmp_2_cfg_a; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_pmp_2_cfg_x; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_pmp_2_cfg_w; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_pmp_2_cfg_r; // @[PTW.scala 439:19]
  wire [29:0] ptw_io_requestor_1_pmp_2_addr; // @[PTW.scala 439:19]
  wire [31:0] ptw_io_requestor_1_pmp_2_mask; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_pmp_3_cfg_l; // @[PTW.scala 439:19]
  wire [1:0] ptw_io_requestor_1_pmp_3_cfg_a; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_pmp_3_cfg_x; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_pmp_3_cfg_w; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_pmp_3_cfg_r; // @[PTW.scala 439:19]
  wire [29:0] ptw_io_requestor_1_pmp_3_addr; // @[PTW.scala 439:19]
  wire [31:0] ptw_io_requestor_1_pmp_3_mask; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_pmp_4_cfg_l; // @[PTW.scala 439:19]
  wire [1:0] ptw_io_requestor_1_pmp_4_cfg_a; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_pmp_4_cfg_x; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_pmp_4_cfg_w; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_pmp_4_cfg_r; // @[PTW.scala 439:19]
  wire [29:0] ptw_io_requestor_1_pmp_4_addr; // @[PTW.scala 439:19]
  wire [31:0] ptw_io_requestor_1_pmp_4_mask; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_pmp_5_cfg_l; // @[PTW.scala 439:19]
  wire [1:0] ptw_io_requestor_1_pmp_5_cfg_a; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_pmp_5_cfg_x; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_pmp_5_cfg_w; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_pmp_5_cfg_r; // @[PTW.scala 439:19]
  wire [29:0] ptw_io_requestor_1_pmp_5_addr; // @[PTW.scala 439:19]
  wire [31:0] ptw_io_requestor_1_pmp_5_mask; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_pmp_6_cfg_l; // @[PTW.scala 439:19]
  wire [1:0] ptw_io_requestor_1_pmp_6_cfg_a; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_pmp_6_cfg_x; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_pmp_6_cfg_w; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_pmp_6_cfg_r; // @[PTW.scala 439:19]
  wire [29:0] ptw_io_requestor_1_pmp_6_addr; // @[PTW.scala 439:19]
  wire [31:0] ptw_io_requestor_1_pmp_6_mask; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_pmp_7_cfg_l; // @[PTW.scala 439:19]
  wire [1:0] ptw_io_requestor_1_pmp_7_cfg_a; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_pmp_7_cfg_x; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_pmp_7_cfg_w; // @[PTW.scala 439:19]
  wire  ptw_io_requestor_1_pmp_7_cfg_r; // @[PTW.scala 439:19]
  wire [29:0] ptw_io_requestor_1_pmp_7_addr; // @[PTW.scala 439:19]
  wire [31:0] ptw_io_requestor_1_pmp_7_mask; // @[PTW.scala 439:19]
  wire [63:0] ptw_io_requestor_1_customCSRs_csrs_0_value; // @[PTW.scala 439:19]
  wire  ptw_io_mem_req_ready; // @[PTW.scala 439:19]
  wire  ptw_io_mem_req_valid; // @[PTW.scala 439:19]
  wire [39:0] ptw_io_mem_req_bits_addr; // @[PTW.scala 439:19]
  wire  ptw_io_mem_s1_kill; // @[PTW.scala 439:19]
  wire  ptw_io_mem_s2_nack; // @[PTW.scala 439:19]
  wire  ptw_io_mem_resp_valid; // @[PTW.scala 439:19]
  wire [63:0] ptw_io_mem_resp_bits_data; // @[PTW.scala 439:19]
  wire  ptw_io_mem_s2_xcpt_ae_ld; // @[PTW.scala 439:19]
  wire [3:0] ptw_io_dpath_ptbr_mode; // @[PTW.scala 439:19]
  wire [43:0] ptw_io_dpath_ptbr_ppn; // @[PTW.scala 439:19]
  wire  ptw_io_dpath_sfence_valid; // @[PTW.scala 439:19]
  wire  ptw_io_dpath_sfence_bits_rs1; // @[PTW.scala 439:19]
  wire  ptw_io_dpath_status_debug; // @[PTW.scala 439:19]
  wire [1:0] ptw_io_dpath_status_dprv; // @[PTW.scala 439:19]
  wire [1:0] ptw_io_dpath_status_prv; // @[PTW.scala 439:19]
  wire  ptw_io_dpath_status_mxr; // @[PTW.scala 439:19]
  wire  ptw_io_dpath_status_sum; // @[PTW.scala 439:19]
  wire  ptw_io_dpath_pmp_0_cfg_l; // @[PTW.scala 439:19]
  wire [1:0] ptw_io_dpath_pmp_0_cfg_a; // @[PTW.scala 439:19]
  wire  ptw_io_dpath_pmp_0_cfg_x; // @[PTW.scala 439:19]
  wire  ptw_io_dpath_pmp_0_cfg_w; // @[PTW.scala 439:19]
  wire  ptw_io_dpath_pmp_0_cfg_r; // @[PTW.scala 439:19]
  wire [29:0] ptw_io_dpath_pmp_0_addr; // @[PTW.scala 439:19]
  wire [31:0] ptw_io_dpath_pmp_0_mask; // @[PTW.scala 439:19]
  wire  ptw_io_dpath_pmp_1_cfg_l; // @[PTW.scala 439:19]
  wire [1:0] ptw_io_dpath_pmp_1_cfg_a; // @[PTW.scala 439:19]
  wire  ptw_io_dpath_pmp_1_cfg_x; // @[PTW.scala 439:19]
  wire  ptw_io_dpath_pmp_1_cfg_w; // @[PTW.scala 439:19]
  wire  ptw_io_dpath_pmp_1_cfg_r; // @[PTW.scala 439:19]
  wire [29:0] ptw_io_dpath_pmp_1_addr; // @[PTW.scala 439:19]
  wire [31:0] ptw_io_dpath_pmp_1_mask; // @[PTW.scala 439:19]
  wire  ptw_io_dpath_pmp_2_cfg_l; // @[PTW.scala 439:19]
  wire [1:0] ptw_io_dpath_pmp_2_cfg_a; // @[PTW.scala 439:19]
  wire  ptw_io_dpath_pmp_2_cfg_x; // @[PTW.scala 439:19]
  wire  ptw_io_dpath_pmp_2_cfg_w; // @[PTW.scala 439:19]
  wire  ptw_io_dpath_pmp_2_cfg_r; // @[PTW.scala 439:19]
  wire [29:0] ptw_io_dpath_pmp_2_addr; // @[PTW.scala 439:19]
  wire [31:0] ptw_io_dpath_pmp_2_mask; // @[PTW.scala 439:19]
  wire  ptw_io_dpath_pmp_3_cfg_l; // @[PTW.scala 439:19]
  wire [1:0] ptw_io_dpath_pmp_3_cfg_a; // @[PTW.scala 439:19]
  wire  ptw_io_dpath_pmp_3_cfg_x; // @[PTW.scala 439:19]
  wire  ptw_io_dpath_pmp_3_cfg_w; // @[PTW.scala 439:19]
  wire  ptw_io_dpath_pmp_3_cfg_r; // @[PTW.scala 439:19]
  wire [29:0] ptw_io_dpath_pmp_3_addr; // @[PTW.scala 439:19]
  wire [31:0] ptw_io_dpath_pmp_3_mask; // @[PTW.scala 439:19]
  wire  ptw_io_dpath_pmp_4_cfg_l; // @[PTW.scala 439:19]
  wire [1:0] ptw_io_dpath_pmp_4_cfg_a; // @[PTW.scala 439:19]
  wire  ptw_io_dpath_pmp_4_cfg_x; // @[PTW.scala 439:19]
  wire  ptw_io_dpath_pmp_4_cfg_w; // @[PTW.scala 439:19]
  wire  ptw_io_dpath_pmp_4_cfg_r; // @[PTW.scala 439:19]
  wire [29:0] ptw_io_dpath_pmp_4_addr; // @[PTW.scala 439:19]
  wire [31:0] ptw_io_dpath_pmp_4_mask; // @[PTW.scala 439:19]
  wire  ptw_io_dpath_pmp_5_cfg_l; // @[PTW.scala 439:19]
  wire [1:0] ptw_io_dpath_pmp_5_cfg_a; // @[PTW.scala 439:19]
  wire  ptw_io_dpath_pmp_5_cfg_x; // @[PTW.scala 439:19]
  wire  ptw_io_dpath_pmp_5_cfg_w; // @[PTW.scala 439:19]
  wire  ptw_io_dpath_pmp_5_cfg_r; // @[PTW.scala 439:19]
  wire [29:0] ptw_io_dpath_pmp_5_addr; // @[PTW.scala 439:19]
  wire [31:0] ptw_io_dpath_pmp_5_mask; // @[PTW.scala 439:19]
  wire  ptw_io_dpath_pmp_6_cfg_l; // @[PTW.scala 439:19]
  wire [1:0] ptw_io_dpath_pmp_6_cfg_a; // @[PTW.scala 439:19]
  wire  ptw_io_dpath_pmp_6_cfg_x; // @[PTW.scala 439:19]
  wire  ptw_io_dpath_pmp_6_cfg_w; // @[PTW.scala 439:19]
  wire  ptw_io_dpath_pmp_6_cfg_r; // @[PTW.scala 439:19]
  wire [29:0] ptw_io_dpath_pmp_6_addr; // @[PTW.scala 439:19]
  wire [31:0] ptw_io_dpath_pmp_6_mask; // @[PTW.scala 439:19]
  wire  ptw_io_dpath_pmp_7_cfg_l; // @[PTW.scala 439:19]
  wire [1:0] ptw_io_dpath_pmp_7_cfg_a; // @[PTW.scala 439:19]
  wire  ptw_io_dpath_pmp_7_cfg_x; // @[PTW.scala 439:19]
  wire  ptw_io_dpath_pmp_7_cfg_w; // @[PTW.scala 439:19]
  wire  ptw_io_dpath_pmp_7_cfg_r; // @[PTW.scala 439:19]
  wire [29:0] ptw_io_dpath_pmp_7_addr; // @[PTW.scala 439:19]
  wire [31:0] ptw_io_dpath_pmp_7_mask; // @[PTW.scala 439:19]
  wire  ptw_io_dpath_perf_l2hit; // @[PTW.scala 439:19]
  wire  ptw_io_dpath_perf_pte_miss; // @[PTW.scala 439:19]
  wire  ptw_io_dpath_perf_pte_hit; // @[PTW.scala 439:19]
  wire [63:0] ptw_io_dpath_customCSRs_csrs_0_value; // @[PTW.scala 439:19]
  wire [29:0] ptw_io_covSum; // @[PTW.scala 439:19]
  wire  ptw_metaAssert; // @[PTW.scala 439:19]
  wire  ptw_metaReset; // @[PTW.scala 439:19]
  wire  core_clock; // @[RocketTile.scala 140:20]
  wire  core_reset; // @[RocketTile.scala 140:20]
  wire  core_io_hartid; // @[RocketTile.scala 140:20]
  wire  core_io_interrupts_debug; // @[RocketTile.scala 140:20]
  wire  core_io_interrupts_mtip; // @[RocketTile.scala 140:20]
  wire  core_io_interrupts_msip; // @[RocketTile.scala 140:20]
  wire  core_io_interrupts_meip; // @[RocketTile.scala 140:20]
  wire  core_io_interrupts_seip; // @[RocketTile.scala 140:20]
  wire  core_io_imem_might_request; // @[RocketTile.scala 140:20]
  wire  core_io_imem_req_valid; // @[RocketTile.scala 140:20]
  wire [39:0] core_io_imem_req_bits_pc; // @[RocketTile.scala 140:20]
  wire  core_io_imem_req_bits_speculative; // @[RocketTile.scala 140:20]
  wire  core_io_imem_sfence_valid; // @[RocketTile.scala 140:20]
  wire  core_io_imem_sfence_bits_rs1; // @[RocketTile.scala 140:20]
  wire  core_io_imem_sfence_bits_rs2; // @[RocketTile.scala 140:20]
  wire [38:0] core_io_imem_sfence_bits_addr; // @[RocketTile.scala 140:20]
  wire  core_io_imem_resp_ready; // @[RocketTile.scala 140:20]
  wire  core_io_imem_resp_valid; // @[RocketTile.scala 140:20]
  wire  core_io_imem_resp_bits_btb_taken; // @[RocketTile.scala 140:20]
  wire  core_io_imem_resp_bits_btb_bridx; // @[RocketTile.scala 140:20]
  wire [4:0] core_io_imem_resp_bits_btb_entry; // @[RocketTile.scala 140:20]
  wire [7:0] core_io_imem_resp_bits_btb_bht_history; // @[RocketTile.scala 140:20]
  wire [39:0] core_io_imem_resp_bits_pc; // @[RocketTile.scala 140:20]
  wire [31:0] core_io_imem_resp_bits_data; // @[RocketTile.scala 140:20]
  wire  core_io_imem_resp_bits_xcpt_pf_inst; // @[RocketTile.scala 140:20]
  wire  core_io_imem_resp_bits_xcpt_ae_inst; // @[RocketTile.scala 140:20]
  wire  core_io_imem_resp_bits_replay; // @[RocketTile.scala 140:20]
  wire  core_io_imem_btb_update_valid; // @[RocketTile.scala 140:20]
  wire [4:0] core_io_imem_btb_update_bits_prediction_entry; // @[RocketTile.scala 140:20]
  wire [38:0] core_io_imem_btb_update_bits_pc; // @[RocketTile.scala 140:20]
  wire  core_io_imem_btb_update_bits_isValid; // @[RocketTile.scala 140:20]
  wire [38:0] core_io_imem_btb_update_bits_br_pc; // @[RocketTile.scala 140:20]
  wire [1:0] core_io_imem_btb_update_bits_cfiType; // @[RocketTile.scala 140:20]
  wire  core_io_imem_bht_update_valid; // @[RocketTile.scala 140:20]
  wire [7:0] core_io_imem_bht_update_bits_prediction_history; // @[RocketTile.scala 140:20]
  wire [38:0] core_io_imem_bht_update_bits_pc; // @[RocketTile.scala 140:20]
  wire  core_io_imem_bht_update_bits_branch; // @[RocketTile.scala 140:20]
  wire  core_io_imem_bht_update_bits_taken; // @[RocketTile.scala 140:20]
  wire  core_io_imem_bht_update_bits_mispredict; // @[RocketTile.scala 140:20]
  wire  core_io_imem_flush_icache; // @[RocketTile.scala 140:20]
  wire  core_io_dmem_req_ready; // @[RocketTile.scala 140:20]
  wire  core_io_dmem_req_valid; // @[RocketTile.scala 140:20]
  wire [39:0] core_io_dmem_req_bits_addr; // @[RocketTile.scala 140:20]
  wire [6:0] core_io_dmem_req_bits_tag; // @[RocketTile.scala 140:20]
  wire [4:0] core_io_dmem_req_bits_cmd; // @[RocketTile.scala 140:20]
  wire [1:0] core_io_dmem_req_bits_size; // @[RocketTile.scala 140:20]
  wire  core_io_dmem_req_bits_signed; // @[RocketTile.scala 140:20]
  wire  core_io_dmem_s1_kill; // @[RocketTile.scala 140:20]
  wire [63:0] core_io_dmem_s1_data_data; // @[RocketTile.scala 140:20]
  wire  core_io_dmem_s2_nack; // @[RocketTile.scala 140:20]
  wire  core_io_dmem_resp_valid; // @[RocketTile.scala 140:20]
  wire [6:0] core_io_dmem_resp_bits_tag; // @[RocketTile.scala 140:20]
  wire [1:0] core_io_dmem_resp_bits_size; // @[RocketTile.scala 140:20]
  wire [63:0] core_io_dmem_resp_bits_data; // @[RocketTile.scala 140:20]
  wire  core_io_dmem_resp_bits_replay; // @[RocketTile.scala 140:20]
  wire  core_io_dmem_resp_bits_has_data; // @[RocketTile.scala 140:20]
  wire [63:0] core_io_dmem_resp_bits_data_word_bypass; // @[RocketTile.scala 140:20]
  wire  core_io_dmem_replay_next; // @[RocketTile.scala 140:20]
  wire  core_io_dmem_s2_xcpt_ma_ld; // @[RocketTile.scala 140:20]
  wire  core_io_dmem_s2_xcpt_ma_st; // @[RocketTile.scala 140:20]
  wire  core_io_dmem_s2_xcpt_pf_ld; // @[RocketTile.scala 140:20]
  wire  core_io_dmem_s2_xcpt_pf_st; // @[RocketTile.scala 140:20]
  wire  core_io_dmem_s2_xcpt_ae_ld; // @[RocketTile.scala 140:20]
  wire  core_io_dmem_s2_xcpt_ae_st; // @[RocketTile.scala 140:20]
  wire  core_io_dmem_ordered; // @[RocketTile.scala 140:20]
  wire  core_io_dmem_perf_release; // @[RocketTile.scala 140:20]
  wire  core_io_dmem_perf_grant; // @[RocketTile.scala 140:20]
  wire [3:0] core_io_ptw_ptbr_mode; // @[RocketTile.scala 140:20]
  wire [43:0] core_io_ptw_ptbr_ppn; // @[RocketTile.scala 140:20]
  wire  core_io_ptw_sfence_valid; // @[RocketTile.scala 140:20]
  wire  core_io_ptw_sfence_bits_rs1; // @[RocketTile.scala 140:20]
  wire  core_io_ptw_status_debug; // @[RocketTile.scala 140:20]
  wire [1:0] core_io_ptw_status_dprv; // @[RocketTile.scala 140:20]
  wire [1:0] core_io_ptw_status_prv; // @[RocketTile.scala 140:20]
  wire  core_io_ptw_status_mxr; // @[RocketTile.scala 140:20]
  wire  core_io_ptw_status_sum; // @[RocketTile.scala 140:20]
  wire  core_io_ptw_pmp_0_cfg_l; // @[RocketTile.scala 140:20]
  wire [1:0] core_io_ptw_pmp_0_cfg_a; // @[RocketTile.scala 140:20]
  wire  core_io_ptw_pmp_0_cfg_x; // @[RocketTile.scala 140:20]
  wire  core_io_ptw_pmp_0_cfg_w; // @[RocketTile.scala 140:20]
  wire  core_io_ptw_pmp_0_cfg_r; // @[RocketTile.scala 140:20]
  wire [29:0] core_io_ptw_pmp_0_addr; // @[RocketTile.scala 140:20]
  wire [31:0] core_io_ptw_pmp_0_mask; // @[RocketTile.scala 140:20]
  wire  core_io_ptw_pmp_1_cfg_l; // @[RocketTile.scala 140:20]
  wire [1:0] core_io_ptw_pmp_1_cfg_a; // @[RocketTile.scala 140:20]
  wire  core_io_ptw_pmp_1_cfg_x; // @[RocketTile.scala 140:20]
  wire  core_io_ptw_pmp_1_cfg_w; // @[RocketTile.scala 140:20]
  wire  core_io_ptw_pmp_1_cfg_r; // @[RocketTile.scala 140:20]
  wire [29:0] core_io_ptw_pmp_1_addr; // @[RocketTile.scala 140:20]
  wire [31:0] core_io_ptw_pmp_1_mask; // @[RocketTile.scala 140:20]
  wire  core_io_ptw_pmp_2_cfg_l; // @[RocketTile.scala 140:20]
  wire [1:0] core_io_ptw_pmp_2_cfg_a; // @[RocketTile.scala 140:20]
  wire  core_io_ptw_pmp_2_cfg_x; // @[RocketTile.scala 140:20]
  wire  core_io_ptw_pmp_2_cfg_w; // @[RocketTile.scala 140:20]
  wire  core_io_ptw_pmp_2_cfg_r; // @[RocketTile.scala 140:20]
  wire [29:0] core_io_ptw_pmp_2_addr; // @[RocketTile.scala 140:20]
  wire [31:0] core_io_ptw_pmp_2_mask; // @[RocketTile.scala 140:20]
  wire  core_io_ptw_pmp_3_cfg_l; // @[RocketTile.scala 140:20]
  wire [1:0] core_io_ptw_pmp_3_cfg_a; // @[RocketTile.scala 140:20]
  wire  core_io_ptw_pmp_3_cfg_x; // @[RocketTile.scala 140:20]
  wire  core_io_ptw_pmp_3_cfg_w; // @[RocketTile.scala 140:20]
  wire  core_io_ptw_pmp_3_cfg_r; // @[RocketTile.scala 140:20]
  wire [29:0] core_io_ptw_pmp_3_addr; // @[RocketTile.scala 140:20]
  wire [31:0] core_io_ptw_pmp_3_mask; // @[RocketTile.scala 140:20]
  wire  core_io_ptw_pmp_4_cfg_l; // @[RocketTile.scala 140:20]
  wire [1:0] core_io_ptw_pmp_4_cfg_a; // @[RocketTile.scala 140:20]
  wire  core_io_ptw_pmp_4_cfg_x; // @[RocketTile.scala 140:20]
  wire  core_io_ptw_pmp_4_cfg_w; // @[RocketTile.scala 140:20]
  wire  core_io_ptw_pmp_4_cfg_r; // @[RocketTile.scala 140:20]
  wire [29:0] core_io_ptw_pmp_4_addr; // @[RocketTile.scala 140:20]
  wire [31:0] core_io_ptw_pmp_4_mask; // @[RocketTile.scala 140:20]
  wire  core_io_ptw_pmp_5_cfg_l; // @[RocketTile.scala 140:20]
  wire [1:0] core_io_ptw_pmp_5_cfg_a; // @[RocketTile.scala 140:20]
  wire  core_io_ptw_pmp_5_cfg_x; // @[RocketTile.scala 140:20]
  wire  core_io_ptw_pmp_5_cfg_w; // @[RocketTile.scala 140:20]
  wire  core_io_ptw_pmp_5_cfg_r; // @[RocketTile.scala 140:20]
  wire [29:0] core_io_ptw_pmp_5_addr; // @[RocketTile.scala 140:20]
  wire [31:0] core_io_ptw_pmp_5_mask; // @[RocketTile.scala 140:20]
  wire  core_io_ptw_pmp_6_cfg_l; // @[RocketTile.scala 140:20]
  wire [1:0] core_io_ptw_pmp_6_cfg_a; // @[RocketTile.scala 140:20]
  wire  core_io_ptw_pmp_6_cfg_x; // @[RocketTile.scala 140:20]
  wire  core_io_ptw_pmp_6_cfg_w; // @[RocketTile.scala 140:20]
  wire  core_io_ptw_pmp_6_cfg_r; // @[RocketTile.scala 140:20]
  wire [29:0] core_io_ptw_pmp_6_addr; // @[RocketTile.scala 140:20]
  wire [31:0] core_io_ptw_pmp_6_mask; // @[RocketTile.scala 140:20]
  wire  core_io_ptw_pmp_7_cfg_l; // @[RocketTile.scala 140:20]
  wire [1:0] core_io_ptw_pmp_7_cfg_a; // @[RocketTile.scala 140:20]
  wire  core_io_ptw_pmp_7_cfg_x; // @[RocketTile.scala 140:20]
  wire  core_io_ptw_pmp_7_cfg_w; // @[RocketTile.scala 140:20]
  wire  core_io_ptw_pmp_7_cfg_r; // @[RocketTile.scala 140:20]
  wire [29:0] core_io_ptw_pmp_7_addr; // @[RocketTile.scala 140:20]
  wire [31:0] core_io_ptw_pmp_7_mask; // @[RocketTile.scala 140:20]
  wire [63:0] core_io_ptw_customCSRs_csrs_0_value; // @[RocketTile.scala 140:20]
  wire [31:0] core_io_fpu_inst; // @[RocketTile.scala 140:20]
  wire [63:0] core_io_fpu_fromint_data; // @[RocketTile.scala 140:20]
  wire [2:0] core_io_fpu_fcsr_rm; // @[RocketTile.scala 140:20]
  wire  core_io_fpu_fcsr_flags_valid; // @[RocketTile.scala 140:20]
  wire [4:0] core_io_fpu_fcsr_flags_bits; // @[RocketTile.scala 140:20]
  wire [63:0] core_io_fpu_store_data; // @[RocketTile.scala 140:20]
  wire [63:0] core_io_fpu_toint_data; // @[RocketTile.scala 140:20]
  wire  core_io_fpu_dmem_resp_val; // @[RocketTile.scala 140:20]
  wire [2:0] core_io_fpu_dmem_resp_type; // @[RocketTile.scala 140:20]
  wire [4:0] core_io_fpu_dmem_resp_tag; // @[RocketTile.scala 140:20]
  wire [63:0] core_io_fpu_dmem_resp_data; // @[RocketTile.scala 140:20]
  wire  core_io_fpu_valid; // @[RocketTile.scala 140:20]
  wire  core_io_fpu_fcsr_rdy; // @[RocketTile.scala 140:20]
  wire  core_io_fpu_nack_mem; // @[RocketTile.scala 140:20]
  wire  core_io_fpu_illegal_rm; // @[RocketTile.scala 140:20]
  wire  core_io_fpu_killx; // @[RocketTile.scala 140:20]
  wire  core_io_fpu_killm; // @[RocketTile.scala 140:20]
  wire  core_io_fpu_dec_wen; // @[RocketTile.scala 140:20]
  wire  core_io_fpu_dec_ren1; // @[RocketTile.scala 140:20]
  wire  core_io_fpu_dec_ren2; // @[RocketTile.scala 140:20]
  wire  core_io_fpu_dec_ren3; // @[RocketTile.scala 140:20]
  wire  core_io_fpu_sboard_set; // @[RocketTile.scala 140:20]
  wire  core_io_fpu_sboard_clr; // @[RocketTile.scala 140:20]
  wire [4:0] core_io_fpu_sboard_clra; // @[RocketTile.scala 140:20]
  wire  core_io_trace_0_valid; // @[RocketTile.scala 140:20]
  wire [39:0] core_io_trace_0_iaddr; // @[RocketTile.scala 140:20]
  wire [31:0] core_io_trace_0_insn; // @[RocketTile.scala 140:20]
  wire [2:0] core_io_trace_0_priv; // @[RocketTile.scala 140:20]
  wire  core_io_trace_0_exception; // @[RocketTile.scala 140:20]
  wire  core_io_trace_0_interrupt; // @[RocketTile.scala 140:20]
  wire [63:0] core_io_trace_0_cause; // @[RocketTile.scala 140:20]
  wire [39:0] core_io_trace_0_tval; // @[RocketTile.scala 140:20]
  wire  core_io_wfi; // @[RocketTile.scala 140:20]
  wire [29:0] core_io_covSum; // @[RocketTile.scala 140:20]
  wire  core_metaAssert; // @[RocketTile.scala 140:20]
  wire  core_metaReset; // @[RocketTile.scala 140:20]
  wire  core_PlusArgTimeout_halt; // @[RocketTile.scala 140:20]
  wire  core_csr_halt; // @[RocketTile.scala 140:20]
  wire  core_ibuf_halt; // @[RocketTile.scala 140:20]
  wire  core_div_halt; // @[RocketTile.scala 140:20]
  reg  bundleOut_0_0_REG; // @[Interrupts.scala 129:36]
  reg [31:0] _RAND_0;
  wire [29:0] RocketTile_covSum;
  wire [29:0] tlMasterXbar_sum;
  wire [29:0] intXbar_sum;
  wire [29:0] fpuOpt_sum;
  wire [29:0] dcacheArb_sum;
  wire [29:0] frontend_sum;
  wire [29:0] dcache_sum;
  wire [29:0] broadcast_3_sum;
  wire [29:0] core_sum;
  wire [29:0] broadcast_sum;
  wire [29:0] broadcast_1_sum;
  wire [29:0] ptw_sum;
  wire  ptw_metaAssert_wire;
  wire  fpuOpt_metaAssert_wire;
  wire  frontend_metaAssert_wire;
  wire  dcacheArb_metaAssert_wire;
  wire  broadcast_1_metaAssert_wire;
  wire  broadcast_3_metaAssert_wire;
  wire  intXbar_metaAssert_wire;
  wire  core_metaAssert_wire;
  wire  tlMasterXbar_metaAssert_wire;
  wire  dcache_metaAssert_wire;
  wire  broadcast_metaAssert_wire;
  wire  RocketTile_or3;
  wire  RocketTile_or10;
  wire  RocketTile_or4;
  wire  RocketTile_or1;
  wire  RocketTile_or12;
  wire  RocketTile_or5;
  wire  RocketTile_or14;
  wire  RocketTile_or6;
  wire  RocketTile_or2;
  wire  RocketTile_or0;
  reg  RocketTile_metaAssert;
  reg [31:0] _RAND_1;
  TLXbar_7 tlMasterXbar ( // @[BaseTile.scala 195:42]
    .clock(tlMasterXbar_clock),
    .reset(tlMasterXbar_reset),
    .auto_in_1_a_ready(tlMasterXbar_auto_in_1_a_ready),
    .auto_in_1_a_valid(tlMasterXbar_auto_in_1_a_valid),
    .auto_in_1_a_bits_address(tlMasterXbar_auto_in_1_a_bits_address),
    .auto_in_1_d_valid(tlMasterXbar_auto_in_1_d_valid),
    .auto_in_1_d_bits_opcode(tlMasterXbar_auto_in_1_d_bits_opcode),
    .auto_in_1_d_bits_size(tlMasterXbar_auto_in_1_d_bits_size),
    .auto_in_1_d_bits_data(tlMasterXbar_auto_in_1_d_bits_data),
    .auto_in_1_d_bits_corrupt(tlMasterXbar_auto_in_1_d_bits_corrupt),
    .auto_in_0_a_ready(tlMasterXbar_auto_in_0_a_ready),
    .auto_in_0_a_valid(tlMasterXbar_auto_in_0_a_valid),
    .auto_in_0_a_bits_opcode(tlMasterXbar_auto_in_0_a_bits_opcode),
    .auto_in_0_a_bits_param(tlMasterXbar_auto_in_0_a_bits_param),
    .auto_in_0_a_bits_size(tlMasterXbar_auto_in_0_a_bits_size),
    .auto_in_0_a_bits_source(tlMasterXbar_auto_in_0_a_bits_source),
    .auto_in_0_a_bits_address(tlMasterXbar_auto_in_0_a_bits_address),
    .auto_in_0_a_bits_mask(tlMasterXbar_auto_in_0_a_bits_mask),
    .auto_in_0_a_bits_data(tlMasterXbar_auto_in_0_a_bits_data),
    .auto_in_0_b_ready(tlMasterXbar_auto_in_0_b_ready),
    .auto_in_0_b_valid(tlMasterXbar_auto_in_0_b_valid),
    .auto_in_0_b_bits_param(tlMasterXbar_auto_in_0_b_bits_param),
    .auto_in_0_b_bits_size(tlMasterXbar_auto_in_0_b_bits_size),
    .auto_in_0_b_bits_source(tlMasterXbar_auto_in_0_b_bits_source),
    .auto_in_0_b_bits_address(tlMasterXbar_auto_in_0_b_bits_address),
    .auto_in_0_c_ready(tlMasterXbar_auto_in_0_c_ready),
    .auto_in_0_c_valid(tlMasterXbar_auto_in_0_c_valid),
    .auto_in_0_c_bits_opcode(tlMasterXbar_auto_in_0_c_bits_opcode),
    .auto_in_0_c_bits_param(tlMasterXbar_auto_in_0_c_bits_param),
    .auto_in_0_c_bits_size(tlMasterXbar_auto_in_0_c_bits_size),
    .auto_in_0_c_bits_source(tlMasterXbar_auto_in_0_c_bits_source),
    .auto_in_0_c_bits_address(tlMasterXbar_auto_in_0_c_bits_address),
    .auto_in_0_c_bits_data(tlMasterXbar_auto_in_0_c_bits_data),
    .auto_in_0_d_ready(tlMasterXbar_auto_in_0_d_ready),
    .auto_in_0_d_valid(tlMasterXbar_auto_in_0_d_valid),
    .auto_in_0_d_bits_opcode(tlMasterXbar_auto_in_0_d_bits_opcode),
    .auto_in_0_d_bits_param(tlMasterXbar_auto_in_0_d_bits_param),
    .auto_in_0_d_bits_size(tlMasterXbar_auto_in_0_d_bits_size),
    .auto_in_0_d_bits_source(tlMasterXbar_auto_in_0_d_bits_source),
    .auto_in_0_d_bits_sink(tlMasterXbar_auto_in_0_d_bits_sink),
    .auto_in_0_d_bits_denied(tlMasterXbar_auto_in_0_d_bits_denied),
    .auto_in_0_d_bits_data(tlMasterXbar_auto_in_0_d_bits_data),
    .auto_in_0_e_ready(tlMasterXbar_auto_in_0_e_ready),
    .auto_in_0_e_valid(tlMasterXbar_auto_in_0_e_valid),
    .auto_in_0_e_bits_sink(tlMasterXbar_auto_in_0_e_bits_sink),
    .auto_out_a_ready(tlMasterXbar_auto_out_a_ready),
    .auto_out_a_valid(tlMasterXbar_auto_out_a_valid),
    .auto_out_a_bits_opcode(tlMasterXbar_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(tlMasterXbar_auto_out_a_bits_param),
    .auto_out_a_bits_size(tlMasterXbar_auto_out_a_bits_size),
    .auto_out_a_bits_source(tlMasterXbar_auto_out_a_bits_source),
    .auto_out_a_bits_address(tlMasterXbar_auto_out_a_bits_address),
    .auto_out_a_bits_mask(tlMasterXbar_auto_out_a_bits_mask),
    .auto_out_a_bits_data(tlMasterXbar_auto_out_a_bits_data),
    .auto_out_b_ready(tlMasterXbar_auto_out_b_ready),
    .auto_out_b_valid(tlMasterXbar_auto_out_b_valid),
    .auto_out_b_bits_opcode(tlMasterXbar_auto_out_b_bits_opcode),
    .auto_out_b_bits_param(tlMasterXbar_auto_out_b_bits_param),
    .auto_out_b_bits_size(tlMasterXbar_auto_out_b_bits_size),
    .auto_out_b_bits_source(tlMasterXbar_auto_out_b_bits_source),
    .auto_out_b_bits_address(tlMasterXbar_auto_out_b_bits_address),
    .auto_out_b_bits_mask(tlMasterXbar_auto_out_b_bits_mask),
    .auto_out_b_bits_corrupt(tlMasterXbar_auto_out_b_bits_corrupt),
    .auto_out_c_ready(tlMasterXbar_auto_out_c_ready),
    .auto_out_c_valid(tlMasterXbar_auto_out_c_valid),
    .auto_out_c_bits_opcode(tlMasterXbar_auto_out_c_bits_opcode),
    .auto_out_c_bits_param(tlMasterXbar_auto_out_c_bits_param),
    .auto_out_c_bits_size(tlMasterXbar_auto_out_c_bits_size),
    .auto_out_c_bits_source(tlMasterXbar_auto_out_c_bits_source),
    .auto_out_c_bits_address(tlMasterXbar_auto_out_c_bits_address),
    .auto_out_c_bits_data(tlMasterXbar_auto_out_c_bits_data),
    .auto_out_d_ready(tlMasterXbar_auto_out_d_ready),
    .auto_out_d_valid(tlMasterXbar_auto_out_d_valid),
    .auto_out_d_bits_opcode(tlMasterXbar_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(tlMasterXbar_auto_out_d_bits_param),
    .auto_out_d_bits_size(tlMasterXbar_auto_out_d_bits_size),
    .auto_out_d_bits_source(tlMasterXbar_auto_out_d_bits_source),
    .auto_out_d_bits_sink(tlMasterXbar_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(tlMasterXbar_auto_out_d_bits_denied),
    .auto_out_d_bits_data(tlMasterXbar_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(tlMasterXbar_auto_out_d_bits_corrupt),
    .auto_out_e_ready(tlMasterXbar_auto_out_e_ready),
    .auto_out_e_valid(tlMasterXbar_auto_out_e_valid),
    .auto_out_e_bits_sink(tlMasterXbar_auto_out_e_bits_sink),
    .io_covSum(tlMasterXbar_io_covSum),
    .metaAssert(tlMasterXbar_metaAssert),
    .metaReset(tlMasterXbar_metaReset),
    .monitor_halt(tlMasterXbar_monitor_halt),
    .monitor_1_halt(tlMasterXbar_monitor_1_halt)
  );
  IntXbar_1 intXbar ( // @[BaseTile.scala 197:37]
    .auto_int_in_3_0(intXbar_auto_int_in_3_0),
    .auto_int_in_2_0(intXbar_auto_int_in_2_0),
    .auto_int_in_1_0(intXbar_auto_int_in_1_0),
    .auto_int_in_1_1(intXbar_auto_int_in_1_1),
    .auto_int_in_0_0(intXbar_auto_int_in_0_0),
    .auto_int_out_0(intXbar_auto_int_out_0),
    .auto_int_out_1(intXbar_auto_int_out_1),
    .auto_int_out_2(intXbar_auto_int_out_2),
    .auto_int_out_3(intXbar_auto_int_out_3),
    .auto_int_out_4(intXbar_auto_int_out_4),
    .io_covSum(intXbar_io_covSum),
    .metaAssert(intXbar_metaAssert)
  );
  BundleBridgeNexus_6 broadcast ( // @[BundleBridge.scala 196:31]
    .auto_in(broadcast_auto_in),
    .auto_out(broadcast_auto_out),
    .io_covSum(broadcast_io_covSum),
    .metaAssert(broadcast_metaAssert)
  );
  BundleBridgeNexus_7 broadcast_1 ( // @[BundleBridge.scala 196:31]
    .auto_in(broadcast_1_auto_in),
    .auto_out_1(broadcast_1_auto_out_1),
    .io_covSum(broadcast_1_io_covSum),
    .metaAssert(broadcast_1_metaAssert)
  );
  BundleBridgeNexus_10 broadcast_3 ( // @[BundleBridge.scala 196:31]
    .auto_in_0_valid(broadcast_3_auto_in_0_valid),
    .auto_in_0_iaddr(broadcast_3_auto_in_0_iaddr),
    .auto_in_0_insn(broadcast_3_auto_in_0_insn),
    .auto_in_0_priv(broadcast_3_auto_in_0_priv),
    .auto_in_0_exception(broadcast_3_auto_in_0_exception),
    .auto_in_0_interrupt(broadcast_3_auto_in_0_interrupt),
    .auto_in_0_cause(broadcast_3_auto_in_0_cause),
    .auto_in_0_tval(broadcast_3_auto_in_0_tval),
    .auto_out_0_valid(broadcast_3_auto_out_0_valid),
    .auto_out_0_iaddr(broadcast_3_auto_out_0_iaddr),
    .auto_out_0_insn(broadcast_3_auto_out_0_insn),
    .auto_out_0_priv(broadcast_3_auto_out_0_priv),
    .auto_out_0_exception(broadcast_3_auto_out_0_exception),
    .auto_out_0_interrupt(broadcast_3_auto_out_0_interrupt),
    .auto_out_0_cause(broadcast_3_auto_out_0_cause),
    .auto_out_0_tval(broadcast_3_auto_out_0_tval),
    .io_covSum(broadcast_3_io_covSum),
    .metaAssert(broadcast_3_metaAssert)
  );
  DCache dcache ( // @[HellaCache.scala 265:43]
    .gated_clock(dcache_gated_clock),
    .reset(dcache_reset),
    .auto_out_a_ready(dcache_auto_out_a_ready),
    .auto_out_a_valid(dcache_auto_out_a_valid),
    .auto_out_a_bits_opcode(dcache_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(dcache_auto_out_a_bits_param),
    .auto_out_a_bits_size(dcache_auto_out_a_bits_size),
    .auto_out_a_bits_source(dcache_auto_out_a_bits_source),
    .auto_out_a_bits_address(dcache_auto_out_a_bits_address),
    .auto_out_a_bits_mask(dcache_auto_out_a_bits_mask),
    .auto_out_a_bits_data(dcache_auto_out_a_bits_data),
    .auto_out_b_ready(dcache_auto_out_b_ready),
    .auto_out_b_valid(dcache_auto_out_b_valid),
    .auto_out_b_bits_param(dcache_auto_out_b_bits_param),
    .auto_out_b_bits_size(dcache_auto_out_b_bits_size),
    .auto_out_b_bits_source(dcache_auto_out_b_bits_source),
    .auto_out_b_bits_address(dcache_auto_out_b_bits_address),
    .auto_out_c_ready(dcache_auto_out_c_ready),
    .auto_out_c_valid(dcache_auto_out_c_valid),
    .auto_out_c_bits_opcode(dcache_auto_out_c_bits_opcode),
    .auto_out_c_bits_param(dcache_auto_out_c_bits_param),
    .auto_out_c_bits_size(dcache_auto_out_c_bits_size),
    .auto_out_c_bits_source(dcache_auto_out_c_bits_source),
    .auto_out_c_bits_address(dcache_auto_out_c_bits_address),
    .auto_out_c_bits_data(dcache_auto_out_c_bits_data),
    .auto_out_d_ready(dcache_auto_out_d_ready),
    .auto_out_d_valid(dcache_auto_out_d_valid),
    .auto_out_d_bits_opcode(dcache_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(dcache_auto_out_d_bits_param),
    .auto_out_d_bits_size(dcache_auto_out_d_bits_size),
    .auto_out_d_bits_source(dcache_auto_out_d_bits_source),
    .auto_out_d_bits_sink(dcache_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(dcache_auto_out_d_bits_denied),
    .auto_out_d_bits_data(dcache_auto_out_d_bits_data),
    .auto_out_e_ready(dcache_auto_out_e_ready),
    .auto_out_e_valid(dcache_auto_out_e_valid),
    .auto_out_e_bits_sink(dcache_auto_out_e_bits_sink),
    .io_cpu_req_ready(dcache_io_cpu_req_ready),
    .io_cpu_req_valid(dcache_io_cpu_req_valid),
    .io_cpu_req_bits_addr(dcache_io_cpu_req_bits_addr),
    .io_cpu_req_bits_tag(dcache_io_cpu_req_bits_tag),
    .io_cpu_req_bits_cmd(dcache_io_cpu_req_bits_cmd),
    .io_cpu_req_bits_size(dcache_io_cpu_req_bits_size),
    .io_cpu_req_bits_signed(dcache_io_cpu_req_bits_signed),
    .io_cpu_req_bits_phys(dcache_io_cpu_req_bits_phys),
    .io_cpu_s1_kill(dcache_io_cpu_s1_kill),
    .io_cpu_s1_data_data(dcache_io_cpu_s1_data_data),
    .io_cpu_s2_nack(dcache_io_cpu_s2_nack),
    .io_cpu_resp_valid(dcache_io_cpu_resp_valid),
    .io_cpu_resp_bits_tag(dcache_io_cpu_resp_bits_tag),
    .io_cpu_resp_bits_size(dcache_io_cpu_resp_bits_size),
    .io_cpu_resp_bits_data(dcache_io_cpu_resp_bits_data),
    .io_cpu_resp_bits_replay(dcache_io_cpu_resp_bits_replay),
    .io_cpu_resp_bits_has_data(dcache_io_cpu_resp_bits_has_data),
    .io_cpu_resp_bits_data_word_bypass(dcache_io_cpu_resp_bits_data_word_bypass),
    .io_cpu_replay_next(dcache_io_cpu_replay_next),
    .io_cpu_s2_xcpt_ma_ld(dcache_io_cpu_s2_xcpt_ma_ld),
    .io_cpu_s2_xcpt_ma_st(dcache_io_cpu_s2_xcpt_ma_st),
    .io_cpu_s2_xcpt_pf_ld(dcache_io_cpu_s2_xcpt_pf_ld),
    .io_cpu_s2_xcpt_pf_st(dcache_io_cpu_s2_xcpt_pf_st),
    .io_cpu_s2_xcpt_ae_ld(dcache_io_cpu_s2_xcpt_ae_ld),
    .io_cpu_s2_xcpt_ae_st(dcache_io_cpu_s2_xcpt_ae_st),
    .io_cpu_ordered(dcache_io_cpu_ordered),
    .io_cpu_perf_release(dcache_io_cpu_perf_release),
    .io_cpu_perf_grant(dcache_io_cpu_perf_grant),
    .io_ptw_req_ready(dcache_io_ptw_req_ready),
    .io_ptw_req_valid(dcache_io_ptw_req_valid),
    .io_ptw_req_bits_bits_addr(dcache_io_ptw_req_bits_bits_addr),
    .io_ptw_resp_valid(dcache_io_ptw_resp_valid),
    .io_ptw_resp_bits_ae(dcache_io_ptw_resp_bits_ae),
    .io_ptw_resp_bits_pte_ppn(dcache_io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_d(dcache_io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_a(dcache_io_ptw_resp_bits_pte_a),
    .io_ptw_resp_bits_pte_g(dcache_io_ptw_resp_bits_pte_g),
    .io_ptw_resp_bits_pte_u(dcache_io_ptw_resp_bits_pte_u),
    .io_ptw_resp_bits_pte_x(dcache_io_ptw_resp_bits_pte_x),
    .io_ptw_resp_bits_pte_w(dcache_io_ptw_resp_bits_pte_w),
    .io_ptw_resp_bits_pte_r(dcache_io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_v(dcache_io_ptw_resp_bits_pte_v),
    .io_ptw_resp_bits_level(dcache_io_ptw_resp_bits_level),
    .io_ptw_resp_bits_homogeneous(dcache_io_ptw_resp_bits_homogeneous),
    .io_ptw_ptbr_mode(dcache_io_ptw_ptbr_mode),
    .io_ptw_status_debug(dcache_io_ptw_status_debug),
    .io_ptw_status_dprv(dcache_io_ptw_status_dprv),
    .io_ptw_status_mxr(dcache_io_ptw_status_mxr),
    .io_ptw_status_sum(dcache_io_ptw_status_sum),
    .io_ptw_pmp_0_cfg_l(dcache_io_ptw_pmp_0_cfg_l),
    .io_ptw_pmp_0_cfg_a(dcache_io_ptw_pmp_0_cfg_a),
    .io_ptw_pmp_0_cfg_x(dcache_io_ptw_pmp_0_cfg_x),
    .io_ptw_pmp_0_cfg_w(dcache_io_ptw_pmp_0_cfg_w),
    .io_ptw_pmp_0_cfg_r(dcache_io_ptw_pmp_0_cfg_r),
    .io_ptw_pmp_0_addr(dcache_io_ptw_pmp_0_addr),
    .io_ptw_pmp_0_mask(dcache_io_ptw_pmp_0_mask),
    .io_ptw_pmp_1_cfg_l(dcache_io_ptw_pmp_1_cfg_l),
    .io_ptw_pmp_1_cfg_a(dcache_io_ptw_pmp_1_cfg_a),
    .io_ptw_pmp_1_cfg_x(dcache_io_ptw_pmp_1_cfg_x),
    .io_ptw_pmp_1_cfg_w(dcache_io_ptw_pmp_1_cfg_w),
    .io_ptw_pmp_1_cfg_r(dcache_io_ptw_pmp_1_cfg_r),
    .io_ptw_pmp_1_addr(dcache_io_ptw_pmp_1_addr),
    .io_ptw_pmp_1_mask(dcache_io_ptw_pmp_1_mask),
    .io_ptw_pmp_2_cfg_l(dcache_io_ptw_pmp_2_cfg_l),
    .io_ptw_pmp_2_cfg_a(dcache_io_ptw_pmp_2_cfg_a),
    .io_ptw_pmp_2_cfg_x(dcache_io_ptw_pmp_2_cfg_x),
    .io_ptw_pmp_2_cfg_w(dcache_io_ptw_pmp_2_cfg_w),
    .io_ptw_pmp_2_cfg_r(dcache_io_ptw_pmp_2_cfg_r),
    .io_ptw_pmp_2_addr(dcache_io_ptw_pmp_2_addr),
    .io_ptw_pmp_2_mask(dcache_io_ptw_pmp_2_mask),
    .io_ptw_pmp_3_cfg_l(dcache_io_ptw_pmp_3_cfg_l),
    .io_ptw_pmp_3_cfg_a(dcache_io_ptw_pmp_3_cfg_a),
    .io_ptw_pmp_3_cfg_x(dcache_io_ptw_pmp_3_cfg_x),
    .io_ptw_pmp_3_cfg_w(dcache_io_ptw_pmp_3_cfg_w),
    .io_ptw_pmp_3_cfg_r(dcache_io_ptw_pmp_3_cfg_r),
    .io_ptw_pmp_3_addr(dcache_io_ptw_pmp_3_addr),
    .io_ptw_pmp_3_mask(dcache_io_ptw_pmp_3_mask),
    .io_ptw_pmp_4_cfg_l(dcache_io_ptw_pmp_4_cfg_l),
    .io_ptw_pmp_4_cfg_a(dcache_io_ptw_pmp_4_cfg_a),
    .io_ptw_pmp_4_cfg_x(dcache_io_ptw_pmp_4_cfg_x),
    .io_ptw_pmp_4_cfg_w(dcache_io_ptw_pmp_4_cfg_w),
    .io_ptw_pmp_4_cfg_r(dcache_io_ptw_pmp_4_cfg_r),
    .io_ptw_pmp_4_addr(dcache_io_ptw_pmp_4_addr),
    .io_ptw_pmp_4_mask(dcache_io_ptw_pmp_4_mask),
    .io_ptw_pmp_5_cfg_l(dcache_io_ptw_pmp_5_cfg_l),
    .io_ptw_pmp_5_cfg_a(dcache_io_ptw_pmp_5_cfg_a),
    .io_ptw_pmp_5_cfg_x(dcache_io_ptw_pmp_5_cfg_x),
    .io_ptw_pmp_5_cfg_w(dcache_io_ptw_pmp_5_cfg_w),
    .io_ptw_pmp_5_cfg_r(dcache_io_ptw_pmp_5_cfg_r),
    .io_ptw_pmp_5_addr(dcache_io_ptw_pmp_5_addr),
    .io_ptw_pmp_5_mask(dcache_io_ptw_pmp_5_mask),
    .io_ptw_pmp_6_cfg_l(dcache_io_ptw_pmp_6_cfg_l),
    .io_ptw_pmp_6_cfg_a(dcache_io_ptw_pmp_6_cfg_a),
    .io_ptw_pmp_6_cfg_x(dcache_io_ptw_pmp_6_cfg_x),
    .io_ptw_pmp_6_cfg_w(dcache_io_ptw_pmp_6_cfg_w),
    .io_ptw_pmp_6_cfg_r(dcache_io_ptw_pmp_6_cfg_r),
    .io_ptw_pmp_6_addr(dcache_io_ptw_pmp_6_addr),
    .io_ptw_pmp_6_mask(dcache_io_ptw_pmp_6_mask),
    .io_ptw_pmp_7_cfg_l(dcache_io_ptw_pmp_7_cfg_l),
    .io_ptw_pmp_7_cfg_a(dcache_io_ptw_pmp_7_cfg_a),
    .io_ptw_pmp_7_cfg_x(dcache_io_ptw_pmp_7_cfg_x),
    .io_ptw_pmp_7_cfg_w(dcache_io_ptw_pmp_7_cfg_w),
    .io_ptw_pmp_7_cfg_r(dcache_io_ptw_pmp_7_cfg_r),
    .io_ptw_pmp_7_addr(dcache_io_ptw_pmp_7_addr),
    .io_ptw_pmp_7_mask(dcache_io_ptw_pmp_7_mask),
    .io_covSum(dcache_io_covSum),
    .metaAssert(dcache_metaAssert),
    .metaReset(dcache_metaReset),
    .data_halt(dcache_data_halt),
    .tlb_halt(dcache_tlb_halt),
    .pma_checker_halt(dcache_pma_checker_halt),
    .lfsr_prng_halt(dcache_lfsr_prng_halt)
  );
  Frontend frontend ( // @[Frontend.scala 350:28]
    .gated_clock(frontend_gated_clock),
    .reset(frontend_reset),
    .auto_icache_master_out_a_ready(frontend_auto_icache_master_out_a_ready),
    .auto_icache_master_out_a_valid(frontend_auto_icache_master_out_a_valid),
    .auto_icache_master_out_a_bits_address(frontend_auto_icache_master_out_a_bits_address),
    .auto_icache_master_out_d_valid(frontend_auto_icache_master_out_d_valid),
    .auto_icache_master_out_d_bits_opcode(frontend_auto_icache_master_out_d_bits_opcode),
    .auto_icache_master_out_d_bits_size(frontend_auto_icache_master_out_d_bits_size),
    .auto_icache_master_out_d_bits_data(frontend_auto_icache_master_out_d_bits_data),
    .auto_icache_master_out_d_bits_corrupt(frontend_auto_icache_master_out_d_bits_corrupt),
    .auto_reset_vector_sink_in(frontend_auto_reset_vector_sink_in),
    .io_cpu_might_request(frontend_io_cpu_might_request),
    .io_cpu_req_valid(frontend_io_cpu_req_valid),
    .io_cpu_req_bits_pc(frontend_io_cpu_req_bits_pc),
    .io_cpu_req_bits_speculative(frontend_io_cpu_req_bits_speculative),
    .io_cpu_sfence_valid(frontend_io_cpu_sfence_valid),
    .io_cpu_sfence_bits_rs1(frontend_io_cpu_sfence_bits_rs1),
    .io_cpu_sfence_bits_rs2(frontend_io_cpu_sfence_bits_rs2),
    .io_cpu_sfence_bits_addr(frontend_io_cpu_sfence_bits_addr),
    .io_cpu_resp_ready(frontend_io_cpu_resp_ready),
    .io_cpu_resp_valid(frontend_io_cpu_resp_valid),
    .io_cpu_resp_bits_btb_taken(frontend_io_cpu_resp_bits_btb_taken),
    .io_cpu_resp_bits_btb_bridx(frontend_io_cpu_resp_bits_btb_bridx),
    .io_cpu_resp_bits_btb_entry(frontend_io_cpu_resp_bits_btb_entry),
    .io_cpu_resp_bits_btb_bht_history(frontend_io_cpu_resp_bits_btb_bht_history),
    .io_cpu_resp_bits_pc(frontend_io_cpu_resp_bits_pc),
    .io_cpu_resp_bits_data(frontend_io_cpu_resp_bits_data),
    .io_cpu_resp_bits_xcpt_pf_inst(frontend_io_cpu_resp_bits_xcpt_pf_inst),
    .io_cpu_resp_bits_xcpt_ae_inst(frontend_io_cpu_resp_bits_xcpt_ae_inst),
    .io_cpu_resp_bits_replay(frontend_io_cpu_resp_bits_replay),
    .io_cpu_btb_update_valid(frontend_io_cpu_btb_update_valid),
    .io_cpu_btb_update_bits_prediction_entry(frontend_io_cpu_btb_update_bits_prediction_entry),
    .io_cpu_btb_update_bits_pc(frontend_io_cpu_btb_update_bits_pc),
    .io_cpu_btb_update_bits_isValid(frontend_io_cpu_btb_update_bits_isValid),
    .io_cpu_btb_update_bits_br_pc(frontend_io_cpu_btb_update_bits_br_pc),
    .io_cpu_btb_update_bits_cfiType(frontend_io_cpu_btb_update_bits_cfiType),
    .io_cpu_bht_update_valid(frontend_io_cpu_bht_update_valid),
    .io_cpu_bht_update_bits_prediction_history(frontend_io_cpu_bht_update_bits_prediction_history),
    .io_cpu_bht_update_bits_pc(frontend_io_cpu_bht_update_bits_pc),
    .io_cpu_bht_update_bits_branch(frontend_io_cpu_bht_update_bits_branch),
    .io_cpu_bht_update_bits_taken(frontend_io_cpu_bht_update_bits_taken),
    .io_cpu_bht_update_bits_mispredict(frontend_io_cpu_bht_update_bits_mispredict),
    .io_cpu_flush_icache(frontend_io_cpu_flush_icache),
    .io_cpu_npc(frontend_io_cpu_npc),
    .io_ptw_req_ready(frontend_io_ptw_req_ready),
    .io_ptw_req_valid(frontend_io_ptw_req_valid),
    .io_ptw_req_bits_valid(frontend_io_ptw_req_bits_valid),
    .io_ptw_req_bits_bits_addr(frontend_io_ptw_req_bits_bits_addr),
    .io_ptw_resp_valid(frontend_io_ptw_resp_valid),
    .io_ptw_resp_bits_ae(frontend_io_ptw_resp_bits_ae),
    .io_ptw_resp_bits_pte_ppn(frontend_io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_d(frontend_io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_a(frontend_io_ptw_resp_bits_pte_a),
    .io_ptw_resp_bits_pte_g(frontend_io_ptw_resp_bits_pte_g),
    .io_ptw_resp_bits_pte_u(frontend_io_ptw_resp_bits_pte_u),
    .io_ptw_resp_bits_pte_x(frontend_io_ptw_resp_bits_pte_x),
    .io_ptw_resp_bits_pte_w(frontend_io_ptw_resp_bits_pte_w),
    .io_ptw_resp_bits_pte_r(frontend_io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_v(frontend_io_ptw_resp_bits_pte_v),
    .io_ptw_resp_bits_level(frontend_io_ptw_resp_bits_level),
    .io_ptw_resp_bits_homogeneous(frontend_io_ptw_resp_bits_homogeneous),
    .io_ptw_ptbr_mode(frontend_io_ptw_ptbr_mode),
    .io_ptw_status_debug(frontend_io_ptw_status_debug),
    .io_ptw_status_prv(frontend_io_ptw_status_prv),
    .io_ptw_pmp_0_cfg_l(frontend_io_ptw_pmp_0_cfg_l),
    .io_ptw_pmp_0_cfg_a(frontend_io_ptw_pmp_0_cfg_a),
    .io_ptw_pmp_0_cfg_x(frontend_io_ptw_pmp_0_cfg_x),
    .io_ptw_pmp_0_cfg_w(frontend_io_ptw_pmp_0_cfg_w),
    .io_ptw_pmp_0_cfg_r(frontend_io_ptw_pmp_0_cfg_r),
    .io_ptw_pmp_0_addr(frontend_io_ptw_pmp_0_addr),
    .io_ptw_pmp_0_mask(frontend_io_ptw_pmp_0_mask),
    .io_ptw_pmp_1_cfg_l(frontend_io_ptw_pmp_1_cfg_l),
    .io_ptw_pmp_1_cfg_a(frontend_io_ptw_pmp_1_cfg_a),
    .io_ptw_pmp_1_cfg_x(frontend_io_ptw_pmp_1_cfg_x),
    .io_ptw_pmp_1_cfg_w(frontend_io_ptw_pmp_1_cfg_w),
    .io_ptw_pmp_1_cfg_r(frontend_io_ptw_pmp_1_cfg_r),
    .io_ptw_pmp_1_addr(frontend_io_ptw_pmp_1_addr),
    .io_ptw_pmp_1_mask(frontend_io_ptw_pmp_1_mask),
    .io_ptw_pmp_2_cfg_l(frontend_io_ptw_pmp_2_cfg_l),
    .io_ptw_pmp_2_cfg_a(frontend_io_ptw_pmp_2_cfg_a),
    .io_ptw_pmp_2_cfg_x(frontend_io_ptw_pmp_2_cfg_x),
    .io_ptw_pmp_2_cfg_w(frontend_io_ptw_pmp_2_cfg_w),
    .io_ptw_pmp_2_cfg_r(frontend_io_ptw_pmp_2_cfg_r),
    .io_ptw_pmp_2_addr(frontend_io_ptw_pmp_2_addr),
    .io_ptw_pmp_2_mask(frontend_io_ptw_pmp_2_mask),
    .io_ptw_pmp_3_cfg_l(frontend_io_ptw_pmp_3_cfg_l),
    .io_ptw_pmp_3_cfg_a(frontend_io_ptw_pmp_3_cfg_a),
    .io_ptw_pmp_3_cfg_x(frontend_io_ptw_pmp_3_cfg_x),
    .io_ptw_pmp_3_cfg_w(frontend_io_ptw_pmp_3_cfg_w),
    .io_ptw_pmp_3_cfg_r(frontend_io_ptw_pmp_3_cfg_r),
    .io_ptw_pmp_3_addr(frontend_io_ptw_pmp_3_addr),
    .io_ptw_pmp_3_mask(frontend_io_ptw_pmp_3_mask),
    .io_ptw_pmp_4_cfg_l(frontend_io_ptw_pmp_4_cfg_l),
    .io_ptw_pmp_4_cfg_a(frontend_io_ptw_pmp_4_cfg_a),
    .io_ptw_pmp_4_cfg_x(frontend_io_ptw_pmp_4_cfg_x),
    .io_ptw_pmp_4_cfg_w(frontend_io_ptw_pmp_4_cfg_w),
    .io_ptw_pmp_4_cfg_r(frontend_io_ptw_pmp_4_cfg_r),
    .io_ptw_pmp_4_addr(frontend_io_ptw_pmp_4_addr),
    .io_ptw_pmp_4_mask(frontend_io_ptw_pmp_4_mask),
    .io_ptw_pmp_5_cfg_l(frontend_io_ptw_pmp_5_cfg_l),
    .io_ptw_pmp_5_cfg_a(frontend_io_ptw_pmp_5_cfg_a),
    .io_ptw_pmp_5_cfg_x(frontend_io_ptw_pmp_5_cfg_x),
    .io_ptw_pmp_5_cfg_w(frontend_io_ptw_pmp_5_cfg_w),
    .io_ptw_pmp_5_cfg_r(frontend_io_ptw_pmp_5_cfg_r),
    .io_ptw_pmp_5_addr(frontend_io_ptw_pmp_5_addr),
    .io_ptw_pmp_5_mask(frontend_io_ptw_pmp_5_mask),
    .io_ptw_pmp_6_cfg_l(frontend_io_ptw_pmp_6_cfg_l),
    .io_ptw_pmp_6_cfg_a(frontend_io_ptw_pmp_6_cfg_a),
    .io_ptw_pmp_6_cfg_x(frontend_io_ptw_pmp_6_cfg_x),
    .io_ptw_pmp_6_cfg_w(frontend_io_ptw_pmp_6_cfg_w),
    .io_ptw_pmp_6_cfg_r(frontend_io_ptw_pmp_6_cfg_r),
    .io_ptw_pmp_6_addr(frontend_io_ptw_pmp_6_addr),
    .io_ptw_pmp_6_mask(frontend_io_ptw_pmp_6_mask),
    .io_ptw_pmp_7_cfg_l(frontend_io_ptw_pmp_7_cfg_l),
    .io_ptw_pmp_7_cfg_a(frontend_io_ptw_pmp_7_cfg_a),
    .io_ptw_pmp_7_cfg_x(frontend_io_ptw_pmp_7_cfg_x),
    .io_ptw_pmp_7_cfg_w(frontend_io_ptw_pmp_7_cfg_w),
    .io_ptw_pmp_7_cfg_r(frontend_io_ptw_pmp_7_cfg_r),
    .io_ptw_pmp_7_addr(frontend_io_ptw_pmp_7_addr),
    .io_ptw_pmp_7_mask(frontend_io_ptw_pmp_7_mask),
    .io_ptw_customCSRs_csrs_0_value(frontend_io_ptw_customCSRs_csrs_0_value),
    .io_covSum(frontend_io_covSum),
    .metaAssert(frontend_metaAssert),
    .metaReset(frontend_metaReset),
    .icache_halt(frontend_icache_halt),
    .fq_halt(frontend_fq_halt),
    .tlb_halt(frontend_tlb_halt),
    .btb_halt(frontend_btb_halt)
  );
  FPU fpuOpt ( // @[RocketTile.scala 202:62]
    .clock(fpuOpt_clock),
    .reset(fpuOpt_reset),
    .io_inst(fpuOpt_io_inst),
    .io_fromint_data(fpuOpt_io_fromint_data),
    .io_fcsr_rm(fpuOpt_io_fcsr_rm),
    .io_fcsr_flags_valid(fpuOpt_io_fcsr_flags_valid),
    .io_fcsr_flags_bits(fpuOpt_io_fcsr_flags_bits),
    .io_store_data(fpuOpt_io_store_data),
    .io_toint_data(fpuOpt_io_toint_data),
    .io_dmem_resp_val(fpuOpt_io_dmem_resp_val),
    .io_dmem_resp_type(fpuOpt_io_dmem_resp_type),
    .io_dmem_resp_tag(fpuOpt_io_dmem_resp_tag),
    .io_dmem_resp_data(fpuOpt_io_dmem_resp_data),
    .io_valid(fpuOpt_io_valid),
    .io_fcsr_rdy(fpuOpt_io_fcsr_rdy),
    .io_nack_mem(fpuOpt_io_nack_mem),
    .io_illegal_rm(fpuOpt_io_illegal_rm),
    .io_killx(fpuOpt_io_killx),
    .io_killm(fpuOpt_io_killm),
    .io_dec_wen(fpuOpt_io_dec_wen),
    .io_dec_ren1(fpuOpt_io_dec_ren1),
    .io_dec_ren2(fpuOpt_io_dec_ren2),
    .io_dec_ren3(fpuOpt_io_dec_ren3),
    .io_sboard_set(fpuOpt_io_sboard_set),
    .io_sboard_clr(fpuOpt_io_sboard_clr),
    .io_sboard_clra(fpuOpt_io_sboard_clra),
    .io_covSum(fpuOpt_io_covSum),
    .metaAssert(fpuOpt_metaAssert),
    .metaReset(fpuOpt_metaReset),
    .fpiu_halt(fpuOpt_fpiu_halt),
    .ifpu_halt(fpuOpt_ifpu_halt),
    .sfma_halt(fpuOpt_sfma_halt),
    .fpmu_halt(fpuOpt_fpmu_halt),
    .divSqrt_1_halt(fpuOpt_divSqrt_1_halt),
    .dfma_halt(fpuOpt_dfma_halt),
    .divSqrt_halt(fpuOpt_divSqrt_halt)
  );
  HellaCacheArbiter dcacheArb ( // @[HellaCache.scala 276:25]
    .clock(dcacheArb_clock),
    .io_requestor_0_req_ready(dcacheArb_io_requestor_0_req_ready),
    .io_requestor_0_req_valid(dcacheArb_io_requestor_0_req_valid),
    .io_requestor_0_req_bits_addr(dcacheArb_io_requestor_0_req_bits_addr),
    .io_requestor_0_s1_kill(dcacheArb_io_requestor_0_s1_kill),
    .io_requestor_0_s2_nack(dcacheArb_io_requestor_0_s2_nack),
    .io_requestor_0_resp_valid(dcacheArb_io_requestor_0_resp_valid),
    .io_requestor_0_resp_bits_data(dcacheArb_io_requestor_0_resp_bits_data),
    .io_requestor_0_s2_xcpt_ae_ld(dcacheArb_io_requestor_0_s2_xcpt_ae_ld),
    .io_requestor_1_req_ready(dcacheArb_io_requestor_1_req_ready),
    .io_requestor_1_req_valid(dcacheArb_io_requestor_1_req_valid),
    .io_requestor_1_req_bits_addr(dcacheArb_io_requestor_1_req_bits_addr),
    .io_requestor_1_req_bits_tag(dcacheArb_io_requestor_1_req_bits_tag),
    .io_requestor_1_req_bits_cmd(dcacheArb_io_requestor_1_req_bits_cmd),
    .io_requestor_1_req_bits_size(dcacheArb_io_requestor_1_req_bits_size),
    .io_requestor_1_req_bits_signed(dcacheArb_io_requestor_1_req_bits_signed),
    .io_requestor_1_s1_kill(dcacheArb_io_requestor_1_s1_kill),
    .io_requestor_1_s1_data_data(dcacheArb_io_requestor_1_s1_data_data),
    .io_requestor_1_s2_nack(dcacheArb_io_requestor_1_s2_nack),
    .io_requestor_1_resp_valid(dcacheArb_io_requestor_1_resp_valid),
    .io_requestor_1_resp_bits_tag(dcacheArb_io_requestor_1_resp_bits_tag),
    .io_requestor_1_resp_bits_size(dcacheArb_io_requestor_1_resp_bits_size),
    .io_requestor_1_resp_bits_data(dcacheArb_io_requestor_1_resp_bits_data),
    .io_requestor_1_resp_bits_replay(dcacheArb_io_requestor_1_resp_bits_replay),
    .io_requestor_1_resp_bits_has_data(dcacheArb_io_requestor_1_resp_bits_has_data),
    .io_requestor_1_resp_bits_data_word_bypass(dcacheArb_io_requestor_1_resp_bits_data_word_bypass),
    .io_requestor_1_replay_next(dcacheArb_io_requestor_1_replay_next),
    .io_requestor_1_s2_xcpt_ma_ld(dcacheArb_io_requestor_1_s2_xcpt_ma_ld),
    .io_requestor_1_s2_xcpt_ma_st(dcacheArb_io_requestor_1_s2_xcpt_ma_st),
    .io_requestor_1_s2_xcpt_pf_ld(dcacheArb_io_requestor_1_s2_xcpt_pf_ld),
    .io_requestor_1_s2_xcpt_pf_st(dcacheArb_io_requestor_1_s2_xcpt_pf_st),
    .io_requestor_1_s2_xcpt_ae_ld(dcacheArb_io_requestor_1_s2_xcpt_ae_ld),
    .io_requestor_1_s2_xcpt_ae_st(dcacheArb_io_requestor_1_s2_xcpt_ae_st),
    .io_requestor_1_ordered(dcacheArb_io_requestor_1_ordered),
    .io_requestor_1_perf_release(dcacheArb_io_requestor_1_perf_release),
    .io_requestor_1_perf_grant(dcacheArb_io_requestor_1_perf_grant),
    .io_mem_req_ready(dcacheArb_io_mem_req_ready),
    .io_mem_req_valid(dcacheArb_io_mem_req_valid),
    .io_mem_req_bits_addr(dcacheArb_io_mem_req_bits_addr),
    .io_mem_req_bits_tag(dcacheArb_io_mem_req_bits_tag),
    .io_mem_req_bits_cmd(dcacheArb_io_mem_req_bits_cmd),
    .io_mem_req_bits_size(dcacheArb_io_mem_req_bits_size),
    .io_mem_req_bits_signed(dcacheArb_io_mem_req_bits_signed),
    .io_mem_req_bits_phys(dcacheArb_io_mem_req_bits_phys),
    .io_mem_s1_kill(dcacheArb_io_mem_s1_kill),
    .io_mem_s1_data_data(dcacheArb_io_mem_s1_data_data),
    .io_mem_s2_nack(dcacheArb_io_mem_s2_nack),
    .io_mem_resp_valid(dcacheArb_io_mem_resp_valid),
    .io_mem_resp_bits_tag(dcacheArb_io_mem_resp_bits_tag),
    .io_mem_resp_bits_size(dcacheArb_io_mem_resp_bits_size),
    .io_mem_resp_bits_data(dcacheArb_io_mem_resp_bits_data),
    .io_mem_resp_bits_replay(dcacheArb_io_mem_resp_bits_replay),
    .io_mem_resp_bits_has_data(dcacheArb_io_mem_resp_bits_has_data),
    .io_mem_resp_bits_data_word_bypass(dcacheArb_io_mem_resp_bits_data_word_bypass),
    .io_mem_replay_next(dcacheArb_io_mem_replay_next),
    .io_mem_s2_xcpt_ma_ld(dcacheArb_io_mem_s2_xcpt_ma_ld),
    .io_mem_s2_xcpt_ma_st(dcacheArb_io_mem_s2_xcpt_ma_st),
    .io_mem_s2_xcpt_pf_ld(dcacheArb_io_mem_s2_xcpt_pf_ld),
    .io_mem_s2_xcpt_pf_st(dcacheArb_io_mem_s2_xcpt_pf_st),
    .io_mem_s2_xcpt_ae_ld(dcacheArb_io_mem_s2_xcpt_ae_ld),
    .io_mem_s2_xcpt_ae_st(dcacheArb_io_mem_s2_xcpt_ae_st),
    .io_mem_ordered(dcacheArb_io_mem_ordered),
    .io_mem_perf_release(dcacheArb_io_mem_perf_release),
    .io_mem_perf_grant(dcacheArb_io_mem_perf_grant),
    .io_covSum(dcacheArb_io_covSum),
    .metaAssert(dcacheArb_metaAssert),
    .metaReset(dcacheArb_metaReset)
  );
  PTW ptw ( // @[PTW.scala 439:19]
    .clock(ptw_clock),
    .reset(ptw_reset),
    .io_requestor_0_req_ready(ptw_io_requestor_0_req_ready),
    .io_requestor_0_req_valid(ptw_io_requestor_0_req_valid),
    .io_requestor_0_req_bits_bits_addr(ptw_io_requestor_0_req_bits_bits_addr),
    .io_requestor_0_resp_valid(ptw_io_requestor_0_resp_valid),
    .io_requestor_0_resp_bits_ae(ptw_io_requestor_0_resp_bits_ae),
    .io_requestor_0_resp_bits_pte_ppn(ptw_io_requestor_0_resp_bits_pte_ppn),
    .io_requestor_0_resp_bits_pte_d(ptw_io_requestor_0_resp_bits_pte_d),
    .io_requestor_0_resp_bits_pte_a(ptw_io_requestor_0_resp_bits_pte_a),
    .io_requestor_0_resp_bits_pte_g(ptw_io_requestor_0_resp_bits_pte_g),
    .io_requestor_0_resp_bits_pte_u(ptw_io_requestor_0_resp_bits_pte_u),
    .io_requestor_0_resp_bits_pte_x(ptw_io_requestor_0_resp_bits_pte_x),
    .io_requestor_0_resp_bits_pte_w(ptw_io_requestor_0_resp_bits_pte_w),
    .io_requestor_0_resp_bits_pte_r(ptw_io_requestor_0_resp_bits_pte_r),
    .io_requestor_0_resp_bits_pte_v(ptw_io_requestor_0_resp_bits_pte_v),
    .io_requestor_0_resp_bits_level(ptw_io_requestor_0_resp_bits_level),
    .io_requestor_0_resp_bits_homogeneous(ptw_io_requestor_0_resp_bits_homogeneous),
    .io_requestor_0_ptbr_mode(ptw_io_requestor_0_ptbr_mode),
    .io_requestor_0_status_debug(ptw_io_requestor_0_status_debug),
    .io_requestor_0_status_dprv(ptw_io_requestor_0_status_dprv),
    .io_requestor_0_status_mxr(ptw_io_requestor_0_status_mxr),
    .io_requestor_0_status_sum(ptw_io_requestor_0_status_sum),
    .io_requestor_0_pmp_0_cfg_l(ptw_io_requestor_0_pmp_0_cfg_l),
    .io_requestor_0_pmp_0_cfg_a(ptw_io_requestor_0_pmp_0_cfg_a),
    .io_requestor_0_pmp_0_cfg_x(ptw_io_requestor_0_pmp_0_cfg_x),
    .io_requestor_0_pmp_0_cfg_w(ptw_io_requestor_0_pmp_0_cfg_w),
    .io_requestor_0_pmp_0_cfg_r(ptw_io_requestor_0_pmp_0_cfg_r),
    .io_requestor_0_pmp_0_addr(ptw_io_requestor_0_pmp_0_addr),
    .io_requestor_0_pmp_0_mask(ptw_io_requestor_0_pmp_0_mask),
    .io_requestor_0_pmp_1_cfg_l(ptw_io_requestor_0_pmp_1_cfg_l),
    .io_requestor_0_pmp_1_cfg_a(ptw_io_requestor_0_pmp_1_cfg_a),
    .io_requestor_0_pmp_1_cfg_x(ptw_io_requestor_0_pmp_1_cfg_x),
    .io_requestor_0_pmp_1_cfg_w(ptw_io_requestor_0_pmp_1_cfg_w),
    .io_requestor_0_pmp_1_cfg_r(ptw_io_requestor_0_pmp_1_cfg_r),
    .io_requestor_0_pmp_1_addr(ptw_io_requestor_0_pmp_1_addr),
    .io_requestor_0_pmp_1_mask(ptw_io_requestor_0_pmp_1_mask),
    .io_requestor_0_pmp_2_cfg_l(ptw_io_requestor_0_pmp_2_cfg_l),
    .io_requestor_0_pmp_2_cfg_a(ptw_io_requestor_0_pmp_2_cfg_a),
    .io_requestor_0_pmp_2_cfg_x(ptw_io_requestor_0_pmp_2_cfg_x),
    .io_requestor_0_pmp_2_cfg_w(ptw_io_requestor_0_pmp_2_cfg_w),
    .io_requestor_0_pmp_2_cfg_r(ptw_io_requestor_0_pmp_2_cfg_r),
    .io_requestor_0_pmp_2_addr(ptw_io_requestor_0_pmp_2_addr),
    .io_requestor_0_pmp_2_mask(ptw_io_requestor_0_pmp_2_mask),
    .io_requestor_0_pmp_3_cfg_l(ptw_io_requestor_0_pmp_3_cfg_l),
    .io_requestor_0_pmp_3_cfg_a(ptw_io_requestor_0_pmp_3_cfg_a),
    .io_requestor_0_pmp_3_cfg_x(ptw_io_requestor_0_pmp_3_cfg_x),
    .io_requestor_0_pmp_3_cfg_w(ptw_io_requestor_0_pmp_3_cfg_w),
    .io_requestor_0_pmp_3_cfg_r(ptw_io_requestor_0_pmp_3_cfg_r),
    .io_requestor_0_pmp_3_addr(ptw_io_requestor_0_pmp_3_addr),
    .io_requestor_0_pmp_3_mask(ptw_io_requestor_0_pmp_3_mask),
    .io_requestor_0_pmp_4_cfg_l(ptw_io_requestor_0_pmp_4_cfg_l),
    .io_requestor_0_pmp_4_cfg_a(ptw_io_requestor_0_pmp_4_cfg_a),
    .io_requestor_0_pmp_4_cfg_x(ptw_io_requestor_0_pmp_4_cfg_x),
    .io_requestor_0_pmp_4_cfg_w(ptw_io_requestor_0_pmp_4_cfg_w),
    .io_requestor_0_pmp_4_cfg_r(ptw_io_requestor_0_pmp_4_cfg_r),
    .io_requestor_0_pmp_4_addr(ptw_io_requestor_0_pmp_4_addr),
    .io_requestor_0_pmp_4_mask(ptw_io_requestor_0_pmp_4_mask),
    .io_requestor_0_pmp_5_cfg_l(ptw_io_requestor_0_pmp_5_cfg_l),
    .io_requestor_0_pmp_5_cfg_a(ptw_io_requestor_0_pmp_5_cfg_a),
    .io_requestor_0_pmp_5_cfg_x(ptw_io_requestor_0_pmp_5_cfg_x),
    .io_requestor_0_pmp_5_cfg_w(ptw_io_requestor_0_pmp_5_cfg_w),
    .io_requestor_0_pmp_5_cfg_r(ptw_io_requestor_0_pmp_5_cfg_r),
    .io_requestor_0_pmp_5_addr(ptw_io_requestor_0_pmp_5_addr),
    .io_requestor_0_pmp_5_mask(ptw_io_requestor_0_pmp_5_mask),
    .io_requestor_0_pmp_6_cfg_l(ptw_io_requestor_0_pmp_6_cfg_l),
    .io_requestor_0_pmp_6_cfg_a(ptw_io_requestor_0_pmp_6_cfg_a),
    .io_requestor_0_pmp_6_cfg_x(ptw_io_requestor_0_pmp_6_cfg_x),
    .io_requestor_0_pmp_6_cfg_w(ptw_io_requestor_0_pmp_6_cfg_w),
    .io_requestor_0_pmp_6_cfg_r(ptw_io_requestor_0_pmp_6_cfg_r),
    .io_requestor_0_pmp_6_addr(ptw_io_requestor_0_pmp_6_addr),
    .io_requestor_0_pmp_6_mask(ptw_io_requestor_0_pmp_6_mask),
    .io_requestor_0_pmp_7_cfg_l(ptw_io_requestor_0_pmp_7_cfg_l),
    .io_requestor_0_pmp_7_cfg_a(ptw_io_requestor_0_pmp_7_cfg_a),
    .io_requestor_0_pmp_7_cfg_x(ptw_io_requestor_0_pmp_7_cfg_x),
    .io_requestor_0_pmp_7_cfg_w(ptw_io_requestor_0_pmp_7_cfg_w),
    .io_requestor_0_pmp_7_cfg_r(ptw_io_requestor_0_pmp_7_cfg_r),
    .io_requestor_0_pmp_7_addr(ptw_io_requestor_0_pmp_7_addr),
    .io_requestor_0_pmp_7_mask(ptw_io_requestor_0_pmp_7_mask),
    .io_requestor_1_req_ready(ptw_io_requestor_1_req_ready),
    .io_requestor_1_req_valid(ptw_io_requestor_1_req_valid),
    .io_requestor_1_req_bits_valid(ptw_io_requestor_1_req_bits_valid),
    .io_requestor_1_req_bits_bits_addr(ptw_io_requestor_1_req_bits_bits_addr),
    .io_requestor_1_resp_valid(ptw_io_requestor_1_resp_valid),
    .io_requestor_1_resp_bits_ae(ptw_io_requestor_1_resp_bits_ae),
    .io_requestor_1_resp_bits_pte_ppn(ptw_io_requestor_1_resp_bits_pte_ppn),
    .io_requestor_1_resp_bits_pte_d(ptw_io_requestor_1_resp_bits_pte_d),
    .io_requestor_1_resp_bits_pte_a(ptw_io_requestor_1_resp_bits_pte_a),
    .io_requestor_1_resp_bits_pte_g(ptw_io_requestor_1_resp_bits_pte_g),
    .io_requestor_1_resp_bits_pte_u(ptw_io_requestor_1_resp_bits_pte_u),
    .io_requestor_1_resp_bits_pte_x(ptw_io_requestor_1_resp_bits_pte_x),
    .io_requestor_1_resp_bits_pte_w(ptw_io_requestor_1_resp_bits_pte_w),
    .io_requestor_1_resp_bits_pte_r(ptw_io_requestor_1_resp_bits_pte_r),
    .io_requestor_1_resp_bits_pte_v(ptw_io_requestor_1_resp_bits_pte_v),
    .io_requestor_1_resp_bits_level(ptw_io_requestor_1_resp_bits_level),
    .io_requestor_1_resp_bits_homogeneous(ptw_io_requestor_1_resp_bits_homogeneous),
    .io_requestor_1_ptbr_mode(ptw_io_requestor_1_ptbr_mode),
    .io_requestor_1_status_debug(ptw_io_requestor_1_status_debug),
    .io_requestor_1_status_prv(ptw_io_requestor_1_status_prv),
    .io_requestor_1_pmp_0_cfg_l(ptw_io_requestor_1_pmp_0_cfg_l),
    .io_requestor_1_pmp_0_cfg_a(ptw_io_requestor_1_pmp_0_cfg_a),
    .io_requestor_1_pmp_0_cfg_x(ptw_io_requestor_1_pmp_0_cfg_x),
    .io_requestor_1_pmp_0_cfg_w(ptw_io_requestor_1_pmp_0_cfg_w),
    .io_requestor_1_pmp_0_cfg_r(ptw_io_requestor_1_pmp_0_cfg_r),
    .io_requestor_1_pmp_0_addr(ptw_io_requestor_1_pmp_0_addr),
    .io_requestor_1_pmp_0_mask(ptw_io_requestor_1_pmp_0_mask),
    .io_requestor_1_pmp_1_cfg_l(ptw_io_requestor_1_pmp_1_cfg_l),
    .io_requestor_1_pmp_1_cfg_a(ptw_io_requestor_1_pmp_1_cfg_a),
    .io_requestor_1_pmp_1_cfg_x(ptw_io_requestor_1_pmp_1_cfg_x),
    .io_requestor_1_pmp_1_cfg_w(ptw_io_requestor_1_pmp_1_cfg_w),
    .io_requestor_1_pmp_1_cfg_r(ptw_io_requestor_1_pmp_1_cfg_r),
    .io_requestor_1_pmp_1_addr(ptw_io_requestor_1_pmp_1_addr),
    .io_requestor_1_pmp_1_mask(ptw_io_requestor_1_pmp_1_mask),
    .io_requestor_1_pmp_2_cfg_l(ptw_io_requestor_1_pmp_2_cfg_l),
    .io_requestor_1_pmp_2_cfg_a(ptw_io_requestor_1_pmp_2_cfg_a),
    .io_requestor_1_pmp_2_cfg_x(ptw_io_requestor_1_pmp_2_cfg_x),
    .io_requestor_1_pmp_2_cfg_w(ptw_io_requestor_1_pmp_2_cfg_w),
    .io_requestor_1_pmp_2_cfg_r(ptw_io_requestor_1_pmp_2_cfg_r),
    .io_requestor_1_pmp_2_addr(ptw_io_requestor_1_pmp_2_addr),
    .io_requestor_1_pmp_2_mask(ptw_io_requestor_1_pmp_2_mask),
    .io_requestor_1_pmp_3_cfg_l(ptw_io_requestor_1_pmp_3_cfg_l),
    .io_requestor_1_pmp_3_cfg_a(ptw_io_requestor_1_pmp_3_cfg_a),
    .io_requestor_1_pmp_3_cfg_x(ptw_io_requestor_1_pmp_3_cfg_x),
    .io_requestor_1_pmp_3_cfg_w(ptw_io_requestor_1_pmp_3_cfg_w),
    .io_requestor_1_pmp_3_cfg_r(ptw_io_requestor_1_pmp_3_cfg_r),
    .io_requestor_1_pmp_3_addr(ptw_io_requestor_1_pmp_3_addr),
    .io_requestor_1_pmp_3_mask(ptw_io_requestor_1_pmp_3_mask),
    .io_requestor_1_pmp_4_cfg_l(ptw_io_requestor_1_pmp_4_cfg_l),
    .io_requestor_1_pmp_4_cfg_a(ptw_io_requestor_1_pmp_4_cfg_a),
    .io_requestor_1_pmp_4_cfg_x(ptw_io_requestor_1_pmp_4_cfg_x),
    .io_requestor_1_pmp_4_cfg_w(ptw_io_requestor_1_pmp_4_cfg_w),
    .io_requestor_1_pmp_4_cfg_r(ptw_io_requestor_1_pmp_4_cfg_r),
    .io_requestor_1_pmp_4_addr(ptw_io_requestor_1_pmp_4_addr),
    .io_requestor_1_pmp_4_mask(ptw_io_requestor_1_pmp_4_mask),
    .io_requestor_1_pmp_5_cfg_l(ptw_io_requestor_1_pmp_5_cfg_l),
    .io_requestor_1_pmp_5_cfg_a(ptw_io_requestor_1_pmp_5_cfg_a),
    .io_requestor_1_pmp_5_cfg_x(ptw_io_requestor_1_pmp_5_cfg_x),
    .io_requestor_1_pmp_5_cfg_w(ptw_io_requestor_1_pmp_5_cfg_w),
    .io_requestor_1_pmp_5_cfg_r(ptw_io_requestor_1_pmp_5_cfg_r),
    .io_requestor_1_pmp_5_addr(ptw_io_requestor_1_pmp_5_addr),
    .io_requestor_1_pmp_5_mask(ptw_io_requestor_1_pmp_5_mask),
    .io_requestor_1_pmp_6_cfg_l(ptw_io_requestor_1_pmp_6_cfg_l),
    .io_requestor_1_pmp_6_cfg_a(ptw_io_requestor_1_pmp_6_cfg_a),
    .io_requestor_1_pmp_6_cfg_x(ptw_io_requestor_1_pmp_6_cfg_x),
    .io_requestor_1_pmp_6_cfg_w(ptw_io_requestor_1_pmp_6_cfg_w),
    .io_requestor_1_pmp_6_cfg_r(ptw_io_requestor_1_pmp_6_cfg_r),
    .io_requestor_1_pmp_6_addr(ptw_io_requestor_1_pmp_6_addr),
    .io_requestor_1_pmp_6_mask(ptw_io_requestor_1_pmp_6_mask),
    .io_requestor_1_pmp_7_cfg_l(ptw_io_requestor_1_pmp_7_cfg_l),
    .io_requestor_1_pmp_7_cfg_a(ptw_io_requestor_1_pmp_7_cfg_a),
    .io_requestor_1_pmp_7_cfg_x(ptw_io_requestor_1_pmp_7_cfg_x),
    .io_requestor_1_pmp_7_cfg_w(ptw_io_requestor_1_pmp_7_cfg_w),
    .io_requestor_1_pmp_7_cfg_r(ptw_io_requestor_1_pmp_7_cfg_r),
    .io_requestor_1_pmp_7_addr(ptw_io_requestor_1_pmp_7_addr),
    .io_requestor_1_pmp_7_mask(ptw_io_requestor_1_pmp_7_mask),
    .io_requestor_1_customCSRs_csrs_0_value(ptw_io_requestor_1_customCSRs_csrs_0_value),
    .io_mem_req_ready(ptw_io_mem_req_ready),
    .io_mem_req_valid(ptw_io_mem_req_valid),
    .io_mem_req_bits_addr(ptw_io_mem_req_bits_addr),
    .io_mem_s1_kill(ptw_io_mem_s1_kill),
    .io_mem_s2_nack(ptw_io_mem_s2_nack),
    .io_mem_resp_valid(ptw_io_mem_resp_valid),
    .io_mem_resp_bits_data(ptw_io_mem_resp_bits_data),
    .io_mem_s2_xcpt_ae_ld(ptw_io_mem_s2_xcpt_ae_ld),
    .io_dpath_ptbr_mode(ptw_io_dpath_ptbr_mode),
    .io_dpath_ptbr_ppn(ptw_io_dpath_ptbr_ppn),
    .io_dpath_sfence_valid(ptw_io_dpath_sfence_valid),
    .io_dpath_sfence_bits_rs1(ptw_io_dpath_sfence_bits_rs1),
    .io_dpath_status_debug(ptw_io_dpath_status_debug),
    .io_dpath_status_dprv(ptw_io_dpath_status_dprv),
    .io_dpath_status_prv(ptw_io_dpath_status_prv),
    .io_dpath_status_mxr(ptw_io_dpath_status_mxr),
    .io_dpath_status_sum(ptw_io_dpath_status_sum),
    .io_dpath_pmp_0_cfg_l(ptw_io_dpath_pmp_0_cfg_l),
    .io_dpath_pmp_0_cfg_a(ptw_io_dpath_pmp_0_cfg_a),
    .io_dpath_pmp_0_cfg_x(ptw_io_dpath_pmp_0_cfg_x),
    .io_dpath_pmp_0_cfg_w(ptw_io_dpath_pmp_0_cfg_w),
    .io_dpath_pmp_0_cfg_r(ptw_io_dpath_pmp_0_cfg_r),
    .io_dpath_pmp_0_addr(ptw_io_dpath_pmp_0_addr),
    .io_dpath_pmp_0_mask(ptw_io_dpath_pmp_0_mask),
    .io_dpath_pmp_1_cfg_l(ptw_io_dpath_pmp_1_cfg_l),
    .io_dpath_pmp_1_cfg_a(ptw_io_dpath_pmp_1_cfg_a),
    .io_dpath_pmp_1_cfg_x(ptw_io_dpath_pmp_1_cfg_x),
    .io_dpath_pmp_1_cfg_w(ptw_io_dpath_pmp_1_cfg_w),
    .io_dpath_pmp_1_cfg_r(ptw_io_dpath_pmp_1_cfg_r),
    .io_dpath_pmp_1_addr(ptw_io_dpath_pmp_1_addr),
    .io_dpath_pmp_1_mask(ptw_io_dpath_pmp_1_mask),
    .io_dpath_pmp_2_cfg_l(ptw_io_dpath_pmp_2_cfg_l),
    .io_dpath_pmp_2_cfg_a(ptw_io_dpath_pmp_2_cfg_a),
    .io_dpath_pmp_2_cfg_x(ptw_io_dpath_pmp_2_cfg_x),
    .io_dpath_pmp_2_cfg_w(ptw_io_dpath_pmp_2_cfg_w),
    .io_dpath_pmp_2_cfg_r(ptw_io_dpath_pmp_2_cfg_r),
    .io_dpath_pmp_2_addr(ptw_io_dpath_pmp_2_addr),
    .io_dpath_pmp_2_mask(ptw_io_dpath_pmp_2_mask),
    .io_dpath_pmp_3_cfg_l(ptw_io_dpath_pmp_3_cfg_l),
    .io_dpath_pmp_3_cfg_a(ptw_io_dpath_pmp_3_cfg_a),
    .io_dpath_pmp_3_cfg_x(ptw_io_dpath_pmp_3_cfg_x),
    .io_dpath_pmp_3_cfg_w(ptw_io_dpath_pmp_3_cfg_w),
    .io_dpath_pmp_3_cfg_r(ptw_io_dpath_pmp_3_cfg_r),
    .io_dpath_pmp_3_addr(ptw_io_dpath_pmp_3_addr),
    .io_dpath_pmp_3_mask(ptw_io_dpath_pmp_3_mask),
    .io_dpath_pmp_4_cfg_l(ptw_io_dpath_pmp_4_cfg_l),
    .io_dpath_pmp_4_cfg_a(ptw_io_dpath_pmp_4_cfg_a),
    .io_dpath_pmp_4_cfg_x(ptw_io_dpath_pmp_4_cfg_x),
    .io_dpath_pmp_4_cfg_w(ptw_io_dpath_pmp_4_cfg_w),
    .io_dpath_pmp_4_cfg_r(ptw_io_dpath_pmp_4_cfg_r),
    .io_dpath_pmp_4_addr(ptw_io_dpath_pmp_4_addr),
    .io_dpath_pmp_4_mask(ptw_io_dpath_pmp_4_mask),
    .io_dpath_pmp_5_cfg_l(ptw_io_dpath_pmp_5_cfg_l),
    .io_dpath_pmp_5_cfg_a(ptw_io_dpath_pmp_5_cfg_a),
    .io_dpath_pmp_5_cfg_x(ptw_io_dpath_pmp_5_cfg_x),
    .io_dpath_pmp_5_cfg_w(ptw_io_dpath_pmp_5_cfg_w),
    .io_dpath_pmp_5_cfg_r(ptw_io_dpath_pmp_5_cfg_r),
    .io_dpath_pmp_5_addr(ptw_io_dpath_pmp_5_addr),
    .io_dpath_pmp_5_mask(ptw_io_dpath_pmp_5_mask),
    .io_dpath_pmp_6_cfg_l(ptw_io_dpath_pmp_6_cfg_l),
    .io_dpath_pmp_6_cfg_a(ptw_io_dpath_pmp_6_cfg_a),
    .io_dpath_pmp_6_cfg_x(ptw_io_dpath_pmp_6_cfg_x),
    .io_dpath_pmp_6_cfg_w(ptw_io_dpath_pmp_6_cfg_w),
    .io_dpath_pmp_6_cfg_r(ptw_io_dpath_pmp_6_cfg_r),
    .io_dpath_pmp_6_addr(ptw_io_dpath_pmp_6_addr),
    .io_dpath_pmp_6_mask(ptw_io_dpath_pmp_6_mask),
    .io_dpath_pmp_7_cfg_l(ptw_io_dpath_pmp_7_cfg_l),
    .io_dpath_pmp_7_cfg_a(ptw_io_dpath_pmp_7_cfg_a),
    .io_dpath_pmp_7_cfg_x(ptw_io_dpath_pmp_7_cfg_x),
    .io_dpath_pmp_7_cfg_w(ptw_io_dpath_pmp_7_cfg_w),
    .io_dpath_pmp_7_cfg_r(ptw_io_dpath_pmp_7_cfg_r),
    .io_dpath_pmp_7_addr(ptw_io_dpath_pmp_7_addr),
    .io_dpath_pmp_7_mask(ptw_io_dpath_pmp_7_mask),
    .io_dpath_perf_l2hit(ptw_io_dpath_perf_l2hit),
    .io_dpath_perf_pte_miss(ptw_io_dpath_perf_pte_miss),
    .io_dpath_perf_pte_hit(ptw_io_dpath_perf_pte_hit),
    .io_dpath_customCSRs_csrs_0_value(ptw_io_dpath_customCSRs_csrs_0_value),
    .io_covSum(ptw_io_covSum),
    .metaAssert(ptw_metaAssert),
    .metaReset(ptw_metaReset)
  );
  Rocket core ( // @[RocketTile.scala 140:20]
    .clock(core_clock),
    .reset(core_reset),
    .io_hartid(core_io_hartid),
    .io_interrupts_debug(core_io_interrupts_debug),
    .io_interrupts_mtip(core_io_interrupts_mtip),
    .io_interrupts_msip(core_io_interrupts_msip),
    .io_interrupts_meip(core_io_interrupts_meip),
    .io_interrupts_seip(core_io_interrupts_seip),
    .io_imem_might_request(core_io_imem_might_request),
    .io_imem_req_valid(core_io_imem_req_valid),
    .io_imem_req_bits_pc(core_io_imem_req_bits_pc),
    .io_imem_req_bits_speculative(core_io_imem_req_bits_speculative),
    .io_imem_sfence_valid(core_io_imem_sfence_valid),
    .io_imem_sfence_bits_rs1(core_io_imem_sfence_bits_rs1),
    .io_imem_sfence_bits_rs2(core_io_imem_sfence_bits_rs2),
    .io_imem_sfence_bits_addr(core_io_imem_sfence_bits_addr),
    .io_imem_resp_ready(core_io_imem_resp_ready),
    .io_imem_resp_valid(core_io_imem_resp_valid),
    .io_imem_resp_bits_btb_taken(core_io_imem_resp_bits_btb_taken),
    .io_imem_resp_bits_btb_bridx(core_io_imem_resp_bits_btb_bridx),
    .io_imem_resp_bits_btb_entry(core_io_imem_resp_bits_btb_entry),
    .io_imem_resp_bits_btb_bht_history(core_io_imem_resp_bits_btb_bht_history),
    .io_imem_resp_bits_pc(core_io_imem_resp_bits_pc),
    .io_imem_resp_bits_data(core_io_imem_resp_bits_data),
    .io_imem_resp_bits_xcpt_pf_inst(core_io_imem_resp_bits_xcpt_pf_inst),
    .io_imem_resp_bits_xcpt_ae_inst(core_io_imem_resp_bits_xcpt_ae_inst),
    .io_imem_resp_bits_replay(core_io_imem_resp_bits_replay),
    .io_imem_btb_update_valid(core_io_imem_btb_update_valid),
    .io_imem_btb_update_bits_prediction_entry(core_io_imem_btb_update_bits_prediction_entry),
    .io_imem_btb_update_bits_pc(core_io_imem_btb_update_bits_pc),
    .io_imem_btb_update_bits_isValid(core_io_imem_btb_update_bits_isValid),
    .io_imem_btb_update_bits_br_pc(core_io_imem_btb_update_bits_br_pc),
    .io_imem_btb_update_bits_cfiType(core_io_imem_btb_update_bits_cfiType),
    .io_imem_bht_update_valid(core_io_imem_bht_update_valid),
    .io_imem_bht_update_bits_prediction_history(core_io_imem_bht_update_bits_prediction_history),
    .io_imem_bht_update_bits_pc(core_io_imem_bht_update_bits_pc),
    .io_imem_bht_update_bits_branch(core_io_imem_bht_update_bits_branch),
    .io_imem_bht_update_bits_taken(core_io_imem_bht_update_bits_taken),
    .io_imem_bht_update_bits_mispredict(core_io_imem_bht_update_bits_mispredict),
    .io_imem_flush_icache(core_io_imem_flush_icache),
    .io_dmem_req_ready(core_io_dmem_req_ready),
    .io_dmem_req_valid(core_io_dmem_req_valid),
    .io_dmem_req_bits_addr(core_io_dmem_req_bits_addr),
    .io_dmem_req_bits_tag(core_io_dmem_req_bits_tag),
    .io_dmem_req_bits_cmd(core_io_dmem_req_bits_cmd),
    .io_dmem_req_bits_size(core_io_dmem_req_bits_size),
    .io_dmem_req_bits_signed(core_io_dmem_req_bits_signed),
    .io_dmem_s1_kill(core_io_dmem_s1_kill),
    .io_dmem_s1_data_data(core_io_dmem_s1_data_data),
    .io_dmem_s2_nack(core_io_dmem_s2_nack),
    .io_dmem_resp_valid(core_io_dmem_resp_valid),
    .io_dmem_resp_bits_tag(core_io_dmem_resp_bits_tag),
    .io_dmem_resp_bits_size(core_io_dmem_resp_bits_size),
    .io_dmem_resp_bits_data(core_io_dmem_resp_bits_data),
    .io_dmem_resp_bits_replay(core_io_dmem_resp_bits_replay),
    .io_dmem_resp_bits_has_data(core_io_dmem_resp_bits_has_data),
    .io_dmem_resp_bits_data_word_bypass(core_io_dmem_resp_bits_data_word_bypass),
    .io_dmem_replay_next(core_io_dmem_replay_next),
    .io_dmem_s2_xcpt_ma_ld(core_io_dmem_s2_xcpt_ma_ld),
    .io_dmem_s2_xcpt_ma_st(core_io_dmem_s2_xcpt_ma_st),
    .io_dmem_s2_xcpt_pf_ld(core_io_dmem_s2_xcpt_pf_ld),
    .io_dmem_s2_xcpt_pf_st(core_io_dmem_s2_xcpt_pf_st),
    .io_dmem_s2_xcpt_ae_ld(core_io_dmem_s2_xcpt_ae_ld),
    .io_dmem_s2_xcpt_ae_st(core_io_dmem_s2_xcpt_ae_st),
    .io_dmem_ordered(core_io_dmem_ordered),
    .io_dmem_perf_release(core_io_dmem_perf_release),
    .io_dmem_perf_grant(core_io_dmem_perf_grant),
    .io_ptw_ptbr_mode(core_io_ptw_ptbr_mode),
    .io_ptw_ptbr_ppn(core_io_ptw_ptbr_ppn),
    .io_ptw_sfence_valid(core_io_ptw_sfence_valid),
    .io_ptw_sfence_bits_rs1(core_io_ptw_sfence_bits_rs1),
    .io_ptw_status_debug(core_io_ptw_status_debug),
    .io_ptw_status_dprv(core_io_ptw_status_dprv),
    .io_ptw_status_prv(core_io_ptw_status_prv),
    .io_ptw_status_mxr(core_io_ptw_status_mxr),
    .io_ptw_status_sum(core_io_ptw_status_sum),
    .io_ptw_pmp_0_cfg_l(core_io_ptw_pmp_0_cfg_l),
    .io_ptw_pmp_0_cfg_a(core_io_ptw_pmp_0_cfg_a),
    .io_ptw_pmp_0_cfg_x(core_io_ptw_pmp_0_cfg_x),
    .io_ptw_pmp_0_cfg_w(core_io_ptw_pmp_0_cfg_w),
    .io_ptw_pmp_0_cfg_r(core_io_ptw_pmp_0_cfg_r),
    .io_ptw_pmp_0_addr(core_io_ptw_pmp_0_addr),
    .io_ptw_pmp_0_mask(core_io_ptw_pmp_0_mask),
    .io_ptw_pmp_1_cfg_l(core_io_ptw_pmp_1_cfg_l),
    .io_ptw_pmp_1_cfg_a(core_io_ptw_pmp_1_cfg_a),
    .io_ptw_pmp_1_cfg_x(core_io_ptw_pmp_1_cfg_x),
    .io_ptw_pmp_1_cfg_w(core_io_ptw_pmp_1_cfg_w),
    .io_ptw_pmp_1_cfg_r(core_io_ptw_pmp_1_cfg_r),
    .io_ptw_pmp_1_addr(core_io_ptw_pmp_1_addr),
    .io_ptw_pmp_1_mask(core_io_ptw_pmp_1_mask),
    .io_ptw_pmp_2_cfg_l(core_io_ptw_pmp_2_cfg_l),
    .io_ptw_pmp_2_cfg_a(core_io_ptw_pmp_2_cfg_a),
    .io_ptw_pmp_2_cfg_x(core_io_ptw_pmp_2_cfg_x),
    .io_ptw_pmp_2_cfg_w(core_io_ptw_pmp_2_cfg_w),
    .io_ptw_pmp_2_cfg_r(core_io_ptw_pmp_2_cfg_r),
    .io_ptw_pmp_2_addr(core_io_ptw_pmp_2_addr),
    .io_ptw_pmp_2_mask(core_io_ptw_pmp_2_mask),
    .io_ptw_pmp_3_cfg_l(core_io_ptw_pmp_3_cfg_l),
    .io_ptw_pmp_3_cfg_a(core_io_ptw_pmp_3_cfg_a),
    .io_ptw_pmp_3_cfg_x(core_io_ptw_pmp_3_cfg_x),
    .io_ptw_pmp_3_cfg_w(core_io_ptw_pmp_3_cfg_w),
    .io_ptw_pmp_3_cfg_r(core_io_ptw_pmp_3_cfg_r),
    .io_ptw_pmp_3_addr(core_io_ptw_pmp_3_addr),
    .io_ptw_pmp_3_mask(core_io_ptw_pmp_3_mask),
    .io_ptw_pmp_4_cfg_l(core_io_ptw_pmp_4_cfg_l),
    .io_ptw_pmp_4_cfg_a(core_io_ptw_pmp_4_cfg_a),
    .io_ptw_pmp_4_cfg_x(core_io_ptw_pmp_4_cfg_x),
    .io_ptw_pmp_4_cfg_w(core_io_ptw_pmp_4_cfg_w),
    .io_ptw_pmp_4_cfg_r(core_io_ptw_pmp_4_cfg_r),
    .io_ptw_pmp_4_addr(core_io_ptw_pmp_4_addr),
    .io_ptw_pmp_4_mask(core_io_ptw_pmp_4_mask),
    .io_ptw_pmp_5_cfg_l(core_io_ptw_pmp_5_cfg_l),
    .io_ptw_pmp_5_cfg_a(core_io_ptw_pmp_5_cfg_a),
    .io_ptw_pmp_5_cfg_x(core_io_ptw_pmp_5_cfg_x),
    .io_ptw_pmp_5_cfg_w(core_io_ptw_pmp_5_cfg_w),
    .io_ptw_pmp_5_cfg_r(core_io_ptw_pmp_5_cfg_r),
    .io_ptw_pmp_5_addr(core_io_ptw_pmp_5_addr),
    .io_ptw_pmp_5_mask(core_io_ptw_pmp_5_mask),
    .io_ptw_pmp_6_cfg_l(core_io_ptw_pmp_6_cfg_l),
    .io_ptw_pmp_6_cfg_a(core_io_ptw_pmp_6_cfg_a),
    .io_ptw_pmp_6_cfg_x(core_io_ptw_pmp_6_cfg_x),
    .io_ptw_pmp_6_cfg_w(core_io_ptw_pmp_6_cfg_w),
    .io_ptw_pmp_6_cfg_r(core_io_ptw_pmp_6_cfg_r),
    .io_ptw_pmp_6_addr(core_io_ptw_pmp_6_addr),
    .io_ptw_pmp_6_mask(core_io_ptw_pmp_6_mask),
    .io_ptw_pmp_7_cfg_l(core_io_ptw_pmp_7_cfg_l),
    .io_ptw_pmp_7_cfg_a(core_io_ptw_pmp_7_cfg_a),
    .io_ptw_pmp_7_cfg_x(core_io_ptw_pmp_7_cfg_x),
    .io_ptw_pmp_7_cfg_w(core_io_ptw_pmp_7_cfg_w),
    .io_ptw_pmp_7_cfg_r(core_io_ptw_pmp_7_cfg_r),
    .io_ptw_pmp_7_addr(core_io_ptw_pmp_7_addr),
    .io_ptw_pmp_7_mask(core_io_ptw_pmp_7_mask),
    .io_ptw_customCSRs_csrs_0_value(core_io_ptw_customCSRs_csrs_0_value),
    .io_fpu_inst(core_io_fpu_inst),
    .io_fpu_fromint_data(core_io_fpu_fromint_data),
    .io_fpu_fcsr_rm(core_io_fpu_fcsr_rm),
    .io_fpu_fcsr_flags_valid(core_io_fpu_fcsr_flags_valid),
    .io_fpu_fcsr_flags_bits(core_io_fpu_fcsr_flags_bits),
    .io_fpu_store_data(core_io_fpu_store_data),
    .io_fpu_toint_data(core_io_fpu_toint_data),
    .io_fpu_dmem_resp_val(core_io_fpu_dmem_resp_val),
    .io_fpu_dmem_resp_type(core_io_fpu_dmem_resp_type),
    .io_fpu_dmem_resp_tag(core_io_fpu_dmem_resp_tag),
    .io_fpu_dmem_resp_data(core_io_fpu_dmem_resp_data),
    .io_fpu_valid(core_io_fpu_valid),
    .io_fpu_fcsr_rdy(core_io_fpu_fcsr_rdy),
    .io_fpu_nack_mem(core_io_fpu_nack_mem),
    .io_fpu_illegal_rm(core_io_fpu_illegal_rm),
    .io_fpu_killx(core_io_fpu_killx),
    .io_fpu_killm(core_io_fpu_killm),
    .io_fpu_dec_wen(core_io_fpu_dec_wen),
    .io_fpu_dec_ren1(core_io_fpu_dec_ren1),
    .io_fpu_dec_ren2(core_io_fpu_dec_ren2),
    .io_fpu_dec_ren3(core_io_fpu_dec_ren3),
    .io_fpu_sboard_set(core_io_fpu_sboard_set),
    .io_fpu_sboard_clr(core_io_fpu_sboard_clr),
    .io_fpu_sboard_clra(core_io_fpu_sboard_clra),
    .io_trace_0_valid(core_io_trace_0_valid),
    .io_trace_0_iaddr(core_io_trace_0_iaddr),
    .io_trace_0_insn(core_io_trace_0_insn),
    .io_trace_0_priv(core_io_trace_0_priv),
    .io_trace_0_exception(core_io_trace_0_exception),
    .io_trace_0_interrupt(core_io_trace_0_interrupt),
    .io_trace_0_cause(core_io_trace_0_cause),
    .io_trace_0_tval(core_io_trace_0_tval),
    .io_wfi(core_io_wfi),
    .io_covSum(core_io_covSum),
    .metaAssert(core_metaAssert),
    .metaReset(core_metaReset),
    .PlusArgTimeout_halt(core_PlusArgTimeout_halt),
    .csr_halt(core_csr_halt),
    .ibuf_halt(core_ibuf_halt),
    .div_halt(core_div_halt)
  );
  assign auto_broadcast_out_0_valid = broadcast_3_auto_out_0_valid; // @[LazyModule.scala 311:12]
  assign auto_broadcast_out_0_iaddr = broadcast_3_auto_out_0_iaddr; // @[LazyModule.scala 311:12]
  assign auto_broadcast_out_0_insn = broadcast_3_auto_out_0_insn; // @[LazyModule.scala 311:12]
  assign auto_broadcast_out_0_priv = broadcast_3_auto_out_0_priv; // @[LazyModule.scala 311:12]
  assign auto_broadcast_out_0_exception = broadcast_3_auto_out_0_exception; // @[LazyModule.scala 311:12]
  assign auto_broadcast_out_0_interrupt = broadcast_3_auto_out_0_interrupt; // @[LazyModule.scala 311:12]
  assign auto_broadcast_out_0_cause = broadcast_3_auto_out_0_cause; // @[LazyModule.scala 311:12]
  assign auto_broadcast_out_0_tval = broadcast_3_auto_out_0_tval; // @[LazyModule.scala 311:12]
  assign auto_wfi_out_0 = bundleOut_0_0_REG; // @[LazyModule.scala 311:12]
  assign auto_cease_out_0 = 1'h0; // @[LazyModule.scala 311:12]
  assign auto_halt_out_0 = 1'h0; // @[LazyModule.scala 311:12]
  assign auto_trace_core_source_out_group_0_iretire = 1'h0; // @[LazyModule.scala 311:12]
  assign auto_trace_core_source_out_group_0_iaddr = 32'h0; // @[LazyModule.scala 311:12]
  assign auto_trace_core_source_out_group_0_itype = 4'h0; // @[LazyModule.scala 311:12]
  assign auto_trace_core_source_out_group_0_ilastsize = 1'h0; // @[LazyModule.scala 311:12]
  assign auto_trace_core_source_out_priv = 4'h0; // @[LazyModule.scala 311:12]
  assign auto_trace_core_source_out_tval = 32'h0; // @[LazyModule.scala 311:12]
  assign auto_trace_core_source_out_cause = 32'h0; // @[LazyModule.scala 311:12]
  assign auto_tl_master_xing_out_a_valid = tlMasterXbar_auto_out_a_valid; // @[LazyModule.scala 311:12]
  assign auto_tl_master_xing_out_a_bits_opcode = tlMasterXbar_auto_out_a_bits_opcode; // @[LazyModule.scala 311:12]
  assign auto_tl_master_xing_out_a_bits_param = tlMasterXbar_auto_out_a_bits_param; // @[LazyModule.scala 311:12]
  assign auto_tl_master_xing_out_a_bits_size = tlMasterXbar_auto_out_a_bits_size; // @[LazyModule.scala 311:12]
  assign auto_tl_master_xing_out_a_bits_source = tlMasterXbar_auto_out_a_bits_source; // @[LazyModule.scala 311:12]
  assign auto_tl_master_xing_out_a_bits_address = tlMasterXbar_auto_out_a_bits_address; // @[LazyModule.scala 311:12]
  assign auto_tl_master_xing_out_a_bits_mask = tlMasterXbar_auto_out_a_bits_mask; // @[LazyModule.scala 311:12]
  assign auto_tl_master_xing_out_a_bits_data = tlMasterXbar_auto_out_a_bits_data; // @[LazyModule.scala 311:12]
  assign auto_tl_master_xing_out_a_bits_corrupt = 1'h0; // @[LazyModule.scala 311:12]
  assign auto_tl_master_xing_out_b_ready = tlMasterXbar_auto_out_b_ready; // @[LazyModule.scala 311:12]
  assign auto_tl_master_xing_out_c_valid = tlMasterXbar_auto_out_c_valid; // @[LazyModule.scala 311:12]
  assign auto_tl_master_xing_out_c_bits_opcode = tlMasterXbar_auto_out_c_bits_opcode; // @[LazyModule.scala 311:12]
  assign auto_tl_master_xing_out_c_bits_param = tlMasterXbar_auto_out_c_bits_param; // @[LazyModule.scala 311:12]
  assign auto_tl_master_xing_out_c_bits_size = tlMasterXbar_auto_out_c_bits_size; // @[LazyModule.scala 311:12]
  assign auto_tl_master_xing_out_c_bits_source = tlMasterXbar_auto_out_c_bits_source; // @[LazyModule.scala 311:12]
  assign auto_tl_master_xing_out_c_bits_address = tlMasterXbar_auto_out_c_bits_address; // @[LazyModule.scala 311:12]
  assign auto_tl_master_xing_out_c_bits_data = tlMasterXbar_auto_out_c_bits_data; // @[LazyModule.scala 311:12]
  assign auto_tl_master_xing_out_c_bits_corrupt = 1'h0; // @[LazyModule.scala 311:12]
  assign auto_tl_master_xing_out_d_ready = tlMasterXbar_auto_out_d_ready; // @[LazyModule.scala 311:12]
  assign auto_tl_master_xing_out_e_valid = tlMasterXbar_auto_out_e_valid; // @[LazyModule.scala 311:12]
  assign auto_tl_master_xing_out_e_bits_sink = tlMasterXbar_auto_out_e_bits_sink; // @[LazyModule.scala 311:12]
  assign tlMasterXbar_clock = clock;
  assign tlMasterXbar_reset = reset;
  assign tlMasterXbar_auto_in_1_a_valid = frontend_auto_icache_master_out_a_valid; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_1_a_bits_address = frontend_auto_icache_master_out_a_bits_address; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_0_a_valid = dcache_auto_out_a_valid; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_0_a_bits_opcode = dcache_auto_out_a_bits_opcode; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_0_a_bits_param = dcache_auto_out_a_bits_param; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_0_a_bits_size = dcache_auto_out_a_bits_size; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_0_a_bits_source = dcache_auto_out_a_bits_source; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_0_a_bits_address = dcache_auto_out_a_bits_address; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_0_a_bits_mask = dcache_auto_out_a_bits_mask; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_0_a_bits_data = dcache_auto_out_a_bits_data; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_0_b_ready = dcache_auto_out_b_ready; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_0_c_valid = dcache_auto_out_c_valid; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_0_c_bits_opcode = dcache_auto_out_c_bits_opcode; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_0_c_bits_param = dcache_auto_out_c_bits_param; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_0_c_bits_size = dcache_auto_out_c_bits_size; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_0_c_bits_source = dcache_auto_out_c_bits_source; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_0_c_bits_address = dcache_auto_out_c_bits_address; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_0_c_bits_data = dcache_auto_out_c_bits_data; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_0_d_ready = dcache_auto_out_d_ready; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_0_e_valid = dcache_auto_out_e_valid; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_in_0_e_bits_sink = dcache_auto_out_e_bits_sink; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_out_a_ready = auto_tl_master_xing_out_a_ready; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_out_b_valid = auto_tl_master_xing_out_b_valid; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_out_b_bits_opcode = auto_tl_master_xing_out_b_bits_opcode; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_out_b_bits_param = auto_tl_master_xing_out_b_bits_param; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_out_b_bits_size = auto_tl_master_xing_out_b_bits_size; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_out_b_bits_source = auto_tl_master_xing_out_b_bits_source; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_out_b_bits_address = auto_tl_master_xing_out_b_bits_address; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_out_b_bits_mask = auto_tl_master_xing_out_b_bits_mask; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_out_b_bits_corrupt = auto_tl_master_xing_out_b_bits_corrupt; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_out_c_ready = auto_tl_master_xing_out_c_ready; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_out_d_valid = auto_tl_master_xing_out_d_valid; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_out_d_bits_opcode = auto_tl_master_xing_out_d_bits_opcode; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_out_d_bits_param = auto_tl_master_xing_out_d_bits_param; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_out_d_bits_size = auto_tl_master_xing_out_d_bits_size; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_out_d_bits_source = auto_tl_master_xing_out_d_bits_source; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_out_d_bits_sink = auto_tl_master_xing_out_d_bits_sink; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_out_d_bits_denied = auto_tl_master_xing_out_d_bits_denied; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_out_d_bits_data = auto_tl_master_xing_out_d_bits_data; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_out_d_bits_corrupt = auto_tl_master_xing_out_d_bits_corrupt; // @[LazyModule.scala 296:16]
  assign tlMasterXbar_auto_out_e_ready = auto_tl_master_xing_out_e_ready; // @[LazyModule.scala 296:16]
  assign intXbar_auto_int_in_3_0 = auto_int_in_xing_in_2_sync_0; // @[LazyModule.scala 298:16]
  assign intXbar_auto_int_in_2_0 = auto_int_in_xing_in_1_sync_0; // @[LazyModule.scala 298:16]
  assign intXbar_auto_int_in_1_0 = auto_int_in_xing_in_0_sync_0; // @[LazyModule.scala 298:16]
  assign intXbar_auto_int_in_1_1 = auto_int_in_xing_in_0_sync_1; // @[LazyModule.scala 298:16]
  assign intXbar_auto_int_in_0_0 = auto_intsink_in_sync_0; // @[LazyModule.scala 298:16]
  assign broadcast_auto_in = auto_hartid_in; // @[LazyModule.scala 298:16]
  assign broadcast_1_auto_in = auto_reset_vector_in; // @[LazyModule.scala 298:16]
  assign broadcast_3_auto_in_0_valid = core_io_trace_0_valid; // @[LazyModule.scala 298:16]
  assign broadcast_3_auto_in_0_iaddr = core_io_trace_0_iaddr; // @[LazyModule.scala 298:16]
  assign broadcast_3_auto_in_0_insn = core_io_trace_0_insn; // @[LazyModule.scala 298:16]
  assign broadcast_3_auto_in_0_priv = core_io_trace_0_priv; // @[LazyModule.scala 298:16]
  assign broadcast_3_auto_in_0_exception = core_io_trace_0_exception; // @[LazyModule.scala 298:16]
  assign broadcast_3_auto_in_0_interrupt = core_io_trace_0_interrupt; // @[LazyModule.scala 298:16]
  assign broadcast_3_auto_in_0_cause = core_io_trace_0_cause; // @[LazyModule.scala 298:16]
  assign broadcast_3_auto_in_0_tval = core_io_trace_0_tval; // @[LazyModule.scala 298:16]
  assign dcache_gated_clock = clock;
  assign dcache_reset = reset;
  assign dcache_auto_out_a_ready = tlMasterXbar_auto_in_0_a_ready; // @[LazyModule.scala 296:16]
  assign dcache_auto_out_b_valid = tlMasterXbar_auto_in_0_b_valid; // @[LazyModule.scala 296:16]
  assign dcache_auto_out_b_bits_param = tlMasterXbar_auto_in_0_b_bits_param; // @[LazyModule.scala 296:16]
  assign dcache_auto_out_b_bits_size = tlMasterXbar_auto_in_0_b_bits_size; // @[LazyModule.scala 296:16]
  assign dcache_auto_out_b_bits_source = tlMasterXbar_auto_in_0_b_bits_source; // @[LazyModule.scala 296:16]
  assign dcache_auto_out_b_bits_address = tlMasterXbar_auto_in_0_b_bits_address; // @[LazyModule.scala 296:16]
  assign dcache_auto_out_c_ready = tlMasterXbar_auto_in_0_c_ready; // @[LazyModule.scala 296:16]
  assign dcache_auto_out_d_valid = tlMasterXbar_auto_in_0_d_valid; // @[LazyModule.scala 296:16]
  assign dcache_auto_out_d_bits_opcode = tlMasterXbar_auto_in_0_d_bits_opcode; // @[LazyModule.scala 296:16]
  assign dcache_auto_out_d_bits_param = tlMasterXbar_auto_in_0_d_bits_param; // @[LazyModule.scala 296:16]
  assign dcache_auto_out_d_bits_size = tlMasterXbar_auto_in_0_d_bits_size; // @[LazyModule.scala 296:16]
  assign dcache_auto_out_d_bits_source = tlMasterXbar_auto_in_0_d_bits_source; // @[LazyModule.scala 296:16]
  assign dcache_auto_out_d_bits_sink = tlMasterXbar_auto_in_0_d_bits_sink; // @[LazyModule.scala 296:16]
  assign dcache_auto_out_d_bits_denied = tlMasterXbar_auto_in_0_d_bits_denied; // @[LazyModule.scala 296:16]
  assign dcache_auto_out_d_bits_data = tlMasterXbar_auto_in_0_d_bits_data; // @[LazyModule.scala 296:16]
  assign dcache_auto_out_e_ready = tlMasterXbar_auto_in_0_e_ready; // @[LazyModule.scala 296:16]
  assign dcache_io_cpu_req_valid = dcacheArb_io_mem_req_valid; // @[HellaCache.scala 277:30]
  assign dcache_io_cpu_req_bits_addr = dcacheArb_io_mem_req_bits_addr; // @[HellaCache.scala 277:30]
  assign dcache_io_cpu_req_bits_tag = dcacheArb_io_mem_req_bits_tag; // @[HellaCache.scala 277:30]
  assign dcache_io_cpu_req_bits_cmd = dcacheArb_io_mem_req_bits_cmd; // @[HellaCache.scala 277:30]
  assign dcache_io_cpu_req_bits_size = dcacheArb_io_mem_req_bits_size; // @[HellaCache.scala 277:30]
  assign dcache_io_cpu_req_bits_signed = dcacheArb_io_mem_req_bits_signed; // @[HellaCache.scala 277:30]
  assign dcache_io_cpu_req_bits_phys = dcacheArb_io_mem_req_bits_phys; // @[HellaCache.scala 277:30]
  assign dcache_io_cpu_s1_kill = dcacheArb_io_mem_s1_kill; // @[HellaCache.scala 277:30]
  assign dcache_io_cpu_s1_data_data = dcacheArb_io_mem_s1_data_data; // @[HellaCache.scala 277:30]
  assign dcache_io_ptw_req_ready = ptw_io_requestor_0_req_ready; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_resp_valid = ptw_io_requestor_0_resp_valid; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_resp_bits_ae = ptw_io_requestor_0_resp_bits_ae; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_resp_bits_pte_ppn = ptw_io_requestor_0_resp_bits_pte_ppn; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_resp_bits_pte_d = ptw_io_requestor_0_resp_bits_pte_d; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_resp_bits_pte_a = ptw_io_requestor_0_resp_bits_pte_a; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_resp_bits_pte_g = ptw_io_requestor_0_resp_bits_pte_g; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_resp_bits_pte_u = ptw_io_requestor_0_resp_bits_pte_u; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_resp_bits_pte_x = ptw_io_requestor_0_resp_bits_pte_x; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_resp_bits_pte_w = ptw_io_requestor_0_resp_bits_pte_w; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_resp_bits_pte_r = ptw_io_requestor_0_resp_bits_pte_r; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_resp_bits_pte_v = ptw_io_requestor_0_resp_bits_pte_v; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_resp_bits_level = ptw_io_requestor_0_resp_bits_level; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_resp_bits_homogeneous = ptw_io_requestor_0_resp_bits_homogeneous; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_ptbr_mode = ptw_io_requestor_0_ptbr_mode; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_status_debug = ptw_io_requestor_0_status_debug; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_status_dprv = ptw_io_requestor_0_status_dprv; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_status_mxr = ptw_io_requestor_0_status_mxr; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_status_sum = ptw_io_requestor_0_status_sum; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_0_cfg_l = ptw_io_requestor_0_pmp_0_cfg_l; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_0_cfg_a = ptw_io_requestor_0_pmp_0_cfg_a; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_0_cfg_x = ptw_io_requestor_0_pmp_0_cfg_x; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_0_cfg_w = ptw_io_requestor_0_pmp_0_cfg_w; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_0_cfg_r = ptw_io_requestor_0_pmp_0_cfg_r; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_0_addr = ptw_io_requestor_0_pmp_0_addr; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_0_mask = ptw_io_requestor_0_pmp_0_mask; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_1_cfg_l = ptw_io_requestor_0_pmp_1_cfg_l; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_1_cfg_a = ptw_io_requestor_0_pmp_1_cfg_a; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_1_cfg_x = ptw_io_requestor_0_pmp_1_cfg_x; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_1_cfg_w = ptw_io_requestor_0_pmp_1_cfg_w; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_1_cfg_r = ptw_io_requestor_0_pmp_1_cfg_r; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_1_addr = ptw_io_requestor_0_pmp_1_addr; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_1_mask = ptw_io_requestor_0_pmp_1_mask; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_2_cfg_l = ptw_io_requestor_0_pmp_2_cfg_l; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_2_cfg_a = ptw_io_requestor_0_pmp_2_cfg_a; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_2_cfg_x = ptw_io_requestor_0_pmp_2_cfg_x; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_2_cfg_w = ptw_io_requestor_0_pmp_2_cfg_w; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_2_cfg_r = ptw_io_requestor_0_pmp_2_cfg_r; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_2_addr = ptw_io_requestor_0_pmp_2_addr; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_2_mask = ptw_io_requestor_0_pmp_2_mask; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_3_cfg_l = ptw_io_requestor_0_pmp_3_cfg_l; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_3_cfg_a = ptw_io_requestor_0_pmp_3_cfg_a; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_3_cfg_x = ptw_io_requestor_0_pmp_3_cfg_x; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_3_cfg_w = ptw_io_requestor_0_pmp_3_cfg_w; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_3_cfg_r = ptw_io_requestor_0_pmp_3_cfg_r; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_3_addr = ptw_io_requestor_0_pmp_3_addr; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_3_mask = ptw_io_requestor_0_pmp_3_mask; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_4_cfg_l = ptw_io_requestor_0_pmp_4_cfg_l; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_4_cfg_a = ptw_io_requestor_0_pmp_4_cfg_a; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_4_cfg_x = ptw_io_requestor_0_pmp_4_cfg_x; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_4_cfg_w = ptw_io_requestor_0_pmp_4_cfg_w; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_4_cfg_r = ptw_io_requestor_0_pmp_4_cfg_r; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_4_addr = ptw_io_requestor_0_pmp_4_addr; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_4_mask = ptw_io_requestor_0_pmp_4_mask; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_5_cfg_l = ptw_io_requestor_0_pmp_5_cfg_l; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_5_cfg_a = ptw_io_requestor_0_pmp_5_cfg_a; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_5_cfg_x = ptw_io_requestor_0_pmp_5_cfg_x; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_5_cfg_w = ptw_io_requestor_0_pmp_5_cfg_w; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_5_cfg_r = ptw_io_requestor_0_pmp_5_cfg_r; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_5_addr = ptw_io_requestor_0_pmp_5_addr; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_5_mask = ptw_io_requestor_0_pmp_5_mask; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_6_cfg_l = ptw_io_requestor_0_pmp_6_cfg_l; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_6_cfg_a = ptw_io_requestor_0_pmp_6_cfg_a; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_6_cfg_x = ptw_io_requestor_0_pmp_6_cfg_x; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_6_cfg_w = ptw_io_requestor_0_pmp_6_cfg_w; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_6_cfg_r = ptw_io_requestor_0_pmp_6_cfg_r; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_6_addr = ptw_io_requestor_0_pmp_6_addr; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_6_mask = ptw_io_requestor_0_pmp_6_mask; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_7_cfg_l = ptw_io_requestor_0_pmp_7_cfg_l; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_7_cfg_a = ptw_io_requestor_0_pmp_7_cfg_a; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_7_cfg_x = ptw_io_requestor_0_pmp_7_cfg_x; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_7_cfg_w = ptw_io_requestor_0_pmp_7_cfg_w; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_7_cfg_r = ptw_io_requestor_0_pmp_7_cfg_r; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_7_addr = ptw_io_requestor_0_pmp_7_addr; // @[RocketTile.scala 198:20]
  assign dcache_io_ptw_pmp_7_mask = ptw_io_requestor_0_pmp_7_mask; // @[RocketTile.scala 198:20]
  assign frontend_gated_clock = clock;
  assign frontend_reset = reset;
  assign frontend_auto_icache_master_out_a_ready = tlMasterXbar_auto_in_1_a_ready; // @[LazyModule.scala 296:16]
  assign frontend_auto_icache_master_out_d_valid = tlMasterXbar_auto_in_1_d_valid; // @[LazyModule.scala 296:16]
  assign frontend_auto_icache_master_out_d_bits_opcode = tlMasterXbar_auto_in_1_d_bits_opcode; // @[LazyModule.scala 296:16]
  assign frontend_auto_icache_master_out_d_bits_size = tlMasterXbar_auto_in_1_d_bits_size; // @[LazyModule.scala 296:16]
  assign frontend_auto_icache_master_out_d_bits_data = tlMasterXbar_auto_in_1_d_bits_data; // @[LazyModule.scala 296:16]
  assign frontend_auto_icache_master_out_d_bits_corrupt = tlMasterXbar_auto_in_1_d_bits_corrupt; // @[LazyModule.scala 296:16]
  assign frontend_auto_reset_vector_sink_in = broadcast_1_auto_out_1; // @[LazyModule.scala 298:16]
  assign frontend_io_cpu_might_request = core_io_imem_might_request; // @[RocketTile.scala 173:32]
  assign frontend_io_cpu_req_valid = core_io_imem_req_valid; // @[RocketTile.scala 173:32]
  assign frontend_io_cpu_req_bits_pc = core_io_imem_req_bits_pc; // @[RocketTile.scala 173:32]
  assign frontend_io_cpu_req_bits_speculative = core_io_imem_req_bits_speculative; // @[RocketTile.scala 173:32]
  assign frontend_io_cpu_sfence_valid = core_io_imem_sfence_valid; // @[RocketTile.scala 173:32]
  assign frontend_io_cpu_sfence_bits_rs1 = core_io_imem_sfence_bits_rs1; // @[RocketTile.scala 173:32]
  assign frontend_io_cpu_sfence_bits_rs2 = core_io_imem_sfence_bits_rs2; // @[RocketTile.scala 173:32]
  assign frontend_io_cpu_sfence_bits_addr = core_io_imem_sfence_bits_addr; // @[RocketTile.scala 173:32]
  assign frontend_io_cpu_resp_ready = core_io_imem_resp_ready; // @[RocketTile.scala 173:32]
  assign frontend_io_cpu_btb_update_valid = core_io_imem_btb_update_valid; // @[RocketTile.scala 173:32]
  assign frontend_io_cpu_btb_update_bits_prediction_entry = core_io_imem_btb_update_bits_prediction_entry; // @[RocketTile.scala 173:32]
  assign frontend_io_cpu_btb_update_bits_pc = core_io_imem_btb_update_bits_pc; // @[RocketTile.scala 173:32]
  assign frontend_io_cpu_btb_update_bits_isValid = core_io_imem_btb_update_bits_isValid; // @[RocketTile.scala 173:32]
  assign frontend_io_cpu_btb_update_bits_br_pc = core_io_imem_btb_update_bits_br_pc; // @[RocketTile.scala 173:32]
  assign frontend_io_cpu_btb_update_bits_cfiType = core_io_imem_btb_update_bits_cfiType; // @[RocketTile.scala 173:32]
  assign frontend_io_cpu_bht_update_valid = core_io_imem_bht_update_valid; // @[RocketTile.scala 173:32]
  assign frontend_io_cpu_bht_update_bits_prediction_history = core_io_imem_bht_update_bits_prediction_history; // @[RocketTile.scala 173:32]
  assign frontend_io_cpu_bht_update_bits_pc = core_io_imem_bht_update_bits_pc; // @[RocketTile.scala 173:32]
  assign frontend_io_cpu_bht_update_bits_branch = core_io_imem_bht_update_bits_branch; // @[RocketTile.scala 173:32]
  assign frontend_io_cpu_bht_update_bits_taken = core_io_imem_bht_update_bits_taken; // @[RocketTile.scala 173:32]
  assign frontend_io_cpu_bht_update_bits_mispredict = core_io_imem_bht_update_bits_mispredict; // @[RocketTile.scala 173:32]
  assign frontend_io_cpu_flush_icache = core_io_imem_flush_icache; // @[RocketTile.scala 173:32]
  assign frontend_io_ptw_req_ready = ptw_io_requestor_1_req_ready; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_resp_valid = ptw_io_requestor_1_resp_valid; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_resp_bits_ae = ptw_io_requestor_1_resp_bits_ae; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_resp_bits_pte_ppn = ptw_io_requestor_1_resp_bits_pte_ppn; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_resp_bits_pte_d = ptw_io_requestor_1_resp_bits_pte_d; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_resp_bits_pte_a = ptw_io_requestor_1_resp_bits_pte_a; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_resp_bits_pte_g = ptw_io_requestor_1_resp_bits_pte_g; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_resp_bits_pte_u = ptw_io_requestor_1_resp_bits_pte_u; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_resp_bits_pte_x = ptw_io_requestor_1_resp_bits_pte_x; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_resp_bits_pte_w = ptw_io_requestor_1_resp_bits_pte_w; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_resp_bits_pte_r = ptw_io_requestor_1_resp_bits_pte_r; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_resp_bits_pte_v = ptw_io_requestor_1_resp_bits_pte_v; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_resp_bits_level = ptw_io_requestor_1_resp_bits_level; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_resp_bits_homogeneous = ptw_io_requestor_1_resp_bits_homogeneous; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_ptbr_mode = ptw_io_requestor_1_ptbr_mode; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_status_debug = ptw_io_requestor_1_status_debug; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_status_prv = ptw_io_requestor_1_status_prv; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_0_cfg_l = ptw_io_requestor_1_pmp_0_cfg_l; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_0_cfg_a = ptw_io_requestor_1_pmp_0_cfg_a; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_0_cfg_x = ptw_io_requestor_1_pmp_0_cfg_x; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_0_cfg_w = ptw_io_requestor_1_pmp_0_cfg_w; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_0_cfg_r = ptw_io_requestor_1_pmp_0_cfg_r; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_0_addr = ptw_io_requestor_1_pmp_0_addr; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_0_mask = ptw_io_requestor_1_pmp_0_mask; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_1_cfg_l = ptw_io_requestor_1_pmp_1_cfg_l; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_1_cfg_a = ptw_io_requestor_1_pmp_1_cfg_a; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_1_cfg_x = ptw_io_requestor_1_pmp_1_cfg_x; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_1_cfg_w = ptw_io_requestor_1_pmp_1_cfg_w; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_1_cfg_r = ptw_io_requestor_1_pmp_1_cfg_r; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_1_addr = ptw_io_requestor_1_pmp_1_addr; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_1_mask = ptw_io_requestor_1_pmp_1_mask; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_2_cfg_l = ptw_io_requestor_1_pmp_2_cfg_l; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_2_cfg_a = ptw_io_requestor_1_pmp_2_cfg_a; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_2_cfg_x = ptw_io_requestor_1_pmp_2_cfg_x; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_2_cfg_w = ptw_io_requestor_1_pmp_2_cfg_w; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_2_cfg_r = ptw_io_requestor_1_pmp_2_cfg_r; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_2_addr = ptw_io_requestor_1_pmp_2_addr; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_2_mask = ptw_io_requestor_1_pmp_2_mask; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_3_cfg_l = ptw_io_requestor_1_pmp_3_cfg_l; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_3_cfg_a = ptw_io_requestor_1_pmp_3_cfg_a; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_3_cfg_x = ptw_io_requestor_1_pmp_3_cfg_x; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_3_cfg_w = ptw_io_requestor_1_pmp_3_cfg_w; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_3_cfg_r = ptw_io_requestor_1_pmp_3_cfg_r; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_3_addr = ptw_io_requestor_1_pmp_3_addr; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_3_mask = ptw_io_requestor_1_pmp_3_mask; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_4_cfg_l = ptw_io_requestor_1_pmp_4_cfg_l; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_4_cfg_a = ptw_io_requestor_1_pmp_4_cfg_a; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_4_cfg_x = ptw_io_requestor_1_pmp_4_cfg_x; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_4_cfg_w = ptw_io_requestor_1_pmp_4_cfg_w; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_4_cfg_r = ptw_io_requestor_1_pmp_4_cfg_r; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_4_addr = ptw_io_requestor_1_pmp_4_addr; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_4_mask = ptw_io_requestor_1_pmp_4_mask; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_5_cfg_l = ptw_io_requestor_1_pmp_5_cfg_l; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_5_cfg_a = ptw_io_requestor_1_pmp_5_cfg_a; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_5_cfg_x = ptw_io_requestor_1_pmp_5_cfg_x; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_5_cfg_w = ptw_io_requestor_1_pmp_5_cfg_w; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_5_cfg_r = ptw_io_requestor_1_pmp_5_cfg_r; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_5_addr = ptw_io_requestor_1_pmp_5_addr; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_5_mask = ptw_io_requestor_1_pmp_5_mask; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_6_cfg_l = ptw_io_requestor_1_pmp_6_cfg_l; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_6_cfg_a = ptw_io_requestor_1_pmp_6_cfg_a; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_6_cfg_x = ptw_io_requestor_1_pmp_6_cfg_x; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_6_cfg_w = ptw_io_requestor_1_pmp_6_cfg_w; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_6_cfg_r = ptw_io_requestor_1_pmp_6_cfg_r; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_6_addr = ptw_io_requestor_1_pmp_6_addr; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_6_mask = ptw_io_requestor_1_pmp_6_mask; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_7_cfg_l = ptw_io_requestor_1_pmp_7_cfg_l; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_7_cfg_a = ptw_io_requestor_1_pmp_7_cfg_a; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_7_cfg_x = ptw_io_requestor_1_pmp_7_cfg_x; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_7_cfg_w = ptw_io_requestor_1_pmp_7_cfg_w; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_7_cfg_r = ptw_io_requestor_1_pmp_7_cfg_r; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_7_addr = ptw_io_requestor_1_pmp_7_addr; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_pmp_7_mask = ptw_io_requestor_1_pmp_7_mask; // @[RocketTile.scala 198:20]
  assign frontend_io_ptw_customCSRs_csrs_0_value = ptw_io_requestor_1_customCSRs_csrs_0_value; // @[RocketTile.scala 198:20]
  assign fpuOpt_clock = clock;
  assign fpuOpt_reset = reset;
  assign fpuOpt_io_inst = core_io_fpu_inst; // @[RocketTile.scala 175:39]
  assign fpuOpt_io_fromint_data = core_io_fpu_fromint_data; // @[RocketTile.scala 175:39]
  assign fpuOpt_io_fcsr_rm = core_io_fpu_fcsr_rm; // @[RocketTile.scala 175:39]
  assign fpuOpt_io_dmem_resp_val = core_io_fpu_dmem_resp_val; // @[RocketTile.scala 175:39]
  assign fpuOpt_io_dmem_resp_type = core_io_fpu_dmem_resp_type; // @[RocketTile.scala 175:39]
  assign fpuOpt_io_dmem_resp_tag = core_io_fpu_dmem_resp_tag; // @[RocketTile.scala 175:39]
  assign fpuOpt_io_dmem_resp_data = core_io_fpu_dmem_resp_data; // @[RocketTile.scala 175:39]
  assign fpuOpt_io_valid = core_io_fpu_valid; // @[RocketTile.scala 175:39]
  assign fpuOpt_io_killx = core_io_fpu_killx; // @[RocketTile.scala 175:39]
  assign fpuOpt_io_killm = core_io_fpu_killm; // @[RocketTile.scala 175:39]
  assign dcacheArb_clock = clock;
  assign dcacheArb_io_requestor_0_req_valid = ptw_io_mem_req_valid; // @[RocketTile.scala 197:26]
  assign dcacheArb_io_requestor_0_req_bits_addr = ptw_io_mem_req_bits_addr; // @[RocketTile.scala 197:26]
  assign dcacheArb_io_requestor_0_s1_kill = ptw_io_mem_s1_kill; // @[RocketTile.scala 197:26]
  assign dcacheArb_io_requestor_1_req_valid = core_io_dmem_req_valid; // @[RocketTile.scala 197:26]
  assign dcacheArb_io_requestor_1_req_bits_addr = core_io_dmem_req_bits_addr; // @[RocketTile.scala 197:26]
  assign dcacheArb_io_requestor_1_req_bits_tag = core_io_dmem_req_bits_tag; // @[RocketTile.scala 197:26]
  assign dcacheArb_io_requestor_1_req_bits_cmd = core_io_dmem_req_bits_cmd; // @[RocketTile.scala 197:26]
  assign dcacheArb_io_requestor_1_req_bits_size = core_io_dmem_req_bits_size; // @[RocketTile.scala 197:26]
  assign dcacheArb_io_requestor_1_req_bits_signed = core_io_dmem_req_bits_signed; // @[RocketTile.scala 197:26]
  assign dcacheArb_io_requestor_1_s1_kill = core_io_dmem_s1_kill; // @[RocketTile.scala 197:26]
  assign dcacheArb_io_requestor_1_s1_data_data = core_io_dmem_s1_data_data; // @[RocketTile.scala 197:26]
  assign dcacheArb_io_mem_req_ready = dcache_io_cpu_req_ready; // @[HellaCache.scala 277:30]
  assign dcacheArb_io_mem_s2_nack = dcache_io_cpu_s2_nack; // @[HellaCache.scala 277:30]
  assign dcacheArb_io_mem_resp_valid = dcache_io_cpu_resp_valid; // @[HellaCache.scala 277:30]
  assign dcacheArb_io_mem_resp_bits_tag = dcache_io_cpu_resp_bits_tag; // @[HellaCache.scala 277:30]
  assign dcacheArb_io_mem_resp_bits_size = dcache_io_cpu_resp_bits_size; // @[HellaCache.scala 277:30]
  assign dcacheArb_io_mem_resp_bits_data = dcache_io_cpu_resp_bits_data; // @[HellaCache.scala 277:30]
  assign dcacheArb_io_mem_resp_bits_replay = dcache_io_cpu_resp_bits_replay; // @[HellaCache.scala 277:30]
  assign dcacheArb_io_mem_resp_bits_has_data = dcache_io_cpu_resp_bits_has_data; // @[HellaCache.scala 277:30]
  assign dcacheArb_io_mem_resp_bits_data_word_bypass = dcache_io_cpu_resp_bits_data_word_bypass; // @[HellaCache.scala 277:30]
  assign dcacheArb_io_mem_replay_next = dcache_io_cpu_replay_next; // @[HellaCache.scala 277:30]
  assign dcacheArb_io_mem_s2_xcpt_ma_ld = dcache_io_cpu_s2_xcpt_ma_ld; // @[HellaCache.scala 277:30]
  assign dcacheArb_io_mem_s2_xcpt_ma_st = dcache_io_cpu_s2_xcpt_ma_st; // @[HellaCache.scala 277:30]
  assign dcacheArb_io_mem_s2_xcpt_pf_ld = dcache_io_cpu_s2_xcpt_pf_ld; // @[HellaCache.scala 277:30]
  assign dcacheArb_io_mem_s2_xcpt_pf_st = dcache_io_cpu_s2_xcpt_pf_st; // @[HellaCache.scala 277:30]
  assign dcacheArb_io_mem_s2_xcpt_ae_ld = dcache_io_cpu_s2_xcpt_ae_ld; // @[HellaCache.scala 277:30]
  assign dcacheArb_io_mem_s2_xcpt_ae_st = dcache_io_cpu_s2_xcpt_ae_st; // @[HellaCache.scala 277:30]
  assign dcacheArb_io_mem_ordered = dcache_io_cpu_ordered; // @[HellaCache.scala 277:30]
  assign dcacheArb_io_mem_perf_release = dcache_io_cpu_perf_release; // @[HellaCache.scala 277:30]
  assign dcacheArb_io_mem_perf_grant = dcache_io_cpu_perf_grant; // @[HellaCache.scala 277:30]
  assign ptw_clock = clock;
  assign ptw_reset = reset;
  assign ptw_io_requestor_0_req_valid = dcache_io_ptw_req_valid; // @[RocketTile.scala 198:20]
  assign ptw_io_requestor_0_req_bits_bits_addr = dcache_io_ptw_req_bits_bits_addr; // @[RocketTile.scala 198:20]
  assign ptw_io_requestor_1_req_valid = frontend_io_ptw_req_valid; // @[RocketTile.scala 198:20]
  assign ptw_io_requestor_1_req_bits_valid = frontend_io_ptw_req_bits_valid; // @[RocketTile.scala 198:20]
  assign ptw_io_requestor_1_req_bits_bits_addr = frontend_io_ptw_req_bits_bits_addr; // @[RocketTile.scala 198:20]
  assign ptw_io_mem_req_ready = dcacheArb_io_requestor_0_req_ready; // @[RocketTile.scala 197:26]
  assign ptw_io_mem_s2_nack = dcacheArb_io_requestor_0_s2_nack; // @[RocketTile.scala 197:26]
  assign ptw_io_mem_resp_valid = dcacheArb_io_requestor_0_resp_valid; // @[RocketTile.scala 197:26]
  assign ptw_io_mem_resp_bits_data = dcacheArb_io_requestor_0_resp_bits_data; // @[RocketTile.scala 197:26]
  assign ptw_io_mem_s2_xcpt_ae_ld = dcacheArb_io_requestor_0_s2_xcpt_ae_ld; // @[RocketTile.scala 197:26]
  assign ptw_io_dpath_ptbr_mode = core_io_ptw_ptbr_mode; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_ptbr_ppn = core_io_ptw_ptbr_ppn; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_sfence_valid = core_io_ptw_sfence_valid; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_sfence_bits_rs1 = core_io_ptw_sfence_bits_rs1; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_status_debug = core_io_ptw_status_debug; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_status_dprv = core_io_ptw_status_dprv; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_status_prv = core_io_ptw_status_prv; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_status_mxr = core_io_ptw_status_mxr; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_status_sum = core_io_ptw_status_sum; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_0_cfg_l = core_io_ptw_pmp_0_cfg_l; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_0_cfg_a = core_io_ptw_pmp_0_cfg_a; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_0_cfg_x = core_io_ptw_pmp_0_cfg_x; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_0_cfg_w = core_io_ptw_pmp_0_cfg_w; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_0_cfg_r = core_io_ptw_pmp_0_cfg_r; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_0_addr = core_io_ptw_pmp_0_addr; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_0_mask = core_io_ptw_pmp_0_mask; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_1_cfg_l = core_io_ptw_pmp_1_cfg_l; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_1_cfg_a = core_io_ptw_pmp_1_cfg_a; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_1_cfg_x = core_io_ptw_pmp_1_cfg_x; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_1_cfg_w = core_io_ptw_pmp_1_cfg_w; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_1_cfg_r = core_io_ptw_pmp_1_cfg_r; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_1_addr = core_io_ptw_pmp_1_addr; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_1_mask = core_io_ptw_pmp_1_mask; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_2_cfg_l = core_io_ptw_pmp_2_cfg_l; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_2_cfg_a = core_io_ptw_pmp_2_cfg_a; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_2_cfg_x = core_io_ptw_pmp_2_cfg_x; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_2_cfg_w = core_io_ptw_pmp_2_cfg_w; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_2_cfg_r = core_io_ptw_pmp_2_cfg_r; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_2_addr = core_io_ptw_pmp_2_addr; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_2_mask = core_io_ptw_pmp_2_mask; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_3_cfg_l = core_io_ptw_pmp_3_cfg_l; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_3_cfg_a = core_io_ptw_pmp_3_cfg_a; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_3_cfg_x = core_io_ptw_pmp_3_cfg_x; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_3_cfg_w = core_io_ptw_pmp_3_cfg_w; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_3_cfg_r = core_io_ptw_pmp_3_cfg_r; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_3_addr = core_io_ptw_pmp_3_addr; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_3_mask = core_io_ptw_pmp_3_mask; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_4_cfg_l = core_io_ptw_pmp_4_cfg_l; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_4_cfg_a = core_io_ptw_pmp_4_cfg_a; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_4_cfg_x = core_io_ptw_pmp_4_cfg_x; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_4_cfg_w = core_io_ptw_pmp_4_cfg_w; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_4_cfg_r = core_io_ptw_pmp_4_cfg_r; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_4_addr = core_io_ptw_pmp_4_addr; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_4_mask = core_io_ptw_pmp_4_mask; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_5_cfg_l = core_io_ptw_pmp_5_cfg_l; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_5_cfg_a = core_io_ptw_pmp_5_cfg_a; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_5_cfg_x = core_io_ptw_pmp_5_cfg_x; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_5_cfg_w = core_io_ptw_pmp_5_cfg_w; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_5_cfg_r = core_io_ptw_pmp_5_cfg_r; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_5_addr = core_io_ptw_pmp_5_addr; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_5_mask = core_io_ptw_pmp_5_mask; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_6_cfg_l = core_io_ptw_pmp_6_cfg_l; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_6_cfg_a = core_io_ptw_pmp_6_cfg_a; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_6_cfg_x = core_io_ptw_pmp_6_cfg_x; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_6_cfg_w = core_io_ptw_pmp_6_cfg_w; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_6_cfg_r = core_io_ptw_pmp_6_cfg_r; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_6_addr = core_io_ptw_pmp_6_addr; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_6_mask = core_io_ptw_pmp_6_mask; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_7_cfg_l = core_io_ptw_pmp_7_cfg_l; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_7_cfg_a = core_io_ptw_pmp_7_cfg_a; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_7_cfg_x = core_io_ptw_pmp_7_cfg_x; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_7_cfg_w = core_io_ptw_pmp_7_cfg_w; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_7_cfg_r = core_io_ptw_pmp_7_cfg_r; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_7_addr = core_io_ptw_pmp_7_addr; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_pmp_7_mask = core_io_ptw_pmp_7_mask; // @[RocketTile.scala 176:15]
  assign ptw_io_dpath_customCSRs_csrs_0_value = core_io_ptw_customCSRs_csrs_0_value; // @[RocketTile.scala 176:15]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_hartid = broadcast_auto_out; // @[RocketTile.scala 168:18]
  assign core_io_interrupts_debug = intXbar_auto_int_out_0; // @[Interrupts.scala 85:93]
  assign core_io_interrupts_mtip = intXbar_auto_int_out_2; // @[Interrupts.scala 85:93]
  assign core_io_interrupts_msip = intXbar_auto_int_out_1; // @[Interrupts.scala 85:93]
  assign core_io_interrupts_meip = intXbar_auto_int_out_3; // @[Interrupts.scala 85:93]
  assign core_io_interrupts_seip = intXbar_auto_int_out_4; // @[Interrupts.scala 85:93]
  assign core_io_imem_resp_valid = frontend_io_cpu_resp_valid; // @[RocketTile.scala 173:32]
  assign core_io_imem_resp_bits_btb_taken = frontend_io_cpu_resp_bits_btb_taken; // @[RocketTile.scala 173:32]
  assign core_io_imem_resp_bits_btb_bridx = frontend_io_cpu_resp_bits_btb_bridx; // @[RocketTile.scala 173:32]
  assign core_io_imem_resp_bits_btb_entry = frontend_io_cpu_resp_bits_btb_entry; // @[RocketTile.scala 173:32]
  assign core_io_imem_resp_bits_btb_bht_history = frontend_io_cpu_resp_bits_btb_bht_history; // @[RocketTile.scala 173:32]
  assign core_io_imem_resp_bits_pc = frontend_io_cpu_resp_bits_pc; // @[RocketTile.scala 173:32]
  assign core_io_imem_resp_bits_data = frontend_io_cpu_resp_bits_data; // @[RocketTile.scala 173:32]
  assign core_io_imem_resp_bits_xcpt_pf_inst = frontend_io_cpu_resp_bits_xcpt_pf_inst; // @[RocketTile.scala 173:32]
  assign core_io_imem_resp_bits_xcpt_ae_inst = frontend_io_cpu_resp_bits_xcpt_ae_inst; // @[RocketTile.scala 173:32]
  assign core_io_imem_resp_bits_replay = frontend_io_cpu_resp_bits_replay; // @[RocketTile.scala 173:32]
  assign core_io_dmem_req_ready = dcacheArb_io_requestor_1_req_ready; // @[RocketTile.scala 197:26]
  assign core_io_dmem_s2_nack = dcacheArb_io_requestor_1_s2_nack; // @[RocketTile.scala 197:26]
  assign core_io_dmem_resp_valid = dcacheArb_io_requestor_1_resp_valid; // @[RocketTile.scala 197:26]
  assign core_io_dmem_resp_bits_tag = dcacheArb_io_requestor_1_resp_bits_tag; // @[RocketTile.scala 197:26]
  assign core_io_dmem_resp_bits_size = dcacheArb_io_requestor_1_resp_bits_size; // @[RocketTile.scala 197:26]
  assign core_io_dmem_resp_bits_data = dcacheArb_io_requestor_1_resp_bits_data; // @[RocketTile.scala 197:26]
  assign core_io_dmem_resp_bits_replay = dcacheArb_io_requestor_1_resp_bits_replay; // @[RocketTile.scala 197:26]
  assign core_io_dmem_resp_bits_has_data = dcacheArb_io_requestor_1_resp_bits_has_data; // @[RocketTile.scala 197:26]
  assign core_io_dmem_resp_bits_data_word_bypass = dcacheArb_io_requestor_1_resp_bits_data_word_bypass; // @[RocketTile.scala 197:26]
  assign core_io_dmem_replay_next = dcacheArb_io_requestor_1_replay_next; // @[RocketTile.scala 197:26]
  assign core_io_dmem_s2_xcpt_ma_ld = dcacheArb_io_requestor_1_s2_xcpt_ma_ld; // @[RocketTile.scala 197:26]
  assign core_io_dmem_s2_xcpt_ma_st = dcacheArb_io_requestor_1_s2_xcpt_ma_st; // @[RocketTile.scala 197:26]
  assign core_io_dmem_s2_xcpt_pf_ld = dcacheArb_io_requestor_1_s2_xcpt_pf_ld; // @[RocketTile.scala 197:26]
  assign core_io_dmem_s2_xcpt_pf_st = dcacheArb_io_requestor_1_s2_xcpt_pf_st; // @[RocketTile.scala 197:26]
  assign core_io_dmem_s2_xcpt_ae_ld = dcacheArb_io_requestor_1_s2_xcpt_ae_ld; // @[RocketTile.scala 197:26]
  assign core_io_dmem_s2_xcpt_ae_st = dcacheArb_io_requestor_1_s2_xcpt_ae_st; // @[RocketTile.scala 197:26]
  assign core_io_dmem_ordered = dcacheArb_io_requestor_1_ordered; // @[RocketTile.scala 197:26]
  assign core_io_dmem_perf_release = dcacheArb_io_requestor_1_perf_release; // @[RocketTile.scala 197:26]
  assign core_io_dmem_perf_grant = dcacheArb_io_requestor_1_perf_grant; // @[RocketTile.scala 197:26]
  assign core_io_fpu_fcsr_flags_valid = fpuOpt_io_fcsr_flags_valid; // @[RocketTile.scala 175:39]
  assign core_io_fpu_fcsr_flags_bits = fpuOpt_io_fcsr_flags_bits; // @[RocketTile.scala 175:39]
  assign core_io_fpu_store_data = fpuOpt_io_store_data; // @[RocketTile.scala 175:39]
  assign core_io_fpu_toint_data = fpuOpt_io_toint_data; // @[RocketTile.scala 175:39]
  assign core_io_fpu_fcsr_rdy = fpuOpt_io_fcsr_rdy; // @[RocketTile.scala 175:39]
  assign core_io_fpu_nack_mem = fpuOpt_io_nack_mem; // @[RocketTile.scala 175:39]
  assign core_io_fpu_illegal_rm = fpuOpt_io_illegal_rm; // @[RocketTile.scala 175:39]
  assign core_io_fpu_dec_wen = fpuOpt_io_dec_wen; // @[RocketTile.scala 175:39]
  assign core_io_fpu_dec_ren1 = fpuOpt_io_dec_ren1; // @[RocketTile.scala 175:39]
  assign core_io_fpu_dec_ren2 = fpuOpt_io_dec_ren2; // @[RocketTile.scala 175:39]
  assign core_io_fpu_dec_ren3 = fpuOpt_io_dec_ren3; // @[RocketTile.scala 175:39]
  assign core_io_fpu_sboard_set = fpuOpt_io_sboard_set; // @[RocketTile.scala 175:39]
  assign core_io_fpu_sboard_clr = fpuOpt_io_sboard_clr; // @[RocketTile.scala 175:39]
  assign core_io_fpu_sboard_clra = fpuOpt_io_sboard_clra; // @[RocketTile.scala 175:39]
  assign RocketTile_covSum = 30'h0;
  assign tlMasterXbar_sum = RocketTile_covSum + tlMasterXbar_io_covSum;
  assign intXbar_sum = tlMasterXbar_sum + intXbar_io_covSum;
  assign fpuOpt_sum = intXbar_sum + fpuOpt_io_covSum;
  assign dcacheArb_sum = fpuOpt_sum + dcacheArb_io_covSum;
  assign frontend_sum = dcacheArb_sum + frontend_io_covSum;
  assign dcache_sum = frontend_sum + dcache_io_covSum;
  assign broadcast_3_sum = dcache_sum + broadcast_3_io_covSum;
  assign core_sum = broadcast_3_sum + core_io_covSum;
  assign broadcast_sum = core_sum + broadcast_io_covSum;
  assign broadcast_1_sum = broadcast_sum + broadcast_1_io_covSum;
  assign ptw_sum = broadcast_1_sum + ptw_io_covSum;
  assign io_covSum = ptw_sum;
  assign broadcast_1_metaAssert_wire = broadcast_1_metaAssert;
  assign core_metaAssert_wire = core_metaAssert;
  assign broadcast_metaAssert_wire = broadcast_metaAssert;
  assign dcache_metaAssert_wire = dcache_metaAssert;
  assign intXbar_metaAssert_wire = intXbar_metaAssert;
  assign tlMasterXbar_metaAssert_wire = tlMasterXbar_metaAssert;
  assign broadcast_3_metaAssert_wire = broadcast_3_metaAssert;
  assign frontend_metaAssert_wire = frontend_metaAssert;
  assign dcacheArb_metaAssert_wire = dcacheArb_metaAssert;
  assign fpuOpt_metaAssert_wire = fpuOpt_metaAssert;
  assign ptw_metaAssert_wire = ptw_metaAssert;
  assign RocketTile_or3 = tlMasterXbar_metaAssert_wire | broadcast_3_metaAssert_wire;
  assign RocketTile_or10 = dcache_metaAssert_wire | fpuOpt_metaAssert_wire;
  assign RocketTile_or4 = frontend_metaAssert_wire | RocketTile_or10;
  assign RocketTile_or1 = RocketTile_or3 | RocketTile_or4;
  assign RocketTile_or12 = intXbar_metaAssert_wire | ptw_metaAssert_wire;
  assign RocketTile_or5 = broadcast_1_metaAssert_wire | RocketTile_or12;
  assign RocketTile_or14 = core_metaAssert_wire | dcacheArb_metaAssert_wire;
  assign RocketTile_or6 = broadcast_metaAssert_wire | RocketTile_or14;
  assign RocketTile_or2 = RocketTile_or5 | RocketTile_or6;
  assign RocketTile_or0 = RocketTile_or1 | RocketTile_or2;
  assign metaAssert = RocketTile_metaAssert;
  assign tlMasterXbar_metaReset = metaReset | tlMasterXbar_halt;
  assign fpuOpt_metaReset = metaReset | fpuOpt_halt;
  assign dcacheArb_metaReset = metaReset | dcacheArb_halt;
  assign frontend_metaReset = metaReset | frontend_halt;
  assign dcache_metaReset = metaReset | dcache_halt;
  assign core_metaReset = metaReset | core_halt;
  assign ptw_metaReset = metaReset | ptw_halt;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  bundleOut_0_0_REG = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  RocketTile_metaAssert = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      bundleOut_0_0_REG <= 1'h0;
    end else if (reset) begin
      bundleOut_0_0_REG <= 1'h0;
    end else begin
      bundleOut_0_0_REG <= core_io_wfi;
    end
    if (metaReset) begin
      RocketTile_metaAssert <= 1'h0;
    end else begin
      RocketTile_metaAssert <= RocketTile_metaAssert | RocketTile_or0;
    end
  end
endmodule
module TLXbar_7(
  input         clock,
  input         reset,
  output        auto_in_1_a_ready,
  input         auto_in_1_a_valid,
  input  [31:0] auto_in_1_a_bits_address,
  output        auto_in_1_d_valid,
  output [2:0]  auto_in_1_d_bits_opcode,
  output [3:0]  auto_in_1_d_bits_size,
  output [63:0] auto_in_1_d_bits_data,
  output        auto_in_1_d_bits_corrupt,
  output        auto_in_0_a_ready,
  input         auto_in_0_a_valid,
  input  [2:0]  auto_in_0_a_bits_opcode,
  input  [2:0]  auto_in_0_a_bits_param,
  input  [3:0]  auto_in_0_a_bits_size,
  input         auto_in_0_a_bits_source,
  input  [31:0] auto_in_0_a_bits_address,
  input  [7:0]  auto_in_0_a_bits_mask,
  input  [63:0] auto_in_0_a_bits_data,
  input         auto_in_0_b_ready,
  output        auto_in_0_b_valid,
  output [1:0]  auto_in_0_b_bits_param,
  output [3:0]  auto_in_0_b_bits_size,
  output        auto_in_0_b_bits_source,
  output [31:0] auto_in_0_b_bits_address,
  output        auto_in_0_c_ready,
  input         auto_in_0_c_valid,
  input  [2:0]  auto_in_0_c_bits_opcode,
  input  [2:0]  auto_in_0_c_bits_param,
  input  [3:0]  auto_in_0_c_bits_size,
  input         auto_in_0_c_bits_source,
  input  [31:0] auto_in_0_c_bits_address,
  input  [63:0] auto_in_0_c_bits_data,
  input         auto_in_0_d_ready,
  output        auto_in_0_d_valid,
  output [2:0]  auto_in_0_d_bits_opcode,
  output [1:0]  auto_in_0_d_bits_param,
  output [3:0]  auto_in_0_d_bits_size,
  output        auto_in_0_d_bits_source,
  output [1:0]  auto_in_0_d_bits_sink,
  output        auto_in_0_d_bits_denied,
  output [63:0] auto_in_0_d_bits_data,
  output        auto_in_0_e_ready,
  input         auto_in_0_e_valid,
  input  [1:0]  auto_in_0_e_bits_sink,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_opcode,
  output [2:0]  auto_out_a_bits_param,
  output [3:0]  auto_out_a_bits_size,
  output [1:0]  auto_out_a_bits_source,
  output [31:0] auto_out_a_bits_address,
  output [7:0]  auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input  [2:0]  auto_out_b_bits_opcode,
  input  [1:0]  auto_out_b_bits_param,
  input  [3:0]  auto_out_b_bits_size,
  input  [1:0]  auto_out_b_bits_source,
  input  [31:0] auto_out_b_bits_address,
  input  [7:0]  auto_out_b_bits_mask,
  input         auto_out_b_bits_corrupt,
  input         auto_out_c_ready,
  output        auto_out_c_valid,
  output [2:0]  auto_out_c_bits_opcode,
  output [2:0]  auto_out_c_bits_param,
  output [3:0]  auto_out_c_bits_size,
  output [1:0]  auto_out_c_bits_source,
  output [31:0] auto_out_c_bits_address,
  output [63:0] auto_out_c_bits_data,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [2:0]  auto_out_d_bits_opcode,
  input  [1:0]  auto_out_d_bits_param,
  input  [3:0]  auto_out_d_bits_size,
  input  [1:0]  auto_out_d_bits_source,
  input  [1:0]  auto_out_d_bits_sink,
  input         auto_out_d_bits_denied,
  input  [63:0] auto_out_d_bits_data,
  input         auto_out_d_bits_corrupt,
  input         auto_out_e_ready,
  output        auto_out_e_valid,
  output [1:0]  auto_out_e_bits_sink,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset,
  input         monitor_halt,
  input         monitor_1_halt
);
  wire  monitor_clock; // @[Nodes.scala 24:25]
  wire  monitor_reset; // @[Nodes.scala 24:25]
  wire  monitor_io_in_a_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_a_valid; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_a_bits_opcode; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_a_bits_param; // @[Nodes.scala 24:25]
  wire [3:0] monitor_io_in_a_bits_size; // @[Nodes.scala 24:25]
  wire  monitor_io_in_a_bits_source; // @[Nodes.scala 24:25]
  wire [31:0] monitor_io_in_a_bits_address; // @[Nodes.scala 24:25]
  wire [7:0] monitor_io_in_a_bits_mask; // @[Nodes.scala 24:25]
  wire  monitor_io_in_b_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_b_valid; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_b_bits_opcode; // @[Nodes.scala 24:25]
  wire [1:0] monitor_io_in_b_bits_param; // @[Nodes.scala 24:25]
  wire [3:0] monitor_io_in_b_bits_size; // @[Nodes.scala 24:25]
  wire  monitor_io_in_b_bits_source; // @[Nodes.scala 24:25]
  wire [31:0] monitor_io_in_b_bits_address; // @[Nodes.scala 24:25]
  wire [7:0] monitor_io_in_b_bits_mask; // @[Nodes.scala 24:25]
  wire  monitor_io_in_b_bits_corrupt; // @[Nodes.scala 24:25]
  wire  monitor_io_in_c_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_c_valid; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_c_bits_opcode; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_c_bits_param; // @[Nodes.scala 24:25]
  wire [3:0] monitor_io_in_c_bits_size; // @[Nodes.scala 24:25]
  wire  monitor_io_in_c_bits_source; // @[Nodes.scala 24:25]
  wire [31:0] monitor_io_in_c_bits_address; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_valid; // @[Nodes.scala 24:25]
  wire [2:0] monitor_io_in_d_bits_opcode; // @[Nodes.scala 24:25]
  wire [1:0] monitor_io_in_d_bits_param; // @[Nodes.scala 24:25]
  wire [3:0] monitor_io_in_d_bits_size; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_bits_source; // @[Nodes.scala 24:25]
  wire [1:0] monitor_io_in_d_bits_sink; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_bits_denied; // @[Nodes.scala 24:25]
  wire  monitor_io_in_d_bits_corrupt; // @[Nodes.scala 24:25]
  wire  monitor_io_in_e_ready; // @[Nodes.scala 24:25]
  wire  monitor_io_in_e_valid; // @[Nodes.scala 24:25]
  wire [1:0] monitor_io_in_e_bits_sink; // @[Nodes.scala 24:25]
  wire [29:0] monitor_io_covSum; // @[Nodes.scala 24:25]
  wire  monitor_metaAssert; // @[Nodes.scala 24:25]
  wire  monitor_metaReset; // @[Nodes.scala 24:25]
  wire  monitor_1_clock; // @[Nodes.scala 24:25]
  wire  monitor_1_reset; // @[Nodes.scala 24:25]
  wire  monitor_1_io_in_a_ready; // @[Nodes.scala 24:25]
  wire  monitor_1_io_in_a_valid; // @[Nodes.scala 24:25]
  wire [31:0] monitor_1_io_in_a_bits_address; // @[Nodes.scala 24:25]
  wire  monitor_1_io_in_d_valid; // @[Nodes.scala 24:25]
  wire [2:0] monitor_1_io_in_d_bits_opcode; // @[Nodes.scala 24:25]
  wire [1:0] monitor_1_io_in_d_bits_param; // @[Nodes.scala 24:25]
  wire [3:0] monitor_1_io_in_d_bits_size; // @[Nodes.scala 24:25]
  wire [1:0] monitor_1_io_in_d_bits_sink; // @[Nodes.scala 24:25]
  wire  monitor_1_io_in_d_bits_denied; // @[Nodes.scala 24:25]
  wire  monitor_1_io_in_d_bits_corrupt; // @[Nodes.scala 24:25]
  wire [29:0] monitor_1_io_covSum; // @[Nodes.scala 24:25]
  wire  monitor_1_metaAssert; // @[Nodes.scala 24:25]
  wire  monitor_1_metaReset; // @[Nodes.scala 24:25]
  wire  requestBOI_0_0; // @[Parameters.scala 54:32]
  wire  requestDOI_0_0; // @[Parameters.scala 54:32]
  wire  requestDOI_0_1; // @[Parameters.scala 46:9]
  wire [26:0] _beatsAI_decode_T_1; // @[package.scala 234:77]
  wire [8:0] beatsAI_decode; // @[Edges.scala 219:59]
  wire  beatsAI_opdata; // @[Edges.scala 91:28]
  wire  _portsDIO_out_0_d_ready_T; // @[Mux.scala 27:72]
  reg [8:0] beatsLeft; // @[Arbiter.scala 87:30]
  reg [31:0] _RAND_0;
  wire  idle; // @[Arbiter.scala 88:28]
  wire  latch; // @[Arbiter.scala 89:24]
  wire [1:0] readys_filter_lo; // @[Cat.scala 30:58]
  wire  _readys_T_1; // @[Arbiter.scala 22:19]
  wire  _readys_T_3; // @[Arbiter.scala 22:12]
  reg [1:0] readys_mask; // @[Arbiter.scala 23:23]
  reg [31:0] _RAND_1;
  wire [1:0] readys_filter_hi; // @[Arbiter.scala 24:28]
  wire [3:0] readys_filter; // @[Cat.scala 30:58]
  wire [3:0] _GEN_1; // @[package.scala 253:43]
  wire [3:0] _readys_unready_T_1; // @[package.scala 253:43]
  wire [3:0] _readys_unready_T_4; // @[Arbiter.scala 25:66]
  wire [3:0] _GEN_2; // @[Arbiter.scala 25:58]
  wire [3:0] readys_unready; // @[Arbiter.scala 25:58]
  wire [1:0] _readys_readys_T_2; // @[Arbiter.scala 26:39]
  wire [1:0] readys_readys; // @[Arbiter.scala 26:18]
  wire  _readys_T_5; // @[Arbiter.scala 27:27]
  wire  _readys_T_6; // @[Arbiter.scala 27:18]
  wire [1:0] _readys_mask_T; // @[Arbiter.scala 28:29]
  wire [2:0] _readys_mask_T_1; // @[package.scala 244:48]
  wire [1:0] _readys_mask_T_3; // @[package.scala 244:43]
  wire  readys_0; // @[Arbiter.scala 95:86]
  wire  readys_1; // @[Arbiter.scala 95:86]
  wire  earlyWinner_0; // @[Arbiter.scala 97:79]
  wire  earlyWinner_1; // @[Arbiter.scala 97:79]
  wire  _prefixOR_T; // @[Arbiter.scala 104:53]
  wire  _T_6; // @[Arbiter.scala 105:64]
  wire  _T_9; // @[Arbiter.scala 105:13]
  wire  _T_11; // @[Arbiter.scala 107:36]
  wire  _T_14; // @[Arbiter.scala 107:41]
  wire  _T_16; // @[Arbiter.scala 107:14]
  wire  _T_21; // @[Arbiter.scala 108:41]
  wire  _T_23; // @[Arbiter.scala 108:14]
  reg  state_0; // @[Arbiter.scala 116:26]
  reg [31:0] _RAND_2;
  wire  muxStateEarly_0; // @[Arbiter.scala 117:30]
  reg  state_1; // @[Arbiter.scala 116:26]
  reg [31:0] _RAND_3;
  wire  muxStateEarly_1; // @[Arbiter.scala 117:30]
  wire  _out_0_a_earlyValid_T_1; // @[Mux.scala 27:72]
  wire  _out_0_a_earlyValid_T_2; // @[Mux.scala 27:72]
  wire  _out_0_a_earlyValid_T_3; // @[Mux.scala 27:72]
  wire  out_2_0_a_earlyValid; // @[Arbiter.scala 125:29]
  wire  _beatsLeft_T_2; // @[ReadyValidCancel.scala 50:33]
  wire [8:0] _GEN_3; // @[Arbiter.scala 113:52]
  wire [8:0] _beatsLeft_T_4; // @[Arbiter.scala 113:52]
  wire  allowed_0; // @[Arbiter.scala 121:24]
  wire  allowed_1; // @[Arbiter.scala 121:24]
  wire [7:0] _T_31; // @[Mux.scala 27:72]
  wire [7:0] _T_32; // @[Mux.scala 27:72]
  wire [31:0] _T_34; // @[Mux.scala 27:72]
  wire [31:0] _T_35; // @[Mux.scala 27:72]
  wire [1:0] in_0_a_bits_source; // @[Xbar.scala 231:18 BundleMap.scala 247:19 Xbar.scala 237:29]
  wire [1:0] _T_37; // @[Mux.scala 27:72]
  wire [1:0] _T_38; // @[Mux.scala 27:72]
  wire [3:0] _T_40; // @[Mux.scala 27:72]
  wire [3:0] _T_41; // @[Mux.scala 27:72]
  wire [2:0] _T_46; // @[Mux.scala 27:72]
  wire [2:0] _T_47; // @[Mux.scala 27:72]
  reg [2:0] TLXbar_7_state; // @[Register tracking TLXbar_7 state]
  reg [31:0] _RAND_4;
  reg  TLXbar_7_cov [0:7]; // @[Coverage map for TLXbar_7]
  reg [31:0] _RAND_5;
  wire  TLXbar_7_cov_read_data; // @[Coverage map for TLXbar_7]
  wire [2:0] TLXbar_7_cov_read_addr; // @[Coverage map for TLXbar_7]
  wire  TLXbar_7_cov_write_data; // @[Coverage map for TLXbar_7]
  wire [2:0] TLXbar_7_cov_write_addr; // @[Coverage map for TLXbar_7]
  wire  TLXbar_7_cov_write_mask; // @[Coverage map for TLXbar_7]
  wire  TLXbar_7_cov_write_en; // @[Coverage map for TLXbar_7]
  reg [29:0] TLXbar_7_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_6;
  wire [1:0] readys_mask_shl;
  wire [2:0] readys_mask_pad;
  wire [2:0] state_0_shl;
  wire [2:0] state_0_pad;
  wire [2:0] state_1_shl;
  wire [2:0] state_1_pad;
  wire [2:0] TLXbar_7_xor2;
  wire [2:0] TLXbar_7_xor0;
  wire [29:0] monitor_sum;
  wire [29:0] monitor_1_sum;
  wire  stopEn0;
  wire  stopEn1;
  wire  stopEn2;
  wire  stopEn3;
  wire  monitor_metaAssert_wire;
  wire  monitor_1_metaAssert_wire;
  wire  TLXbar_7_or4;
  wire  TLXbar_7_or1;
  wire  TLXbar_7_or6;
  wire  TLXbar_7_or2;
  wire  TLXbar_7_or0;
  reg  TLXbar_7_metaAssert;
  reg [31:0] _RAND_7;
  TLMonitor_23 monitor ( // @[Nodes.scala 24:25]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_a_ready(monitor_io_in_a_ready),
    .io_in_a_valid(monitor_io_in_a_valid),
    .io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(monitor_io_in_a_bits_param),
    .io_in_a_bits_size(monitor_io_in_a_bits_size),
    .io_in_a_bits_source(monitor_io_in_a_bits_source),
    .io_in_a_bits_address(monitor_io_in_a_bits_address),
    .io_in_a_bits_mask(monitor_io_in_a_bits_mask),
    .io_in_b_ready(monitor_io_in_b_ready),
    .io_in_b_valid(monitor_io_in_b_valid),
    .io_in_b_bits_opcode(monitor_io_in_b_bits_opcode),
    .io_in_b_bits_param(monitor_io_in_b_bits_param),
    .io_in_b_bits_size(monitor_io_in_b_bits_size),
    .io_in_b_bits_source(monitor_io_in_b_bits_source),
    .io_in_b_bits_address(monitor_io_in_b_bits_address),
    .io_in_b_bits_mask(monitor_io_in_b_bits_mask),
    .io_in_b_bits_corrupt(monitor_io_in_b_bits_corrupt),
    .io_in_c_ready(monitor_io_in_c_ready),
    .io_in_c_valid(monitor_io_in_c_valid),
    .io_in_c_bits_opcode(monitor_io_in_c_bits_opcode),
    .io_in_c_bits_param(monitor_io_in_c_bits_param),
    .io_in_c_bits_size(monitor_io_in_c_bits_size),
    .io_in_c_bits_source(monitor_io_in_c_bits_source),
    .io_in_c_bits_address(monitor_io_in_c_bits_address),
    .io_in_d_ready(monitor_io_in_d_ready),
    .io_in_d_valid(monitor_io_in_d_valid),
    .io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(monitor_io_in_d_bits_param),
    .io_in_d_bits_size(monitor_io_in_d_bits_size),
    .io_in_d_bits_source(monitor_io_in_d_bits_source),
    .io_in_d_bits_sink(monitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(monitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt),
    .io_in_e_ready(monitor_io_in_e_ready),
    .io_in_e_valid(monitor_io_in_e_valid),
    .io_in_e_bits_sink(monitor_io_in_e_bits_sink),
    .io_covSum(monitor_io_covSum),
    .metaAssert(monitor_metaAssert),
    .metaReset(monitor_metaReset)
  );
  TLMonitor_24 monitor_1 ( // @[Nodes.scala 24:25]
    .clock(monitor_1_clock),
    .reset(monitor_1_reset),
    .io_in_a_ready(monitor_1_io_in_a_ready),
    .io_in_a_valid(monitor_1_io_in_a_valid),
    .io_in_a_bits_address(monitor_1_io_in_a_bits_address),
    .io_in_d_valid(monitor_1_io_in_d_valid),
    .io_in_d_bits_opcode(monitor_1_io_in_d_bits_opcode),
    .io_in_d_bits_param(monitor_1_io_in_d_bits_param),
    .io_in_d_bits_size(monitor_1_io_in_d_bits_size),
    .io_in_d_bits_sink(monitor_1_io_in_d_bits_sink),
    .io_in_d_bits_denied(monitor_1_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(monitor_1_io_in_d_bits_corrupt),
    .io_covSum(monitor_1_io_covSum),
    .metaAssert(monitor_1_metaAssert),
    .metaReset(monitor_1_metaReset)
  );
  assign requestBOI_0_0 = ~auto_out_b_bits_source[1]; // @[Parameters.scala 54:32]
  assign requestDOI_0_0 = ~auto_out_d_bits_source[1]; // @[Parameters.scala 54:32]
  assign requestDOI_0_1 = auto_out_d_bits_source == 2'h2; // @[Parameters.scala 46:9]
  assign _beatsAI_decode_T_1 = 27'hfff << auto_in_0_a_bits_size; // @[package.scala 234:77]
  assign beatsAI_decode = ~_beatsAI_decode_T_1[11:3]; // @[Edges.scala 219:59]
  assign beatsAI_opdata = ~auto_in_0_a_bits_opcode[2]; // @[Edges.scala 91:28]
  assign _portsDIO_out_0_d_ready_T = requestDOI_0_0 & auto_in_0_d_ready; // @[Mux.scala 27:72]
  assign idle = beatsLeft == 9'h0; // @[Arbiter.scala 88:28]
  assign latch = idle & auto_out_a_ready; // @[Arbiter.scala 89:24]
  assign readys_filter_lo = {auto_in_1_a_valid,auto_in_0_a_valid}; // @[Cat.scala 30:58]
  assign _readys_T_1 = readys_filter_lo == readys_filter_lo; // @[Arbiter.scala 22:19]
  assign _readys_T_3 = _readys_T_1 | reset; // @[Arbiter.scala 22:12]
  assign readys_filter_hi = readys_filter_lo & ~readys_mask; // @[Arbiter.scala 24:28]
  assign readys_filter = {readys_filter_hi,auto_in_1_a_valid,auto_in_0_a_valid}; // @[Cat.scala 30:58]
  assign _GEN_1 = {{1'd0}, readys_filter[3:1]}; // @[package.scala 253:43]
  assign _readys_unready_T_1 = readys_filter | _GEN_1; // @[package.scala 253:43]
  assign _readys_unready_T_4 = {readys_mask, 2'h0}; // @[Arbiter.scala 25:66]
  assign _GEN_2 = {{1'd0}, _readys_unready_T_1[3:1]}; // @[Arbiter.scala 25:58]
  assign readys_unready = _GEN_2 | _readys_unready_T_4; // @[Arbiter.scala 25:58]
  assign _readys_readys_T_2 = readys_unready[3:2] & readys_unready[1:0]; // @[Arbiter.scala 26:39]
  assign readys_readys = ~_readys_readys_T_2; // @[Arbiter.scala 26:18]
  assign _readys_T_5 = |readys_filter_lo; // @[Arbiter.scala 27:27]
  assign _readys_T_6 = latch & _readys_T_5; // @[Arbiter.scala 27:18]
  assign _readys_mask_T = readys_readys & readys_filter_lo; // @[Arbiter.scala 28:29]
  assign _readys_mask_T_1 = {_readys_mask_T, 1'h0}; // @[package.scala 244:48]
  assign _readys_mask_T_3 = _readys_mask_T | _readys_mask_T_1[1:0]; // @[package.scala 244:43]
  assign readys_0 = readys_readys[0]; // @[Arbiter.scala 95:86]
  assign readys_1 = readys_readys[1]; // @[Arbiter.scala 95:86]
  assign earlyWinner_0 = readys_0 & auto_in_0_a_valid; // @[Arbiter.scala 97:79]
  assign earlyWinner_1 = readys_1 & auto_in_1_a_valid; // @[Arbiter.scala 97:79]
  assign _prefixOR_T = earlyWinner_0 | earlyWinner_1; // @[Arbiter.scala 104:53]
  assign _T_6 = ~earlyWinner_0 | ~earlyWinner_1; // @[Arbiter.scala 105:64]
  assign _T_9 = _T_6 | reset; // @[Arbiter.scala 105:13]
  assign _T_11 = auto_in_0_a_valid | auto_in_1_a_valid; // @[Arbiter.scala 107:36]
  assign _T_14 = ~_T_11 | _prefixOR_T; // @[Arbiter.scala 107:41]
  assign _T_16 = _T_14 | reset; // @[Arbiter.scala 107:14]
  assign _T_21 = ~_T_11 | _T_11; // @[Arbiter.scala 108:41]
  assign _T_23 = _T_21 | reset; // @[Arbiter.scala 108:14]
  assign muxStateEarly_0 = idle ? earlyWinner_0 : state_0; // @[Arbiter.scala 117:30]
  assign muxStateEarly_1 = idle ? earlyWinner_1 : state_1; // @[Arbiter.scala 117:30]
  assign _out_0_a_earlyValid_T_1 = state_0 & auto_in_0_a_valid; // @[Mux.scala 27:72]
  assign _out_0_a_earlyValid_T_2 = state_1 & auto_in_1_a_valid; // @[Mux.scala 27:72]
  assign _out_0_a_earlyValid_T_3 = _out_0_a_earlyValid_T_1 | _out_0_a_earlyValid_T_2; // @[Mux.scala 27:72]
  assign out_2_0_a_earlyValid = idle ? _T_11 : _out_0_a_earlyValid_T_3; // @[Arbiter.scala 125:29]
  assign _beatsLeft_T_2 = auto_out_a_ready & out_2_0_a_earlyValid; // @[ReadyValidCancel.scala 50:33]
  assign _GEN_3 = {{8'd0}, _beatsLeft_T_2}; // @[Arbiter.scala 113:52]
  assign _beatsLeft_T_4 = beatsLeft - _GEN_3; // @[Arbiter.scala 113:52]
  assign allowed_0 = idle ? readys_0 : state_0; // @[Arbiter.scala 121:24]
  assign allowed_1 = idle ? readys_1 : state_1; // @[Arbiter.scala 121:24]
  assign _T_31 = muxStateEarly_0 ? auto_in_0_a_bits_mask : 8'h0; // @[Mux.scala 27:72]
  assign _T_32 = muxStateEarly_1 ? 8'hff : 8'h0; // @[Mux.scala 27:72]
  assign _T_34 = muxStateEarly_0 ? auto_in_0_a_bits_address : 32'h0; // @[Mux.scala 27:72]
  assign _T_35 = muxStateEarly_1 ? auto_in_1_a_bits_address : 32'h0; // @[Mux.scala 27:72]
  assign in_0_a_bits_source = {{1'd0}, auto_in_0_a_bits_source}; // @[Xbar.scala 231:18 BundleMap.scala 247:19 Xbar.scala 237:29]
  assign _T_37 = muxStateEarly_0 ? in_0_a_bits_source : 2'h0; // @[Mux.scala 27:72]
  assign _T_38 = muxStateEarly_1 ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  assign _T_40 = muxStateEarly_0 ? auto_in_0_a_bits_size : 4'h0; // @[Mux.scala 27:72]
  assign _T_41 = muxStateEarly_1 ? 4'h6 : 4'h0; // @[Mux.scala 27:72]
  assign _T_46 = muxStateEarly_0 ? auto_in_0_a_bits_opcode : 3'h0; // @[Mux.scala 27:72]
  assign _T_47 = muxStateEarly_1 ? 3'h4 : 3'h0; // @[Mux.scala 27:72]
  assign auto_in_1_a_ready = auto_out_a_ready & allowed_1; // @[LazyModule.scala 309:16]
  assign auto_in_1_d_valid = auto_out_d_valid & requestDOI_0_1; // @[LazyModule.scala 309:16]
  assign auto_in_1_d_bits_opcode = auto_out_d_bits_opcode; // @[LazyModule.scala 309:16]
  assign auto_in_1_d_bits_size = auto_out_d_bits_size; // @[LazyModule.scala 309:16]
  assign auto_in_1_d_bits_data = auto_out_d_bits_data; // @[LazyModule.scala 309:16]
  assign auto_in_1_d_bits_corrupt = auto_out_d_bits_corrupt; // @[LazyModule.scala 309:16]
  assign auto_in_0_a_ready = auto_out_a_ready & allowed_0; // @[LazyModule.scala 309:16]
  assign auto_in_0_b_valid = auto_out_b_valid & requestBOI_0_0; // @[LazyModule.scala 309:16]
  assign auto_in_0_b_bits_param = auto_out_b_bits_param; // @[LazyModule.scala 309:16]
  assign auto_in_0_b_bits_size = auto_out_b_bits_size; // @[LazyModule.scala 309:16]
  assign auto_in_0_b_bits_source = auto_out_b_bits_source[0]; // @[LazyModule.scala 309:16]
  assign auto_in_0_b_bits_address = auto_out_b_bits_address; // @[LazyModule.scala 309:16]
  assign auto_in_0_c_ready = auto_out_c_ready; // @[LazyModule.scala 309:16]
  assign auto_in_0_d_valid = auto_out_d_valid & requestDOI_0_0; // @[LazyModule.scala 309:16]
  assign auto_in_0_d_bits_opcode = auto_out_d_bits_opcode; // @[LazyModule.scala 309:16]
  assign auto_in_0_d_bits_param = auto_out_d_bits_param; // @[LazyModule.scala 309:16]
  assign auto_in_0_d_bits_size = auto_out_d_bits_size; // @[LazyModule.scala 309:16]
  assign auto_in_0_d_bits_source = auto_out_d_bits_source[0]; // @[LazyModule.scala 309:16]
  assign auto_in_0_d_bits_sink = auto_out_d_bits_sink; // @[LazyModule.scala 309:16]
  assign auto_in_0_d_bits_denied = auto_out_d_bits_denied; // @[LazyModule.scala 309:16]
  assign auto_in_0_d_bits_data = auto_out_d_bits_data; // @[LazyModule.scala 309:16]
  assign auto_in_0_e_ready = auto_out_e_ready; // @[LazyModule.scala 309:16]
  assign auto_out_a_valid = idle ? _T_11 : _out_0_a_earlyValid_T_3; // @[LazyModule.scala 311:12]
  assign auto_out_a_bits_opcode = _T_46 | _T_47; // @[LazyModule.scala 311:12]
  assign auto_out_a_bits_param = muxStateEarly_0 ? auto_in_0_a_bits_param : 3'h0; // @[LazyModule.scala 311:12]
  assign auto_out_a_bits_size = _T_40 | _T_41; // @[LazyModule.scala 311:12]
  assign auto_out_a_bits_source = _T_37 | _T_38; // @[LazyModule.scala 311:12]
  assign auto_out_a_bits_address = _T_34 | _T_35; // @[LazyModule.scala 311:12]
  assign auto_out_a_bits_mask = _T_31 | _T_32; // @[LazyModule.scala 311:12]
  assign auto_out_a_bits_data = muxStateEarly_0 ? auto_in_0_a_bits_data : 64'h0; // @[LazyModule.scala 311:12]
  assign auto_out_b_ready = requestBOI_0_0 & auto_in_0_b_ready; // @[LazyModule.scala 311:12]
  assign auto_out_c_valid = auto_in_0_c_valid; // @[LazyModule.scala 311:12]
  assign auto_out_c_bits_opcode = auto_in_0_c_bits_opcode; // @[LazyModule.scala 311:12]
  assign auto_out_c_bits_param = auto_in_0_c_bits_param; // @[LazyModule.scala 311:12]
  assign auto_out_c_bits_size = auto_in_0_c_bits_size; // @[LazyModule.scala 311:12]
  assign auto_out_c_bits_source = {{1'd0}, auto_in_0_c_bits_source}; // @[LazyModule.scala 311:12]
  assign auto_out_c_bits_address = auto_in_0_c_bits_address; // @[LazyModule.scala 311:12]
  assign auto_out_c_bits_data = auto_in_0_c_bits_data; // @[LazyModule.scala 311:12]
  assign auto_out_d_ready = _portsDIO_out_0_d_ready_T | requestDOI_0_1; // @[LazyModule.scala 311:12]
  assign auto_out_e_valid = auto_in_0_e_valid; // @[LazyModule.scala 311:12]
  assign auto_out_e_bits_sink = auto_in_0_e_bits_sink; // @[LazyModule.scala 311:12]
  assign monitor_clock = clock;
  assign monitor_reset = reset;
  assign monitor_io_in_a_ready = auto_out_a_ready & allowed_0; // @[Nodes.scala 25:19]
  assign monitor_io_in_a_valid = auto_in_0_a_valid; // @[Nodes.scala 25:19]
  assign monitor_io_in_a_bits_opcode = auto_in_0_a_bits_opcode; // @[Nodes.scala 25:19]
  assign monitor_io_in_a_bits_param = auto_in_0_a_bits_param; // @[Nodes.scala 25:19]
  assign monitor_io_in_a_bits_size = auto_in_0_a_bits_size; // @[Nodes.scala 25:19]
  assign monitor_io_in_a_bits_source = auto_in_0_a_bits_source; // @[Nodes.scala 25:19]
  assign monitor_io_in_a_bits_address = auto_in_0_a_bits_address; // @[Nodes.scala 25:19]
  assign monitor_io_in_a_bits_mask = auto_in_0_a_bits_mask; // @[Nodes.scala 25:19]
  assign monitor_io_in_b_ready = auto_in_0_b_ready; // @[Nodes.scala 25:19]
  assign monitor_io_in_b_valid = auto_out_b_valid & requestBOI_0_0; // @[Nodes.scala 25:19]
  assign monitor_io_in_b_bits_opcode = auto_out_b_bits_opcode; // @[Nodes.scala 25:19]
  assign monitor_io_in_b_bits_param = auto_out_b_bits_param; // @[Nodes.scala 25:19]
  assign monitor_io_in_b_bits_size = auto_out_b_bits_size; // @[Nodes.scala 25:19]
  assign monitor_io_in_b_bits_source = auto_out_b_bits_source[0]; // @[Nodes.scala 25:19]
  assign monitor_io_in_b_bits_address = auto_out_b_bits_address; // @[Nodes.scala 25:19]
  assign monitor_io_in_b_bits_mask = auto_out_b_bits_mask; // @[Nodes.scala 25:19]
  assign monitor_io_in_b_bits_corrupt = auto_out_b_bits_corrupt; // @[Nodes.scala 25:19]
  assign monitor_io_in_c_ready = auto_out_c_ready; // @[Nodes.scala 25:19]
  assign monitor_io_in_c_valid = auto_in_0_c_valid; // @[Nodes.scala 25:19]
  assign monitor_io_in_c_bits_opcode = auto_in_0_c_bits_opcode; // @[Nodes.scala 25:19]
  assign monitor_io_in_c_bits_param = auto_in_0_c_bits_param; // @[Nodes.scala 25:19]
  assign monitor_io_in_c_bits_size = auto_in_0_c_bits_size; // @[Nodes.scala 25:19]
  assign monitor_io_in_c_bits_source = auto_in_0_c_bits_source; // @[Nodes.scala 25:19]
  assign monitor_io_in_c_bits_address = auto_in_0_c_bits_address; // @[Nodes.scala 25:19]
  assign monitor_io_in_d_ready = auto_in_0_d_ready; // @[Nodes.scala 25:19]
  assign monitor_io_in_d_valid = auto_out_d_valid & requestDOI_0_0; // @[Nodes.scala 25:19]
  assign monitor_io_in_d_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 25:19]
  assign monitor_io_in_d_bits_param = auto_out_d_bits_param; // @[Nodes.scala 25:19]
  assign monitor_io_in_d_bits_size = auto_out_d_bits_size; // @[Nodes.scala 25:19]
  assign monitor_io_in_d_bits_source = auto_out_d_bits_source[0]; // @[Nodes.scala 25:19]
  assign monitor_io_in_d_bits_sink = auto_out_d_bits_sink; // @[Nodes.scala 25:19]
  assign monitor_io_in_d_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 25:19]
  assign monitor_io_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[Nodes.scala 25:19]
  assign monitor_io_in_e_ready = auto_out_e_ready; // @[Nodes.scala 25:19]
  assign monitor_io_in_e_valid = auto_in_0_e_valid; // @[Nodes.scala 25:19]
  assign monitor_io_in_e_bits_sink = auto_in_0_e_bits_sink; // @[Nodes.scala 25:19]
  assign monitor_1_clock = clock;
  assign monitor_1_reset = reset;
  assign monitor_1_io_in_a_ready = auto_out_a_ready & allowed_1; // @[Nodes.scala 25:19]
  assign monitor_1_io_in_a_valid = auto_in_1_a_valid; // @[Nodes.scala 25:19]
  assign monitor_1_io_in_a_bits_address = auto_in_1_a_bits_address; // @[Nodes.scala 25:19]
  assign monitor_1_io_in_d_valid = auto_out_d_valid & requestDOI_0_1; // @[Nodes.scala 25:19]
  assign monitor_1_io_in_d_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 25:19]
  assign monitor_1_io_in_d_bits_param = auto_out_d_bits_param; // @[Nodes.scala 25:19]
  assign monitor_1_io_in_d_bits_size = auto_out_d_bits_size; // @[Nodes.scala 25:19]
  assign monitor_1_io_in_d_bits_sink = auto_out_d_bits_sink; // @[Nodes.scala 25:19]
  assign monitor_1_io_in_d_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 25:19]
  assign monitor_1_io_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[Nodes.scala 25:19]
  assign TLXbar_7_cov_read_addr = TLXbar_7_state;
  assign TLXbar_7_cov_read_data = TLXbar_7_cov[TLXbar_7_cov_read_addr]; // @[Coverage map for TLXbar_7]
  assign TLXbar_7_cov_write_data = 1'h1;
  assign TLXbar_7_cov_write_addr = TLXbar_7_state;
  assign TLXbar_7_cov_write_mask = 1'h1;
  assign TLXbar_7_cov_write_en = 1'h1;
  assign readys_mask_shl = readys_mask;
  assign readys_mask_pad = {1'h0,readys_mask_shl};
  assign state_0_shl = {state_0, 2'h0};
  assign state_0_pad = state_0_shl;
  assign state_1_shl = {state_1, 2'h0};
  assign state_1_pad = state_1_shl;
  assign TLXbar_7_xor2 = state_0_pad ^ state_1_pad;
  assign TLXbar_7_xor0 = readys_mask_pad ^ TLXbar_7_xor2;
  assign monitor_sum = TLXbar_7_covSum + monitor_io_covSum;
  assign monitor_1_sum = monitor_sum + monitor_1_io_covSum;
  assign io_covSum = monitor_1_sum;
  assign stopEn0 = ~_readys_T_3;
  assign stopEn1 = ~_T_9;
  assign stopEn2 = ~_T_16;
  assign stopEn3 = ~_T_23;
  assign monitor_metaAssert_wire = monitor_metaAssert;
  assign monitor_1_metaAssert_wire = monitor_1_metaAssert;
  assign TLXbar_7_or4 = stopEn1 | stopEn2;
  assign TLXbar_7_or1 = stopEn0 | TLXbar_7_or4;
  assign TLXbar_7_or6 = monitor_metaAssert_wire | monitor_1_metaAssert_wire;
  assign TLXbar_7_or2 = stopEn3 | TLXbar_7_or6;
  assign TLXbar_7_or0 = TLXbar_7_or1 | TLXbar_7_or2;
  assign metaAssert = TLXbar_7_metaAssert;
  assign monitor_metaReset = metaReset | monitor_halt;
  assign monitor_1_metaReset = metaReset | monitor_1_halt;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  beatsLeft = _RAND_0[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  readys_mask = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  state_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  state_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  TLXbar_7_state = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    TLXbar_7_cov[initvar] = _RAND_5[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  TLXbar_7_covSum = _RAND_6[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  TLXbar_7_metaAssert = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      beatsLeft <= 9'h0;
    end else if (reset) begin
      beatsLeft <= 9'h0;
    end else if (latch) begin
      if (earlyWinner_0) begin
        if (beatsAI_opdata) begin
          beatsLeft <= beatsAI_decode;
        end else begin
          beatsLeft <= 9'h0;
        end
      end else begin
        beatsLeft <= 9'h0;
      end
    end else begin
      beatsLeft <= _beatsLeft_T_4;
    end
    if (metaReset) begin
      readys_mask <= 2'h0;
    end else if (reset) begin
      readys_mask <= 2'h3;
    end else if (_readys_T_6) begin
      readys_mask <= _readys_mask_T_3;
    end
    if (metaReset) begin
      state_0 <= 1'h0;
    end else if (reset) begin
      state_0 <= 1'h0;
    end else if (idle) begin
      state_0 <= earlyWinner_0;
    end
    if (metaReset) begin
      state_1 <= 1'h0;
    end else if (reset) begin
      state_1 <= 1'h0;
    end else if (idle) begin
      state_1 <= earlyWinner_1;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_readys_T_3) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:22 assert (valid === valids)\n"); // @[Arbiter.scala 22:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_readys_T_3) begin
          $fatal; // @[Arbiter.scala 22:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_9) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:105 assert((prefixOR zip earlyWinner) map { case (p,w) => !p || !w } reduce {_ && _})\n"); // @[Arbiter.scala 105:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_9) begin
          $fatal; // @[Arbiter.scala 105:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_16) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:107 assert (!earlyValids.reduce(_||_) || earlyWinner.reduce(_||_))\n"); // @[Arbiter.scala 107:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_16) begin
          $fatal; // @[Arbiter.scala 107:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_23) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:108 assert (!validQuals .reduce(_||_) || validQuals .reduce(_||_))\n"); // @[Arbiter.scala 108:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_23) begin
          $fatal; // @[Arbiter.scala 108:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    TLXbar_7_state <= TLXbar_7_xor0;
    if (!(TLXbar_7_cov_read_data)) begin
      TLXbar_7_covSum <= TLXbar_7_covSum + 1'h1;
    end
    if (metaReset) begin
      TLXbar_7_metaAssert <= 1'h0;
    end else begin
      TLXbar_7_metaAssert <= TLXbar_7_metaAssert | TLXbar_7_or0;
    end
  end
  always @(posedge clock) begin
    if(TLXbar_7_cov_write_en & TLXbar_7_cov_write_mask) begin
      TLXbar_7_cov[TLXbar_7_cov_write_addr] <= TLXbar_7_cov_write_data; // @[Coverage map for TLXbar_7]
    end
  end
endmodule
module IntXbar_1(
  input         auto_int_in_3_0,
  input         auto_int_in_2_0,
  input         auto_int_in_1_0,
  input         auto_int_in_1_1,
  input         auto_int_in_0_0,
  output        auto_int_out_0,
  output        auto_int_out_1,
  output        auto_int_out_2,
  output        auto_int_out_3,
  output        auto_int_out_4,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire [29:0] IntXbar_1_covSum;
  assign auto_int_out_0 = auto_int_in_0_0; // @[LazyModule.scala 311:12]
  assign auto_int_out_1 = auto_int_in_1_0; // @[LazyModule.scala 311:12]
  assign auto_int_out_2 = auto_int_in_1_1; // @[LazyModule.scala 311:12]
  assign auto_int_out_3 = auto_int_in_2_0; // @[LazyModule.scala 311:12]
  assign auto_int_out_4 = auto_int_in_3_0; // @[LazyModule.scala 311:12]
  assign IntXbar_1_covSum = 30'h0;
  assign io_covSum = IntXbar_1_covSum;
  assign metaAssert = 1'h0;
endmodule
module BundleBridgeNexus_6(
  input         auto_in,
  output        auto_out,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire [29:0] BundleBridgeNexus_6_covSum;
  assign auto_out = auto_in; // @[LazyModule.scala 311:12]
  assign BundleBridgeNexus_6_covSum = 30'h0;
  assign io_covSum = BundleBridgeNexus_6_covSum;
  assign metaAssert = 1'h0;
endmodule
module BundleBridgeNexus_7(
  input  [31:0] auto_in,
  output [31:0] auto_out_1,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire [29:0] BundleBridgeNexus_7_covSum;
  assign auto_out_1 = auto_in; // @[LazyModule.scala 311:12]
  assign BundleBridgeNexus_7_covSum = 30'h0;
  assign io_covSum = BundleBridgeNexus_7_covSum;
  assign metaAssert = 1'h0;
endmodule
module BundleBridgeNexus_10(
  input         auto_in_0_valid,
  input  [39:0] auto_in_0_iaddr,
  input  [31:0] auto_in_0_insn,
  input  [2:0]  auto_in_0_priv,
  input         auto_in_0_exception,
  input         auto_in_0_interrupt,
  input  [63:0] auto_in_0_cause,
  input  [39:0] auto_in_0_tval,
  output        auto_out_0_valid,
  output [39:0] auto_out_0_iaddr,
  output [31:0] auto_out_0_insn,
  output [2:0]  auto_out_0_priv,
  output        auto_out_0_exception,
  output        auto_out_0_interrupt,
  output [63:0] auto_out_0_cause,
  output [39:0] auto_out_0_tval,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire [29:0] BundleBridgeNexus_10_covSum;
  assign auto_out_0_valid = auto_in_0_valid; // @[LazyModule.scala 311:12]
  assign auto_out_0_iaddr = auto_in_0_iaddr; // @[LazyModule.scala 311:12]
  assign auto_out_0_insn = auto_in_0_insn; // @[LazyModule.scala 311:12]
  assign auto_out_0_priv = auto_in_0_priv; // @[LazyModule.scala 311:12]
  assign auto_out_0_exception = auto_in_0_exception; // @[LazyModule.scala 311:12]
  assign auto_out_0_interrupt = auto_in_0_interrupt; // @[LazyModule.scala 311:12]
  assign auto_out_0_cause = auto_in_0_cause; // @[LazyModule.scala 311:12]
  assign auto_out_0_tval = auto_in_0_tval; // @[LazyModule.scala 311:12]
  assign BundleBridgeNexus_10_covSum = 30'h0;
  assign io_covSum = BundleBridgeNexus_10_covSum;
  assign metaAssert = 1'h0;
endmodule
module DCache(
  input         gated_clock,
  input         reset,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_opcode,
  output [2:0]  auto_out_a_bits_param,
  output [3:0]  auto_out_a_bits_size,
  output        auto_out_a_bits_source,
  output [31:0] auto_out_a_bits_address,
  output [7:0]  auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input  [1:0]  auto_out_b_bits_param,
  input  [3:0]  auto_out_b_bits_size,
  input         auto_out_b_bits_source,
  input  [31:0] auto_out_b_bits_address,
  input         auto_out_c_ready,
  output        auto_out_c_valid,
  output [2:0]  auto_out_c_bits_opcode,
  output [2:0]  auto_out_c_bits_param,
  output [3:0]  auto_out_c_bits_size,
  output        auto_out_c_bits_source,
  output [31:0] auto_out_c_bits_address,
  output [63:0] auto_out_c_bits_data,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [2:0]  auto_out_d_bits_opcode,
  input  [1:0]  auto_out_d_bits_param,
  input  [3:0]  auto_out_d_bits_size,
  input         auto_out_d_bits_source,
  input  [1:0]  auto_out_d_bits_sink,
  input         auto_out_d_bits_denied,
  input  [63:0] auto_out_d_bits_data,
  input         auto_out_e_ready,
  output        auto_out_e_valid,
  output [1:0]  auto_out_e_bits_sink,
  output        io_cpu_req_ready,
  input         io_cpu_req_valid,
  input  [39:0] io_cpu_req_bits_addr,
  input  [6:0]  io_cpu_req_bits_tag,
  input  [4:0]  io_cpu_req_bits_cmd,
  input  [1:0]  io_cpu_req_bits_size,
  input         io_cpu_req_bits_signed,
  input         io_cpu_req_bits_phys,
  input         io_cpu_s1_kill,
  input  [63:0] io_cpu_s1_data_data,
  output        io_cpu_s2_nack,
  output        io_cpu_resp_valid,
  output [6:0]  io_cpu_resp_bits_tag,
  output [1:0]  io_cpu_resp_bits_size,
  output [63:0] io_cpu_resp_bits_data,
  output        io_cpu_resp_bits_replay,
  output        io_cpu_resp_bits_has_data,
  output [63:0] io_cpu_resp_bits_data_word_bypass,
  output        io_cpu_replay_next,
  output        io_cpu_s2_xcpt_ma_ld,
  output        io_cpu_s2_xcpt_ma_st,
  output        io_cpu_s2_xcpt_pf_ld,
  output        io_cpu_s2_xcpt_pf_st,
  output        io_cpu_s2_xcpt_ae_ld,
  output        io_cpu_s2_xcpt_ae_st,
  output        io_cpu_ordered,
  output        io_cpu_perf_release,
  output        io_cpu_perf_grant,
  input         io_ptw_req_ready,
  output        io_ptw_req_valid,
  output [26:0] io_ptw_req_bits_bits_addr,
  input         io_ptw_resp_valid,
  input         io_ptw_resp_bits_ae,
  input  [53:0] io_ptw_resp_bits_pte_ppn,
  input         io_ptw_resp_bits_pte_d,
  input         io_ptw_resp_bits_pte_a,
  input         io_ptw_resp_bits_pte_g,
  input         io_ptw_resp_bits_pte_u,
  input         io_ptw_resp_bits_pte_x,
  input         io_ptw_resp_bits_pte_w,
  input         io_ptw_resp_bits_pte_r,
  input         io_ptw_resp_bits_pte_v,
  input  [1:0]  io_ptw_resp_bits_level,
  input         io_ptw_resp_bits_homogeneous,
  input  [3:0]  io_ptw_ptbr_mode,
  input         io_ptw_status_debug,
  input  [1:0]  io_ptw_status_dprv,
  input         io_ptw_status_mxr,
  input         io_ptw_status_sum,
  input         io_ptw_pmp_0_cfg_l,
  input  [1:0]  io_ptw_pmp_0_cfg_a,
  input         io_ptw_pmp_0_cfg_x,
  input         io_ptw_pmp_0_cfg_w,
  input         io_ptw_pmp_0_cfg_r,
  input  [29:0] io_ptw_pmp_0_addr,
  input  [31:0] io_ptw_pmp_0_mask,
  input         io_ptw_pmp_1_cfg_l,
  input  [1:0]  io_ptw_pmp_1_cfg_a,
  input         io_ptw_pmp_1_cfg_x,
  input         io_ptw_pmp_1_cfg_w,
  input         io_ptw_pmp_1_cfg_r,
  input  [29:0] io_ptw_pmp_1_addr,
  input  [31:0] io_ptw_pmp_1_mask,
  input         io_ptw_pmp_2_cfg_l,
  input  [1:0]  io_ptw_pmp_2_cfg_a,
  input         io_ptw_pmp_2_cfg_x,
  input         io_ptw_pmp_2_cfg_w,
  input         io_ptw_pmp_2_cfg_r,
  input  [29:0] io_ptw_pmp_2_addr,
  input  [31:0] io_ptw_pmp_2_mask,
  input         io_ptw_pmp_3_cfg_l,
  input  [1:0]  io_ptw_pmp_3_cfg_a,
  input         io_ptw_pmp_3_cfg_x,
  input         io_ptw_pmp_3_cfg_w,
  input         io_ptw_pmp_3_cfg_r,
  input  [29:0] io_ptw_pmp_3_addr,
  input  [31:0] io_ptw_pmp_3_mask,
  input         io_ptw_pmp_4_cfg_l,
  input  [1:0]  io_ptw_pmp_4_cfg_a,
  input         io_ptw_pmp_4_cfg_x,
  input         io_ptw_pmp_4_cfg_w,
  input         io_ptw_pmp_4_cfg_r,
  input  [29:0] io_ptw_pmp_4_addr,
  input  [31:0] io_ptw_pmp_4_mask,
  input         io_ptw_pmp_5_cfg_l,
  input  [1:0]  io_ptw_pmp_5_cfg_a,
  input         io_ptw_pmp_5_cfg_x,
  input         io_ptw_pmp_5_cfg_w,
  input         io_ptw_pmp_5_cfg_r,
  input  [29:0] io_ptw_pmp_5_addr,
  input  [31:0] io_ptw_pmp_5_mask,
  input         io_ptw_pmp_6_cfg_l,
  input  [1:0]  io_ptw_pmp_6_cfg_a,
  input         io_ptw_pmp_6_cfg_x,
  input         io_ptw_pmp_6_cfg_w,
  input         io_ptw_pmp_6_cfg_r,
  input  [29:0] io_ptw_pmp_6_addr,
  input  [31:0] io_ptw_pmp_6_mask,
  input         io_ptw_pmp_7_cfg_l,
  input  [1:0]  io_ptw_pmp_7_cfg_a,
  input         io_ptw_pmp_7_cfg_x,
  input         io_ptw_pmp_7_cfg_w,
  input         io_ptw_pmp_7_cfg_r,
  input  [29:0] io_ptw_pmp_7_addr,
  input  [31:0] io_ptw_pmp_7_mask,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset,
  input         data_halt,
  input         tlb_halt,
  input         pma_checker_halt,
  input         lfsr_prng_halt
);
  wire  tlb_clock; // @[DCache.scala 117:19]
  wire  tlb_reset; // @[DCache.scala 117:19]
  wire  tlb_io_req_ready; // @[DCache.scala 117:19]
  wire  tlb_io_req_valid; // @[DCache.scala 117:19]
  wire [39:0] tlb_io_req_bits_vaddr; // @[DCache.scala 117:19]
  wire  tlb_io_req_bits_passthrough; // @[DCache.scala 117:19]
  wire [1:0] tlb_io_req_bits_size; // @[DCache.scala 117:19]
  wire [4:0] tlb_io_req_bits_cmd; // @[DCache.scala 117:19]
  wire  tlb_io_resp_miss; // @[DCache.scala 117:19]
  wire [31:0] tlb_io_resp_paddr; // @[DCache.scala 117:19]
  wire  tlb_io_resp_pf_ld; // @[DCache.scala 117:19]
  wire  tlb_io_resp_pf_st; // @[DCache.scala 117:19]
  wire  tlb_io_resp_ae_ld; // @[DCache.scala 117:19]
  wire  tlb_io_resp_ae_st; // @[DCache.scala 117:19]
  wire  tlb_io_resp_ma_ld; // @[DCache.scala 117:19]
  wire  tlb_io_resp_ma_st; // @[DCache.scala 117:19]
  wire  tlb_io_resp_cacheable; // @[DCache.scala 117:19]
  wire  tlb_io_sfence_valid; // @[DCache.scala 117:19]
  wire  tlb_io_sfence_bits_rs1; // @[DCache.scala 117:19]
  wire  tlb_io_sfence_bits_rs2; // @[DCache.scala 117:19]
  wire [38:0] tlb_io_sfence_bits_addr; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_req_ready; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_req_valid; // @[DCache.scala 117:19]
  wire [26:0] tlb_io_ptw_req_bits_bits_addr; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_resp_valid; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_resp_bits_ae; // @[DCache.scala 117:19]
  wire [53:0] tlb_io_ptw_resp_bits_pte_ppn; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_resp_bits_pte_d; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_resp_bits_pte_a; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_resp_bits_pte_g; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_resp_bits_pte_u; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_resp_bits_pte_x; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_resp_bits_pte_w; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_resp_bits_pte_r; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_resp_bits_pte_v; // @[DCache.scala 117:19]
  wire [1:0] tlb_io_ptw_resp_bits_level; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_resp_bits_homogeneous; // @[DCache.scala 117:19]
  wire [3:0] tlb_io_ptw_ptbr_mode; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_status_debug; // @[DCache.scala 117:19]
  wire [1:0] tlb_io_ptw_status_dprv; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_status_mxr; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_status_sum; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_pmp_0_cfg_l; // @[DCache.scala 117:19]
  wire [1:0] tlb_io_ptw_pmp_0_cfg_a; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_pmp_0_cfg_x; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_pmp_0_cfg_w; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_pmp_0_cfg_r; // @[DCache.scala 117:19]
  wire [29:0] tlb_io_ptw_pmp_0_addr; // @[DCache.scala 117:19]
  wire [31:0] tlb_io_ptw_pmp_0_mask; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_pmp_1_cfg_l; // @[DCache.scala 117:19]
  wire [1:0] tlb_io_ptw_pmp_1_cfg_a; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_pmp_1_cfg_x; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_pmp_1_cfg_w; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_pmp_1_cfg_r; // @[DCache.scala 117:19]
  wire [29:0] tlb_io_ptw_pmp_1_addr; // @[DCache.scala 117:19]
  wire [31:0] tlb_io_ptw_pmp_1_mask; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_pmp_2_cfg_l; // @[DCache.scala 117:19]
  wire [1:0] tlb_io_ptw_pmp_2_cfg_a; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_pmp_2_cfg_x; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_pmp_2_cfg_w; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_pmp_2_cfg_r; // @[DCache.scala 117:19]
  wire [29:0] tlb_io_ptw_pmp_2_addr; // @[DCache.scala 117:19]
  wire [31:0] tlb_io_ptw_pmp_2_mask; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_pmp_3_cfg_l; // @[DCache.scala 117:19]
  wire [1:0] tlb_io_ptw_pmp_3_cfg_a; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_pmp_3_cfg_x; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_pmp_3_cfg_w; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_pmp_3_cfg_r; // @[DCache.scala 117:19]
  wire [29:0] tlb_io_ptw_pmp_3_addr; // @[DCache.scala 117:19]
  wire [31:0] tlb_io_ptw_pmp_3_mask; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_pmp_4_cfg_l; // @[DCache.scala 117:19]
  wire [1:0] tlb_io_ptw_pmp_4_cfg_a; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_pmp_4_cfg_x; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_pmp_4_cfg_w; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_pmp_4_cfg_r; // @[DCache.scala 117:19]
  wire [29:0] tlb_io_ptw_pmp_4_addr; // @[DCache.scala 117:19]
  wire [31:0] tlb_io_ptw_pmp_4_mask; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_pmp_5_cfg_l; // @[DCache.scala 117:19]
  wire [1:0] tlb_io_ptw_pmp_5_cfg_a; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_pmp_5_cfg_x; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_pmp_5_cfg_w; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_pmp_5_cfg_r; // @[DCache.scala 117:19]
  wire [29:0] tlb_io_ptw_pmp_5_addr; // @[DCache.scala 117:19]
  wire [31:0] tlb_io_ptw_pmp_5_mask; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_pmp_6_cfg_l; // @[DCache.scala 117:19]
  wire [1:0] tlb_io_ptw_pmp_6_cfg_a; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_pmp_6_cfg_x; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_pmp_6_cfg_w; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_pmp_6_cfg_r; // @[DCache.scala 117:19]
  wire [29:0] tlb_io_ptw_pmp_6_addr; // @[DCache.scala 117:19]
  wire [31:0] tlb_io_ptw_pmp_6_mask; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_pmp_7_cfg_l; // @[DCache.scala 117:19]
  wire [1:0] tlb_io_ptw_pmp_7_cfg_a; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_pmp_7_cfg_x; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_pmp_7_cfg_w; // @[DCache.scala 117:19]
  wire  tlb_io_ptw_pmp_7_cfg_r; // @[DCache.scala 117:19]
  wire [29:0] tlb_io_ptw_pmp_7_addr; // @[DCache.scala 117:19]
  wire [31:0] tlb_io_ptw_pmp_7_mask; // @[DCache.scala 117:19]
  wire [29:0] tlb_io_covSum; // @[DCache.scala 117:19]
  wire  tlb_metaAssert; // @[DCache.scala 117:19]
  wire  tlb_metaReset; // @[DCache.scala 117:19]
  wire  pma_checker_clock; // @[DCache.scala 118:27]
  wire  pma_checker_reset; // @[DCache.scala 118:27]
  wire  pma_checker_io_req_ready; // @[DCache.scala 118:27]
  wire  pma_checker_io_req_valid; // @[DCache.scala 118:27]
  wire [39:0] pma_checker_io_req_bits_vaddr; // @[DCache.scala 118:27]
  wire  pma_checker_io_req_bits_passthrough; // @[DCache.scala 118:27]
  wire [1:0] pma_checker_io_req_bits_size; // @[DCache.scala 118:27]
  wire [4:0] pma_checker_io_req_bits_cmd; // @[DCache.scala 118:27]
  wire  pma_checker_io_resp_miss; // @[DCache.scala 118:27]
  wire [31:0] pma_checker_io_resp_paddr; // @[DCache.scala 118:27]
  wire  pma_checker_io_resp_pf_ld; // @[DCache.scala 118:27]
  wire  pma_checker_io_resp_pf_st; // @[DCache.scala 118:27]
  wire  pma_checker_io_resp_ae_ld; // @[DCache.scala 118:27]
  wire  pma_checker_io_resp_ae_st; // @[DCache.scala 118:27]
  wire  pma_checker_io_resp_ma_ld; // @[DCache.scala 118:27]
  wire  pma_checker_io_resp_ma_st; // @[DCache.scala 118:27]
  wire  pma_checker_io_resp_cacheable; // @[DCache.scala 118:27]
  wire  pma_checker_io_sfence_valid; // @[DCache.scala 118:27]
  wire  pma_checker_io_sfence_bits_rs1; // @[DCache.scala 118:27]
  wire  pma_checker_io_sfence_bits_rs2; // @[DCache.scala 118:27]
  wire [38:0] pma_checker_io_sfence_bits_addr; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_req_ready; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_req_valid; // @[DCache.scala 118:27]
  wire [26:0] pma_checker_io_ptw_req_bits_bits_addr; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_resp_valid; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_resp_bits_ae; // @[DCache.scala 118:27]
  wire [53:0] pma_checker_io_ptw_resp_bits_pte_ppn; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_resp_bits_pte_d; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_resp_bits_pte_a; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_resp_bits_pte_g; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_resp_bits_pte_u; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_resp_bits_pte_x; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_resp_bits_pte_w; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_resp_bits_pte_r; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_resp_bits_pte_v; // @[DCache.scala 118:27]
  wire [1:0] pma_checker_io_ptw_resp_bits_level; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_resp_bits_homogeneous; // @[DCache.scala 118:27]
  wire [3:0] pma_checker_io_ptw_ptbr_mode; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_status_debug; // @[DCache.scala 118:27]
  wire [1:0] pma_checker_io_ptw_status_dprv; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_status_mxr; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_status_sum; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_pmp_0_cfg_l; // @[DCache.scala 118:27]
  wire [1:0] pma_checker_io_ptw_pmp_0_cfg_a; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_pmp_0_cfg_x; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_pmp_0_cfg_w; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_pmp_0_cfg_r; // @[DCache.scala 118:27]
  wire [29:0] pma_checker_io_ptw_pmp_0_addr; // @[DCache.scala 118:27]
  wire [31:0] pma_checker_io_ptw_pmp_0_mask; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_pmp_1_cfg_l; // @[DCache.scala 118:27]
  wire [1:0] pma_checker_io_ptw_pmp_1_cfg_a; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_pmp_1_cfg_x; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_pmp_1_cfg_w; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_pmp_1_cfg_r; // @[DCache.scala 118:27]
  wire [29:0] pma_checker_io_ptw_pmp_1_addr; // @[DCache.scala 118:27]
  wire [31:0] pma_checker_io_ptw_pmp_1_mask; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_pmp_2_cfg_l; // @[DCache.scala 118:27]
  wire [1:0] pma_checker_io_ptw_pmp_2_cfg_a; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_pmp_2_cfg_x; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_pmp_2_cfg_w; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_pmp_2_cfg_r; // @[DCache.scala 118:27]
  wire [29:0] pma_checker_io_ptw_pmp_2_addr; // @[DCache.scala 118:27]
  wire [31:0] pma_checker_io_ptw_pmp_2_mask; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_pmp_3_cfg_l; // @[DCache.scala 118:27]
  wire [1:0] pma_checker_io_ptw_pmp_3_cfg_a; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_pmp_3_cfg_x; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_pmp_3_cfg_w; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_pmp_3_cfg_r; // @[DCache.scala 118:27]
  wire [29:0] pma_checker_io_ptw_pmp_3_addr; // @[DCache.scala 118:27]
  wire [31:0] pma_checker_io_ptw_pmp_3_mask; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_pmp_4_cfg_l; // @[DCache.scala 118:27]
  wire [1:0] pma_checker_io_ptw_pmp_4_cfg_a; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_pmp_4_cfg_x; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_pmp_4_cfg_w; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_pmp_4_cfg_r; // @[DCache.scala 118:27]
  wire [29:0] pma_checker_io_ptw_pmp_4_addr; // @[DCache.scala 118:27]
  wire [31:0] pma_checker_io_ptw_pmp_4_mask; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_pmp_5_cfg_l; // @[DCache.scala 118:27]
  wire [1:0] pma_checker_io_ptw_pmp_5_cfg_a; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_pmp_5_cfg_x; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_pmp_5_cfg_w; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_pmp_5_cfg_r; // @[DCache.scala 118:27]
  wire [29:0] pma_checker_io_ptw_pmp_5_addr; // @[DCache.scala 118:27]
  wire [31:0] pma_checker_io_ptw_pmp_5_mask; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_pmp_6_cfg_l; // @[DCache.scala 118:27]
  wire [1:0] pma_checker_io_ptw_pmp_6_cfg_a; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_pmp_6_cfg_x; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_pmp_6_cfg_w; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_pmp_6_cfg_r; // @[DCache.scala 118:27]
  wire [29:0] pma_checker_io_ptw_pmp_6_addr; // @[DCache.scala 118:27]
  wire [31:0] pma_checker_io_ptw_pmp_6_mask; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_pmp_7_cfg_l; // @[DCache.scala 118:27]
  wire [1:0] pma_checker_io_ptw_pmp_7_cfg_a; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_pmp_7_cfg_x; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_pmp_7_cfg_w; // @[DCache.scala 118:27]
  wire  pma_checker_io_ptw_pmp_7_cfg_r; // @[DCache.scala 118:27]
  wire [29:0] pma_checker_io_ptw_pmp_7_addr; // @[DCache.scala 118:27]
  wire [31:0] pma_checker_io_ptw_pmp_7_mask; // @[DCache.scala 118:27]
  wire [29:0] pma_checker_io_covSum; // @[DCache.scala 118:27]
  wire  pma_checker_metaAssert; // @[DCache.scala 118:27]
  wire  pma_checker_metaReset; // @[DCache.scala 118:27]
  wire  lfsr_prng_clock; // @[PRNG.scala 82:22]
  wire  lfsr_prng_reset; // @[PRNG.scala 82:22]
  wire  lfsr_prng_io_increment; // @[PRNG.scala 82:22]
  wire  lfsr_prng_io_out_0; // @[PRNG.scala 82:22]
  wire  lfsr_prng_io_out_1; // @[PRNG.scala 82:22]
  wire  lfsr_prng_io_out_2; // @[PRNG.scala 82:22]
  wire  lfsr_prng_io_out_3; // @[PRNG.scala 82:22]
  wire  lfsr_prng_io_out_4; // @[PRNG.scala 82:22]
  wire  lfsr_prng_io_out_5; // @[PRNG.scala 82:22]
  wire  lfsr_prng_io_out_6; // @[PRNG.scala 82:22]
  wire  lfsr_prng_io_out_7; // @[PRNG.scala 82:22]
  wire  lfsr_prng_io_out_8; // @[PRNG.scala 82:22]
  wire  lfsr_prng_io_out_9; // @[PRNG.scala 82:22]
  wire  lfsr_prng_io_out_10; // @[PRNG.scala 82:22]
  wire  lfsr_prng_io_out_11; // @[PRNG.scala 82:22]
  wire  lfsr_prng_io_out_12; // @[PRNG.scala 82:22]
  wire  lfsr_prng_io_out_13; // @[PRNG.scala 82:22]
  wire  lfsr_prng_io_out_14; // @[PRNG.scala 82:22]
  wire  lfsr_prng_io_out_15; // @[PRNG.scala 82:22]
  wire [29:0] lfsr_prng_io_covSum; // @[PRNG.scala 82:22]
  wire  lfsr_prng_metaAssert; // @[PRNG.scala 82:22]
  wire  lfsr_prng_metaReset; // @[PRNG.scala 82:22]
  wire  metaArb_io_in_0_valid; // @[DCache.scala 122:23]
  wire [39:0] metaArb_io_in_0_bits_addr; // @[DCache.scala 122:23]
  wire [5:0] metaArb_io_in_0_bits_idx; // @[DCache.scala 122:23]
  wire  metaArb_io_in_1_valid; // @[DCache.scala 122:23]
  wire [39:0] metaArb_io_in_1_bits_addr; // @[DCache.scala 122:23]
  wire [5:0] metaArb_io_in_1_bits_idx; // @[DCache.scala 122:23]
  wire [21:0] metaArb_io_in_1_bits_data; // @[DCache.scala 122:23]
  wire  metaArb_io_in_2_valid; // @[DCache.scala 122:23]
  wire [39:0] metaArb_io_in_2_bits_addr; // @[DCache.scala 122:23]
  wire [5:0] metaArb_io_in_2_bits_idx; // @[DCache.scala 122:23]
  wire [3:0] metaArb_io_in_2_bits_way_en; // @[DCache.scala 122:23]
  wire [21:0] metaArb_io_in_2_bits_data; // @[DCache.scala 122:23]
  wire  metaArb_io_in_3_valid; // @[DCache.scala 122:23]
  wire [39:0] metaArb_io_in_3_bits_addr; // @[DCache.scala 122:23]
  wire [5:0] metaArb_io_in_3_bits_idx; // @[DCache.scala 122:23]
  wire [3:0] metaArb_io_in_3_bits_way_en; // @[DCache.scala 122:23]
  wire [21:0] metaArb_io_in_3_bits_data; // @[DCache.scala 122:23]
  wire  metaArb_io_in_4_ready; // @[DCache.scala 122:23]
  wire  metaArb_io_in_4_valid; // @[DCache.scala 122:23]
  wire [39:0] metaArb_io_in_4_bits_addr; // @[DCache.scala 122:23]
  wire [5:0] metaArb_io_in_4_bits_idx; // @[DCache.scala 122:23]
  wire [3:0] metaArb_io_in_4_bits_way_en; // @[DCache.scala 122:23]
  wire [21:0] metaArb_io_in_4_bits_data; // @[DCache.scala 122:23]
  wire  metaArb_io_in_5_ready; // @[DCache.scala 122:23]
  wire  metaArb_io_in_5_valid; // @[DCache.scala 122:23]
  wire [39:0] metaArb_io_in_5_bits_addr; // @[DCache.scala 122:23]
  wire [5:0] metaArb_io_in_5_bits_idx; // @[DCache.scala 122:23]
  wire  metaArb_io_in_6_ready; // @[DCache.scala 122:23]
  wire  metaArb_io_in_6_valid; // @[DCache.scala 122:23]
  wire [39:0] metaArb_io_in_6_bits_addr; // @[DCache.scala 122:23]
  wire [5:0] metaArb_io_in_6_bits_idx; // @[DCache.scala 122:23]
  wire [3:0] metaArb_io_in_6_bits_way_en; // @[DCache.scala 122:23]
  wire [21:0] metaArb_io_in_6_bits_data; // @[DCache.scala 122:23]
  wire  metaArb_io_in_7_ready; // @[DCache.scala 122:23]
  wire  metaArb_io_in_7_valid; // @[DCache.scala 122:23]
  wire [39:0] metaArb_io_in_7_bits_addr; // @[DCache.scala 122:23]
  wire [5:0] metaArb_io_in_7_bits_idx; // @[DCache.scala 122:23]
  wire [3:0] metaArb_io_in_7_bits_way_en; // @[DCache.scala 122:23]
  wire [21:0] metaArb_io_in_7_bits_data; // @[DCache.scala 122:23]
  wire  metaArb_io_out_valid; // @[DCache.scala 122:23]
  wire  metaArb_io_out_bits_write; // @[DCache.scala 122:23]
  wire [39:0] metaArb_io_out_bits_addr; // @[DCache.scala 122:23]
  wire [5:0] metaArb_io_out_bits_idx; // @[DCache.scala 122:23]
  wire [3:0] metaArb_io_out_bits_way_en; // @[DCache.scala 122:23]
  wire [21:0] metaArb_io_out_bits_data; // @[DCache.scala 122:23]
  wire [29:0] metaArb_io_covSum; // @[DCache.scala 122:23]
  wire  metaArb_metaAssert; // @[DCache.scala 122:23]
  reg [21:0] tag_array_0 [0:63]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_0;
  wire [21:0] tag_array_0_s1_meta_data; // @[DescribedSRAM.scala 19:26]
  wire [5:0] tag_array_0_s1_meta_addr; // @[DescribedSRAM.scala 19:26]
  wire [21:0] tag_array_0_MPORT_data; // @[DescribedSRAM.scala 19:26]
  wire [5:0] tag_array_0_MPORT_addr; // @[DescribedSRAM.scala 19:26]
  wire  tag_array_0_MPORT_mask; // @[DescribedSRAM.scala 19:26]
  wire  tag_array_0_MPORT_en; // @[DescribedSRAM.scala 19:26]
  reg  tag_array_0_s1_meta_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [5:0] tag_array_0_s1_meta_addr_pipe_0;
  reg [31:0] _RAND_2;
  reg [21:0] tag_array_1 [0:63]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_3;
  wire [21:0] tag_array_1_s1_meta_data; // @[DescribedSRAM.scala 19:26]
  wire [5:0] tag_array_1_s1_meta_addr; // @[DescribedSRAM.scala 19:26]
  wire [21:0] tag_array_1_MPORT_data; // @[DescribedSRAM.scala 19:26]
  wire [5:0] tag_array_1_MPORT_addr; // @[DescribedSRAM.scala 19:26]
  wire  tag_array_1_MPORT_mask; // @[DescribedSRAM.scala 19:26]
  wire  tag_array_1_MPORT_en; // @[DescribedSRAM.scala 19:26]
  reg  tag_array_1_s1_meta_en_pipe_0;
  reg [31:0] _RAND_4;
  reg [5:0] tag_array_1_s1_meta_addr_pipe_0;
  reg [31:0] _RAND_5;
  reg [21:0] tag_array_2 [0:63]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_6;
  wire [21:0] tag_array_2_s1_meta_data; // @[DescribedSRAM.scala 19:26]
  wire [5:0] tag_array_2_s1_meta_addr; // @[DescribedSRAM.scala 19:26]
  wire [21:0] tag_array_2_MPORT_data; // @[DescribedSRAM.scala 19:26]
  wire [5:0] tag_array_2_MPORT_addr; // @[DescribedSRAM.scala 19:26]
  wire  tag_array_2_MPORT_mask; // @[DescribedSRAM.scala 19:26]
  wire  tag_array_2_MPORT_en; // @[DescribedSRAM.scala 19:26]
  reg  tag_array_2_s1_meta_en_pipe_0;
  reg [31:0] _RAND_7;
  reg [5:0] tag_array_2_s1_meta_addr_pipe_0;
  reg [31:0] _RAND_8;
  reg [21:0] tag_array_3 [0:63]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_9;
  wire [21:0] tag_array_3_s1_meta_data; // @[DescribedSRAM.scala 19:26]
  wire [5:0] tag_array_3_s1_meta_addr; // @[DescribedSRAM.scala 19:26]
  wire [21:0] tag_array_3_MPORT_data; // @[DescribedSRAM.scala 19:26]
  wire [5:0] tag_array_3_MPORT_addr; // @[DescribedSRAM.scala 19:26]
  wire  tag_array_3_MPORT_mask; // @[DescribedSRAM.scala 19:26]
  wire  tag_array_3_MPORT_en; // @[DescribedSRAM.scala 19:26]
  reg  tag_array_3_s1_meta_en_pipe_0;
  reg [31:0] _RAND_10;
  reg [5:0] tag_array_3_s1_meta_addr_pipe_0;
  reg [31:0] _RAND_11;
  wire  data_clock; // @[DCache.scala 132:20]
  wire  data_io_req_valid; // @[DCache.scala 132:20]
  wire [11:0] data_io_req_bits_addr; // @[DCache.scala 132:20]
  wire  data_io_req_bits_write; // @[DCache.scala 132:20]
  wire [63:0] data_io_req_bits_wdata; // @[DCache.scala 132:20]
  wire [7:0] data_io_req_bits_eccMask; // @[DCache.scala 132:20]
  wire [3:0] data_io_req_bits_way_en; // @[DCache.scala 132:20]
  wire [63:0] data_io_resp_0; // @[DCache.scala 132:20]
  wire [63:0] data_io_resp_1; // @[DCache.scala 132:20]
  wire [63:0] data_io_resp_2; // @[DCache.scala 132:20]
  wire [63:0] data_io_resp_3; // @[DCache.scala 132:20]
  wire [29:0] data_io_covSum; // @[DCache.scala 132:20]
  wire  data_metaAssert; // @[DCache.scala 132:20]
  wire  data_metaReset; // @[DCache.scala 132:20]
  wire  dataArb_io_in_0_valid; // @[DCache.scala 133:23]
  wire [11:0] dataArb_io_in_0_bits_addr; // @[DCache.scala 133:23]
  wire  dataArb_io_in_0_bits_write; // @[DCache.scala 133:23]
  wire [63:0] dataArb_io_in_0_bits_wdata; // @[DCache.scala 133:23]
  wire [7:0] dataArb_io_in_0_bits_eccMask; // @[DCache.scala 133:23]
  wire [3:0] dataArb_io_in_0_bits_way_en; // @[DCache.scala 133:23]
  wire  dataArb_io_in_1_ready; // @[DCache.scala 133:23]
  wire  dataArb_io_in_1_valid; // @[DCache.scala 133:23]
  wire [11:0] dataArb_io_in_1_bits_addr; // @[DCache.scala 133:23]
  wire  dataArb_io_in_1_bits_write; // @[DCache.scala 133:23]
  wire [63:0] dataArb_io_in_1_bits_wdata; // @[DCache.scala 133:23]
  wire [3:0] dataArb_io_in_1_bits_way_en; // @[DCache.scala 133:23]
  wire  dataArb_io_in_2_ready; // @[DCache.scala 133:23]
  wire  dataArb_io_in_2_valid; // @[DCache.scala 133:23]
  wire [11:0] dataArb_io_in_2_bits_addr; // @[DCache.scala 133:23]
  wire [63:0] dataArb_io_in_2_bits_wdata; // @[DCache.scala 133:23]
  wire  dataArb_io_in_3_ready; // @[DCache.scala 133:23]
  wire  dataArb_io_in_3_valid; // @[DCache.scala 133:23]
  wire [11:0] dataArb_io_in_3_bits_addr; // @[DCache.scala 133:23]
  wire [63:0] dataArb_io_in_3_bits_wdata; // @[DCache.scala 133:23]
  wire  dataArb_io_in_3_bits_wordMask; // @[DCache.scala 133:23]
  wire  dataArb_io_out_valid; // @[DCache.scala 133:23]
  wire [11:0] dataArb_io_out_bits_addr; // @[DCache.scala 133:23]
  wire  dataArb_io_out_bits_write; // @[DCache.scala 133:23]
  wire [63:0] dataArb_io_out_bits_wdata; // @[DCache.scala 133:23]
  wire [7:0] dataArb_io_out_bits_eccMask; // @[DCache.scala 133:23]
  wire [3:0] dataArb_io_out_bits_way_en; // @[DCache.scala 133:23]
  wire [29:0] dataArb_io_covSum; // @[DCache.scala 133:23]
  wire  dataArb_metaAssert; // @[DCache.scala 133:23]
  wire [7:0] amoalu_io_mask; // @[DCache.scala 950:26]
  wire [4:0] amoalu_io_cmd; // @[DCache.scala 950:26]
  wire [63:0] amoalu_io_lhs; // @[DCache.scala 950:26]
  wire [63:0] amoalu_io_rhs; // @[DCache.scala 950:26]
  wire [63:0] amoalu_io_out; // @[DCache.scala 950:26]
  wire [29:0] amoalu_io_covSum; // @[DCache.scala 950:26]
  wire  amoalu_metaAssert; // @[DCache.scala 950:26]
  wire [7:0] lfsr_lo; // @[PRNG.scala 86:17]
  wire [15:0] lfsr; // @[PRNG.scala 86:17]
  wire  s1_valid_x9; // @[Decoupled.scala 40:37]
  reg  s1_valid; // @[DCache.scala 162:21]
  reg [31:0] _RAND_12;
  reg [2:0] blockProbeAfterGrantCount; // @[DCache.scala 639:38]
  reg [31:0] _RAND_13;
  wire  _block_probe_for_core_progress_T; // @[DCache.scala 737:65]
  reg [6:0] lrscCount; // @[DCache.scala 443:22]
  reg [31:0] _RAND_14;
  wire  lrscValid; // @[DCache.scala 444:29]
  wire  block_probe_for_core_progress; // @[DCache.scala 737:69]
  reg  s1_probe; // @[DCache.scala 163:21]
  reg [31:0] _RAND_15;
  reg  s2_probe; // @[DCache.scala 304:21]
  reg [31:0] _RAND_16;
  wire  _releaseInFlight_T; // @[DCache.scala 305:34]
  reg [3:0] release_state; // @[DCache.scala 206:26]
  reg [31:0] _RAND_17;
  wire  _releaseInFlight_T_1; // @[DCache.scala 305:63]
  wire  releaseInFlight; // @[DCache.scala 305:46]
  reg  release_ack_wait; // @[DCache.scala 204:29]
  reg [31:0] _RAND_18;
  reg [31:0] release_ack_addr; // @[DCache.scala 205:29]
  reg [31:0] _RAND_19;
  wire [31:0] _block_probe_for_pending_release_ack_T; // @[DCache.scala 738:88]
  wire  _block_probe_for_pending_release_ack_T_2; // @[DCache.scala 738:163]
  wire  block_probe_for_pending_release_ack; // @[DCache.scala 738:62]
  wire  _block_probe_for_ordering_T; // @[DCache.scala 739:50]
  reg  grantInProgress; // @[DCache.scala 638:28]
  reg [31:0] _RAND_20;
  wire  block_probe_for_ordering; // @[DCache.scala 739:89]
  wire  _bundleOut_0_b_ready_T; // @[DCache.scala 741:79]
  wire  _bundleOut_0_b_ready_T_1; // @[DCache.scala 741:107]
  reg  s2_valid; // @[DCache.scala 302:21]
  reg [31:0] _RAND_21;
  wire  _bundleOut_0_b_ready_T_2; // @[DCache.scala 741:119]
  wire  tl_out__b_ready; // @[DCache.scala 741:44]
  wire  s1_probe_x12; // @[Decoupled.scala 40:37]
  reg [1:0] probe_bits_param; // @[Reg.scala 15:16]
  reg [31:0] _RAND_22;
  reg [3:0] probe_bits_size; // @[Reg.scala 15:16]
  reg [31:0] _RAND_23;
  reg  probe_bits_source; // @[Reg.scala 15:16]
  reg [31:0] _RAND_24;
  reg [31:0] probe_bits_address; // @[Reg.scala 15:16]
  reg [31:0] _RAND_25;
  wire  s1_valid_masked; // @[DCache.scala 166:34]
  wire  s2_meta_error; // @[DCache.scala 333:83]
  reg [1:0] s2_probe_state_state; // @[Reg.scala 15:16]
  reg [31:0] _RAND_26;
  wire [3:0] _T_118; // @[Cat.scala 30:58]
  wire  _T_175; // @[Misc.scala 55:20]
  wire  _T_171; // @[Misc.scala 55:20]
  wire  _T_167; // @[Misc.scala 55:20]
  wire  _T_163; // @[Misc.scala 55:20]
  wire  _T_159; // @[Misc.scala 55:20]
  wire  _T_155; // @[Misc.scala 55:20]
  wire  _T_151; // @[Misc.scala 55:20]
  wire  _T_147; // @[Misc.scala 55:20]
  wire  _T_143; // @[Misc.scala 55:20]
  wire  _T_139; // @[Misc.scala 55:20]
  wire  _T_135; // @[Misc.scala 55:20]
  wire  _T_131; // @[Misc.scala 55:20]
  wire  _T_148; // @[Misc.scala 37:9]
  wire  _T_152; // @[Misc.scala 37:9]
  wire  _T_156; // @[Misc.scala 37:9]
  wire  _T_160; // @[Misc.scala 37:9]
  wire  _T_164; // @[Misc.scala 37:9]
  wire  _T_168; // @[Misc.scala 37:9]
  wire  _T_172; // @[Misc.scala 37:9]
  wire  s2_prb_ack_data; // @[Misc.scala 37:9]
  wire  _T_303; // @[Metadata.scala 49:45]
  reg [8:0] counter_1; // @[Edges.scala 228:27]
  reg [31:0] _RAND_27;
  wire  _last_T_2; // @[Edges.scala 231:25]
  wire  _T_308; // @[package.scala 15:47]
  wire  _T_309; // @[package.scala 15:47]
  wire  _T_311; // @[package.scala 72:59]
  wire  _T_310; // @[package.scala 15:47]
  wire  _T_312; // @[package.scala 72:59]
  wire [2:0] _GEN_323; // @[DCache.scala 835:52]
  wire  _T_307; // @[DCache.scala 830:25]
  wire  _T_306; // @[DCache.scala 825:25]
  wire [2:0] _GEN_315; // @[DCache.scala 830:48]
  wire [2:0] tl_out__c_bits_opcode; // @[DCache.scala 834:102]
  wire  beats1_opdata_1; // @[Edges.scala 101:36]
  wire [3:0] tl_out__c_bits_size; // @[DCache.scala 834:102]
  wire [26:0] _beats1_decode_T_5; // @[package.scala 234:77]
  wire [8:0] beats1_decode_1; // @[Edges.scala 219:59]
  wire [8:0] beats1_1; // @[Edges.scala 220:14]
  wire  _last_T_3; // @[Edges.scala 231:47]
  wire  c_last; // @[Edges.scala 231:37]
  wire  _T_305; // @[DCache.scala 821:25]
  reg  s2_release_data_valid; // @[DCache.scala 773:34]
  reg [31:0] _RAND_28;
  wire  c_first; // @[Edges.scala 230:25]
  wire  _bundleOut_0_c_valid_T_3; // @[DCache.scala 781:128]
  wire  _bundleOut_0_c_valid_T_5; // @[DCache.scala 781:115]
  wire  _GEN_264; // @[DCache.scala 799:36]
  wire  _GEN_274; // @[DCache.scala 797:28]
  wire  _GEN_285; // @[DCache.scala 795:21]
  wire  _GEN_302; // @[DCache.scala 821:47]
  wire  tl_out__c_valid; // @[DCache.scala 825:48]
  wire  _T_297; // @[Decoupled.scala 40:37]
  wire  releaseDone; // @[Edges.scala 232:22]
  wire  _GEN_262; // @[DCache.scala 801:45]
  wire  _GEN_272; // @[DCache.scala 799:36]
  wire  probeNack; // @[DCache.scala 797:28]
  reg [4:0] s1_req_cmd; // @[Reg.scala 15:16]
  reg [31:0] _RAND_29;
  wire  _s1_read_T; // @[Consts.scala 81:31]
  wire  _s1_read_T_1; // @[Consts.scala 81:48]
  wire  _s1_read_T_2; // @[Consts.scala 81:41]
  wire  _s1_read_T_3; // @[Consts.scala 81:65]
  wire  _s1_read_T_4; // @[Consts.scala 81:58]
  wire  _s1_read_T_5; // @[package.scala 15:47]
  wire  _s1_read_T_6; // @[package.scala 15:47]
  wire  _s1_read_T_9; // @[package.scala 72:59]
  wire  _s1_read_T_7; // @[package.scala 15:47]
  wire  _s1_read_T_10; // @[package.scala 72:59]
  wire  _s1_read_T_8; // @[package.scala 15:47]
  wire  _s1_read_T_11; // @[package.scala 72:59]
  wire  _s1_read_T_12; // @[package.scala 15:47]
  wire  _s1_read_T_13; // @[package.scala 15:47]
  wire  _s1_read_T_17; // @[package.scala 72:59]
  wire  _s1_read_T_14; // @[package.scala 15:47]
  wire  _s1_read_T_18; // @[package.scala 72:59]
  wire  _s1_read_T_15; // @[package.scala 15:47]
  wire  _s1_read_T_19; // @[package.scala 72:59]
  wire  _s1_read_T_16; // @[package.scala 15:47]
  wire  _s1_read_T_20; // @[package.scala 72:59]
  wire  _s1_read_T_21; // @[Consts.scala 79:44]
  wire  s1_read; // @[Consts.scala 81:75]
  reg [4:0] s2_req_cmd; // @[DCache.scala 310:19]
  reg [31:0] _RAND_30;
  wire  _s2_write_T; // @[Consts.scala 82:32]
  wire  _s2_write_T_1; // @[Consts.scala 82:49]
  wire  _s2_write_T_2; // @[Consts.scala 82:42]
  wire  _s2_write_T_3; // @[Consts.scala 82:66]
  wire  _s2_write_T_4; // @[Consts.scala 82:59]
  wire  _s2_write_T_5; // @[package.scala 15:47]
  wire  _s2_write_T_6; // @[package.scala 15:47]
  wire  _s2_write_T_9; // @[package.scala 72:59]
  wire  _s2_write_T_7; // @[package.scala 15:47]
  wire  _s2_write_T_10; // @[package.scala 72:59]
  wire  _s2_write_T_8; // @[package.scala 15:47]
  wire  _s2_write_T_11; // @[package.scala 72:59]
  wire  _s2_write_T_12; // @[package.scala 15:47]
  wire  _s2_write_T_13; // @[package.scala 15:47]
  wire  _s2_write_T_17; // @[package.scala 72:59]
  wire  _s2_write_T_14; // @[package.scala 15:47]
  wire  _s2_write_T_18; // @[package.scala 72:59]
  wire  _s2_write_T_15; // @[package.scala 15:47]
  wire  _s2_write_T_19; // @[package.scala 72:59]
  wire  _s2_write_T_16; // @[package.scala 15:47]
  wire  _s2_write_T_20; // @[package.scala 72:59]
  wire  _s2_write_T_21; // @[Consts.scala 79:44]
  wire  s2_write; // @[Consts.scala 82:76]
  wire  _pstore1_valid_likely_T; // @[DCache.scala 476:39]
  reg  pstore1_held; // @[DCache.scala 475:29]
  reg [31:0] _RAND_31;
  wire  pstore1_valid_likely; // @[DCache.scala 476:51]
  reg [39:0] pstore1_addr; // @[Reg.scala 15:16]
  reg [63:0] _RAND_32;
  reg [39:0] s1_req_addr; // @[Reg.scala 15:16]
  reg [63:0] _RAND_33;
  wire [27:0] s1_vaddr_hi; // @[DCache.scala 177:56]
  wire [11:0] s1_vaddr_lo; // @[DCache.scala 177:78]
  wire [39:0] s1_vaddr; // @[Cat.scala 30:58]
  wire  _s1_hazard_T_2; // @[DCache.scala 532:31]
  wire  _s1_write_T; // @[Consts.scala 82:32]
  wire  _s1_write_T_1; // @[Consts.scala 82:49]
  wire  _s1_write_T_2; // @[Consts.scala 82:42]
  wire  _s1_write_T_4; // @[Consts.scala 82:59]
  wire  s1_write; // @[Consts.scala 82:76]
  reg [7:0] pstore1_mask; // @[Reg.scala 15:16]
  reg [31:0] _RAND_34;
  wire  s1_hazard_hi_hi_hi; // @[DCache.scala 1149:66]
  wire  s1_hazard_hi_hi_lo; // @[DCache.scala 1149:66]
  wire  s1_hazard_hi_lo_hi; // @[DCache.scala 1149:66]
  wire  s1_hazard_hi_lo_lo; // @[DCache.scala 1149:66]
  wire  s1_hazard_lo_hi_hi; // @[DCache.scala 1149:66]
  wire  s1_hazard_lo_hi_lo; // @[DCache.scala 1149:66]
  wire  s1_hazard_lo_lo_hi; // @[DCache.scala 1149:66]
  wire  s1_hazard_lo_lo_lo; // @[DCache.scala 1149:66]
  wire [7:0] _s1_hazard_T_11; // @[Cat.scala 30:58]
  wire  s1_hazard_hi_hi_hi_1; // @[Bitwise.scala 26:51]
  wire  s1_hazard_hi_hi_lo_1; // @[Bitwise.scala 26:51]
  wire  s1_hazard_hi_lo_hi_1; // @[Bitwise.scala 26:51]
  wire  s1_hazard_hi_lo_lo_1; // @[Bitwise.scala 26:51]
  wire  s1_hazard_lo_hi_hi_1; // @[Bitwise.scala 26:51]
  wire  s1_hazard_lo_hi_lo_1; // @[Bitwise.scala 26:51]
  wire  s1_hazard_lo_lo_hi_1; // @[Bitwise.scala 26:51]
  wire  s1_hazard_lo_lo_lo_1; // @[Bitwise.scala 26:51]
  wire [7:0] _s1_hazard_T_12; // @[Cat.scala 30:58]
  reg [1:0] s1_req_size; // @[Reg.scala 15:16]
  reg [31:0] _RAND_35;
  wire  _s1_mask_xwr_upper_T_2; // @[AMOALU.scala 17:57]
  wire  s1_mask_xwr_hi; // @[AMOALU.scala 17:46]
  wire  s1_mask_xwr_lo; // @[AMOALU.scala 18:22]
  wire [1:0] _s1_mask_xwr_T; // @[Cat.scala 30:58]
  wire [1:0] _s1_mask_xwr_upper_T_5; // @[AMOALU.scala 17:22]
  wire  _s1_mask_xwr_upper_T_6; // @[AMOALU.scala 17:57]
  wire [1:0] _s1_mask_xwr_upper_T_7; // @[AMOALU.scala 17:51]
  wire [1:0] s1_mask_xwr_hi_1; // @[AMOALU.scala 17:46]
  wire [1:0] s1_mask_xwr_lo_1; // @[AMOALU.scala 18:22]
  wire [3:0] _s1_mask_xwr_T_1; // @[Cat.scala 30:58]
  wire [3:0] _s1_mask_xwr_upper_T_9; // @[AMOALU.scala 17:22]
  wire  _s1_mask_xwr_upper_T_10; // @[AMOALU.scala 17:57]
  wire [3:0] _s1_mask_xwr_upper_T_11; // @[AMOALU.scala 17:51]
  wire [3:0] s1_mask_xwr_hi_2; // @[AMOALU.scala 17:46]
  wire [3:0] s1_mask_xwr_lo_2; // @[AMOALU.scala 18:22]
  wire [7:0] s1_mask_xwr; // @[Cat.scala 30:58]
  wire  s1_hazard_hi_hi_hi_2; // @[DCache.scala 1149:66]
  wire  s1_hazard_hi_hi_lo_2; // @[DCache.scala 1149:66]
  wire  s1_hazard_hi_lo_hi_2; // @[DCache.scala 1149:66]
  wire  s1_hazard_hi_lo_lo_2; // @[DCache.scala 1149:66]
  wire  s1_hazard_lo_hi_hi_2; // @[DCache.scala 1149:66]
  wire  s1_hazard_lo_hi_lo_2; // @[DCache.scala 1149:66]
  wire  s1_hazard_lo_lo_hi_2; // @[DCache.scala 1149:66]
  wire  s1_hazard_lo_lo_lo_2; // @[DCache.scala 1149:66]
  wire [7:0] _s1_hazard_T_21; // @[Cat.scala 30:58]
  wire  s1_hazard_hi_hi_hi_3; // @[Bitwise.scala 26:51]
  wire  s1_hazard_hi_hi_lo_3; // @[Bitwise.scala 26:51]
  wire  s1_hazard_hi_lo_hi_3; // @[Bitwise.scala 26:51]
  wire  s1_hazard_hi_lo_lo_3; // @[Bitwise.scala 26:51]
  wire  s1_hazard_lo_hi_hi_3; // @[Bitwise.scala 26:51]
  wire  s1_hazard_lo_hi_lo_3; // @[Bitwise.scala 26:51]
  wire  s1_hazard_lo_lo_hi_3; // @[Bitwise.scala 26:51]
  wire  s1_hazard_lo_lo_lo_3; // @[Bitwise.scala 26:51]
  wire [7:0] _s1_hazard_T_22; // @[Cat.scala 30:58]
  wire [7:0] _s1_hazard_T_23; // @[DCache.scala 533:38]
  wire  _s1_hazard_T_24; // @[DCache.scala 533:66]
  wire [7:0] _s1_hazard_T_25; // @[DCache.scala 533:77]
  wire  _s1_hazard_T_26; // @[DCache.scala 533:92]
  wire  _s1_hazard_T_27; // @[DCache.scala 533:8]
  wire  _s1_hazard_T_28; // @[DCache.scala 532:65]
  wire  _s1_hazard_T_29; // @[DCache.scala 535:27]
  reg  pstore2_valid; // @[DCache.scala 472:30]
  reg [31:0] _RAND_36;
  reg [39:0] pstore2_addr; // @[Reg.scala 15:16]
  reg [63:0] _RAND_37;
  wire  _s1_hazard_T_32; // @[DCache.scala 532:31]
  reg [7:0] mask; // @[DCache.scala 502:19]
  reg [31:0] _RAND_38;
  wire  s1_hazard_hi_hi_hi_4; // @[DCache.scala 1149:66]
  wire  s1_hazard_hi_hi_lo_4; // @[DCache.scala 1149:66]
  wire  s1_hazard_hi_lo_hi_4; // @[DCache.scala 1149:66]
  wire  s1_hazard_hi_lo_lo_4; // @[DCache.scala 1149:66]
  wire  s1_hazard_lo_hi_hi_4; // @[DCache.scala 1149:66]
  wire  s1_hazard_lo_hi_lo_4; // @[DCache.scala 1149:66]
  wire  s1_hazard_lo_lo_hi_4; // @[DCache.scala 1149:66]
  wire  s1_hazard_lo_lo_lo_4; // @[DCache.scala 1149:66]
  wire [7:0] _s1_hazard_T_41; // @[Cat.scala 30:58]
  wire  s1_hazard_hi_hi_hi_5; // @[Bitwise.scala 26:51]
  wire  s1_hazard_hi_hi_lo_5; // @[Bitwise.scala 26:51]
  wire  s1_hazard_hi_lo_hi_5; // @[Bitwise.scala 26:51]
  wire  s1_hazard_hi_lo_lo_5; // @[Bitwise.scala 26:51]
  wire  s1_hazard_lo_hi_hi_5; // @[Bitwise.scala 26:51]
  wire  s1_hazard_lo_hi_lo_5; // @[Bitwise.scala 26:51]
  wire  s1_hazard_lo_lo_hi_5; // @[Bitwise.scala 26:51]
  wire  s1_hazard_lo_lo_lo_5; // @[Bitwise.scala 26:51]
  wire [7:0] _s1_hazard_T_42; // @[Cat.scala 30:58]
  wire [7:0] _s1_hazard_T_53; // @[DCache.scala 533:38]
  wire  _s1_hazard_T_54; // @[DCache.scala 533:66]
  wire [7:0] _s1_hazard_T_55; // @[DCache.scala 533:77]
  wire  _s1_hazard_T_56; // @[DCache.scala 533:92]
  wire  _s1_hazard_T_57; // @[DCache.scala 533:8]
  wire  _s1_hazard_T_58; // @[DCache.scala 532:65]
  wire  _s1_hazard_T_59; // @[DCache.scala 536:21]
  wire  s1_hazard; // @[DCache.scala 535:69]
  wire  s1_raw_hazard; // @[DCache.scala 537:31]
  wire  _T_262; // @[DCache.scala 542:18]
  wire [5:0] _s2_valid_no_xcpt_T; // @[DCache.scala 303:54]
  wire  _s2_valid_no_xcpt_T_1; // @[DCache.scala 303:61]
  wire  s2_valid_no_xcpt; // @[DCache.scala 303:35]
  reg  s2_not_nacked_in_s1; // @[DCache.scala 306:36]
  reg [31:0] _RAND_39;
  wire  s2_valid_masked; // @[DCache.scala 308:42]
  wire  _s2_valid_hit_maybe_flush_pre_data_ecc_and_waw_T_1; // @[DCache.scala 368:71]
  wire  _c_cat_T_45; // @[Consts.scala 83:54]
  wire  _c_cat_T_46; // @[Consts.scala 83:47]
  wire  _c_cat_T_47; // @[Consts.scala 83:71]
  wire  c_cat_lo; // @[Consts.scala 83:64]
  reg [1:0] s2_hit_state_state; // @[Reg.scala 15:16]
  reg [31:0] _RAND_40;
  wire [3:0] _T_71; // @[Cat.scala 30:58]
  wire  _T_117; // @[Misc.scala 48:20]
  wire  _T_114; // @[Misc.scala 48:20]
  wire  _T_111; // @[Misc.scala 48:20]
  wire  _T_108; // @[Misc.scala 48:20]
  wire  _T_105; // @[Misc.scala 48:20]
  wire  _T_102; // @[Misc.scala 48:20]
  wire  _T_99; // @[Misc.scala 48:20]
  wire  _T_96; // @[Misc.scala 48:20]
  wire  _T_93; // @[Misc.scala 48:20]
  wire  _T_90; // @[Misc.scala 48:20]
  wire  _T_87; // @[Misc.scala 48:20]
  wire  _T_84; // @[Misc.scala 48:20]
  wire  _T_103; // @[Misc.scala 34:9]
  wire  _T_106; // @[Misc.scala 34:9]
  wire  _T_109; // @[Misc.scala 34:9]
  wire  _T_112; // @[Misc.scala 34:9]
  wire  _T_115; // @[Misc.scala 34:9]
  wire  s2_hit; // @[Misc.scala 34:9]
  wire  s2_valid_hit_maybe_flush_pre_data_ecc_and_waw; // @[DCache.scala 368:89]
  wire  _s2_read_T; // @[Consts.scala 81:31]
  wire  _s2_read_T_2; // @[Consts.scala 81:41]
  wire  _s2_read_T_4; // @[Consts.scala 81:58]
  wire  s2_read; // @[Consts.scala 81:75]
  wire  s2_readwrite; // @[DCache.scala 325:30]
  wire  s2_valid_hit_pre_data_ecc_and_waw; // @[DCache.scala 389:89]
  wire [1:0] _T_86; // @[Misc.scala 34:36]
  wire [1:0] _T_89; // @[Misc.scala 34:36]
  wire [1:0] _T_92; // @[Misc.scala 34:36]
  wire [1:0] _T_95; // @[Misc.scala 34:36]
  wire [1:0] _T_98; // @[Misc.scala 34:36]
  wire [1:0] _T_101; // @[Misc.scala 34:36]
  wire [1:0] _T_104; // @[Misc.scala 34:36]
  wire [1:0] _T_107; // @[Misc.scala 34:36]
  wire [1:0] _T_110; // @[Misc.scala 34:36]
  wire [1:0] _T_113; // @[Misc.scala 34:36]
  wire [1:0] _T_116; // @[Misc.scala 34:36]
  wire [1:0] s2_grow_param; // @[Misc.scala 34:36]
  wire  _s2_update_meta_T; // @[Metadata.scala 45:46]
  wire  s2_update_meta; // @[Metadata.scala 46:40]
  wire  _T_241; // @[DCache.scala 417:62]
  wire  _T_242; // @[DCache.scala 417:24]
  wire  s1_readwrite; // @[DCache.scala 190:30]
  wire  _s1_flush_line_T; // @[DCache.scala 192:34]
  wire  s1_flush_line; // @[DCache.scala 192:50]
  wire  _s1_cmd_uses_tlb_T; // @[DCache.scala 248:38]
  wire  _s1_cmd_uses_tlb_T_1; // @[DCache.scala 248:69]
  wire  s1_cmd_uses_tlb; // @[DCache.scala 248:55]
  wire  _T_13; // @[DCache.scala 254:39]
  wire  _T_14; // @[DCache.scala 254:58]
  wire  _GEN_117; // @[DCache.scala 417:82]
  wire  _GEN_141; // @[DCache.scala 542:36]
  wire  _GEN_283; // @[DCache.scala 810:24]
  wire  s1_nack; // @[DCache.scala 795:21]
  wire  s1_valid_not_nacked; // @[DCache.scala 167:38]
  wire  s0_clk_en; // @[DCache.scala 170:40]
  wire [33:0] s0_req_addr_hi; // @[DCache.scala 173:47]
  wire [5:0] s0_req_addr_lo; // @[DCache.scala 173:84]
  wire [39:0] s0_req_addr; // @[Cat.scala 30:58]
  wire  s0_req_phys; // @[DCache.scala 175:34]
  reg [6:0] s1_req_tag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_41;
  reg  s1_req_signed; // @[Reg.scala 15:16]
  reg [31:0] _RAND_42;
  reg [39:0] s1_tlb_req_vaddr; // @[Reg.scala 15:16]
  reg [63:0] _RAND_43;
  reg  s1_tlb_req_passthrough; // @[Reg.scala 15:16]
  reg [31:0] _RAND_44;
  reg [1:0] s1_tlb_req_size; // @[Reg.scala 15:16]
  reg [31:0] _RAND_45;
  reg [4:0] s1_tlb_req_cmd; // @[Reg.scala 15:16]
  reg [31:0] _RAND_46;
  wire  s1_sfence; // @[DCache.scala 191:30]
  reg  s1_flush_valid; // @[DCache.scala 193:27]
  reg [31:0] _RAND_47;
  reg  cached_grant_wait; // @[DCache.scala 201:30]
  reg [31:0] _RAND_48;
  reg  resetting; // @[DCache.scala 202:26]
  reg [31:0] _RAND_49;
  reg [7:0] flushCounter; // @[DCache.scala 203:25]
  reg [31:0] _RAND_50;
  reg [3:0] refill_way; // @[DCache.scala 207:23]
  reg [31:0] _RAND_51;
  wire  inWriteback; // @[package.scala 72:59]
  wire  _io_cpu_req_ready_T; // @[DCache.scala 211:38]
  wire  _io_cpu_req_ready_T_2; // @[DCache.scala 211:51]
  wire  _io_cpu_req_ready_T_4; // @[DCache.scala 211:73]
  reg  uncachedInFlight_0; // @[DCache.scala 214:33]
  reg [31:0] _RAND_52;
  reg [39:0] uncachedReqs_0_addr; // @[DCache.scala 215:25]
  reg [63:0] _RAND_53;
  reg [6:0] uncachedReqs_0_tag; // @[DCache.scala 215:25]
  reg [31:0] _RAND_54;
  reg [1:0] uncachedReqs_0_size; // @[DCache.scala 215:25]
  reg [31:0] _RAND_55;
  reg  uncachedReqs_0_signed; // @[DCache.scala 215:25]
  reg [31:0] _RAND_56;
  wire  _s0_read_T; // @[Consts.scala 81:31]
  wire  _s0_read_T_1; // @[Consts.scala 81:48]
  wire  _s0_read_T_2; // @[Consts.scala 81:41]
  wire  _s0_read_T_3; // @[Consts.scala 81:65]
  wire  _s0_read_T_4; // @[Consts.scala 81:58]
  wire  _s0_read_T_5; // @[package.scala 15:47]
  wire  _s0_read_T_6; // @[package.scala 15:47]
  wire  _s0_read_T_7; // @[package.scala 15:47]
  wire  _s0_read_T_8; // @[package.scala 15:47]
  wire  _s0_read_T_9; // @[package.scala 72:59]
  wire  _s0_read_T_10; // @[package.scala 72:59]
  wire  _s0_read_T_11; // @[package.scala 72:59]
  wire  _s0_read_T_12; // @[package.scala 15:47]
  wire  _s0_read_T_13; // @[package.scala 15:47]
  wire  _s0_read_T_14; // @[package.scala 15:47]
  wire  _s0_read_T_15; // @[package.scala 15:47]
  wire  _s0_read_T_16; // @[package.scala 15:47]
  wire  _s0_read_T_17; // @[package.scala 72:59]
  wire  _s0_read_T_18; // @[package.scala 72:59]
  wire  _s0_read_T_19; // @[package.scala 72:59]
  wire  _s0_read_T_20; // @[package.scala 72:59]
  wire  _s0_read_T_21; // @[Consts.scala 79:44]
  wire  s0_read; // @[Consts.scala 81:75]
  wire  _dataArb_io_in_3_valid_res_T; // @[package.scala 15:47]
  wire  _dataArb_io_in_3_valid_res_T_1; // @[package.scala 15:47]
  wire  _dataArb_io_in_3_valid_res_T_2; // @[package.scala 72:59]
  wire  res; // @[DCache.scala 1153:15]
  wire  _dataArb_io_in_3_valid_T_24; // @[Consts.scala 82:49]
  wire  _dataArb_io_in_3_valid_T_25; // @[Consts.scala 82:42]
  wire  _dataArb_io_in_3_valid_T_27; // @[Consts.scala 82:59]
  wire  _dataArb_io_in_3_valid_T_45; // @[Consts.scala 82:76]
  wire  _dataArb_io_in_3_valid_T_49; // @[DCache.scala 1159:23]
  wire  _dataArb_io_in_3_valid_T_50; // @[DCache.scala 1158:21]
  wire  _dataArb_io_in_3_valid_T_52; // @[DCache.scala 1154:28]
  wire  _dataArb_io_in_3_valid_T_54; // @[DCache.scala 1154:11]
  wire  _dataArb_io_in_3_valid_T_56; // @[DCache.scala 220:46]
  wire [27:0] dataArb_io_in_3_bits_addr_hi; // @[DCache.scala 223:89]
  wire [11:0] dataArb_io_in_3_bits_addr_lo; // @[DCache.scala 223:120]
  wire [39:0] _dataArb_io_in_3_bits_addr_T; // @[Cat.scala 30:58]
  wire  _T_4; // @[DCache.scala 236:33]
  wire  _GEN_28; // @[DCache.scala 236:45]
  wire  _s1_did_read_T_51; // @[DCache.scala 237:75]
  wire  _s1_did_read_T_52; // @[DCache.scala 237:54]
  reg  s1_did_read; // @[Reg.scala 15:16]
  reg [31:0] _RAND_57;
  reg  s1_read_mask; // @[Reg.scala 15:16]
  reg [31:0] _RAND_58;
  wire  _GEN_31; // @[DCache.scala 245:34]
  wire  _T_8; // @[DCache.scala 253:27]
  wire  _T_10; // @[DCache.scala 253:53]
  wire  _GEN_32; // @[DCache.scala 253:79]
  wire [19:0] s1_paddr_hi; // @[DCache.scala 269:99]
  wire [31:0] s1_paddr; // @[Cat.scala 30:58]
  wire [21:0] _WIRE_2;
  wire [19:0] s1_meta_uncorrected_0_tag; // @[DCache.scala 286:80]
  wire [1:0] s1_meta_uncorrected_0_coh_state; // @[DCache.scala 286:80]
  wire [21:0] _WIRE_3;
  wire [19:0] s1_meta_uncorrected_1_tag; // @[DCache.scala 286:80]
  wire [1:0] s1_meta_uncorrected_1_coh_state; // @[DCache.scala 286:80]
  wire [21:0] _WIRE_4;
  wire [19:0] s1_meta_uncorrected_2_tag; // @[DCache.scala 286:80]
  wire [1:0] s1_meta_uncorrected_2_coh_state; // @[DCache.scala 286:80]
  wire [21:0] _WIRE_5;
  wire [19:0] s1_meta_uncorrected_3_tag; // @[DCache.scala 286:80]
  wire [1:0] s1_meta_uncorrected_3_coh_state; // @[DCache.scala 286:80]
  wire [19:0] s1_tag; // @[DCache.scala 287:29]
  wire  _T_32; // @[Metadata.scala 49:45]
  wire  _T_33; // @[DCache.scala 288:83]
  wire  lo_lo; // @[DCache.scala 288:74]
  wire  _T_34; // @[Metadata.scala 49:45]
  wire  _T_35; // @[DCache.scala 288:83]
  wire  lo_hi; // @[DCache.scala 288:74]
  wire  _T_36; // @[Metadata.scala 49:45]
  wire  _T_37; // @[DCache.scala 288:83]
  wire  hi_lo; // @[DCache.scala 288:74]
  wire  _T_38; // @[Metadata.scala 49:45]
  wire  _T_39; // @[DCache.scala 288:83]
  wire  hi_hi; // @[DCache.scala 288:74]
  wire [3:0] s1_meta_hit_way; // @[Cat.scala 30:58]
  wire  _T_42; // @[DCache.scala 290:59]
  wire [1:0] _T_43; // @[DCache.scala 290:41]
  wire  _T_46; // @[DCache.scala 290:59]
  wire [1:0] _T_47; // @[DCache.scala 290:41]
  wire  _T_50; // @[DCache.scala 290:59]
  wire [1:0] _T_51; // @[DCache.scala 290:41]
  wire  _T_54; // @[DCache.scala 290:59]
  wire [1:0] _T_55; // @[DCache.scala 290:41]
  wire [1:0] _T_56; // @[DCache.scala 291:19]
  wire [1:0] _T_57; // @[DCache.scala 291:19]
  wire [1:0] s1_meta_hit_state_state; // @[DCache.scala 291:19]
  wire  s2_hit_valid; // @[Metadata.scala 49:45]
  reg [3:0] s2_hit_way; // @[Reg.scala 15:16]
  reg [31:0] _RAND_59;
  reg [1:0] s2_victim_way_r; // @[Reg.scala 15:16]
  reg [31:0] _RAND_60;
  wire [3:0] s2_victim_way; // @[OneHot.scala 58:35]
  wire [3:0] s2_victim_or_hit_way; // @[DCache.scala 403:33]
  reg [3:0] s2_probe_way; // @[Reg.scala 15:16]
  reg [31:0] _RAND_61;
  wire [3:0] releaseWay; // @[DCache.scala 834:102]
  wire [3:0] s1_data_way_x35; // @[DCache.scala 294:61]
  wire [7:0] tl_d_data_encoded_lo_lo_lo; // @[package.scala 202:50]
  wire [7:0] tl_d_data_encoded_lo_lo_hi; // @[package.scala 202:50]
  wire [7:0] tl_d_data_encoded_lo_hi_lo; // @[package.scala 202:50]
  wire [7:0] tl_d_data_encoded_lo_hi_hi; // @[package.scala 202:50]
  wire [7:0] tl_d_data_encoded_hi_lo_lo; // @[package.scala 202:50]
  wire [7:0] tl_d_data_encoded_hi_lo_hi; // @[package.scala 202:50]
  wire [7:0] tl_d_data_encoded_hi_hi_lo; // @[package.scala 202:50]
  wire [7:0] tl_d_data_encoded_hi_hi_hi; // @[package.scala 202:50]
  wire [31:0] tl_d_data_encoded_lo; // @[Cat.scala 30:58]
  wire [31:0] tl_d_data_encoded_hi; // @[Cat.scala 30:58]
  wire [63:0] _tl_d_data_encoded_T; // @[Cat.scala 30:58]
  wire  _T_61; // @[DCache.scala 300:28]
  wire  _T_65; // @[DCache.scala 300:93]
  wire  _T_66; // @[DCache.scala 300:53]
  wire  _T_68; // @[DCache.scala 300:9]
  wire  s2_valid_x37; // @[DCache.scala 302:43]
  reg [39:0] s2_req_addr; // @[DCache.scala 310:19]
  reg [63:0] _RAND_62;
  reg [6:0] s2_req_tag; // @[DCache.scala 310:19]
  reg [31:0] _RAND_63;
  reg [1:0] s2_req_size; // @[DCache.scala 310:19]
  reg [31:0] _RAND_64;
  reg  s2_req_signed; // @[DCache.scala 310:19]
  reg [31:0] _RAND_65;
  wire  _s2_cmd_flush_all_T; // @[DCache.scala 311:37]
  wire  s2_cmd_flush_line; // @[DCache.scala 312:54]
  reg  s2_tlb_xcpt_pf_ld; // @[DCache.scala 313:24]
  reg [31:0] _RAND_66;
  reg  s2_tlb_xcpt_pf_st; // @[DCache.scala 313:24]
  reg [31:0] _RAND_67;
  reg  s2_tlb_xcpt_ae_ld; // @[DCache.scala 313:24]
  reg [31:0] _RAND_68;
  reg  s2_tlb_xcpt_ae_st; // @[DCache.scala 313:24]
  reg [31:0] _RAND_69;
  reg  s2_tlb_xcpt_ma_ld; // @[DCache.scala 313:24]
  reg [31:0] _RAND_70;
  reg  s2_tlb_xcpt_ma_st; // @[DCache.scala 313:24]
  reg [31:0] _RAND_71;
  reg  s2_pma_cacheable; // @[DCache.scala 314:19]
  reg [31:0] _RAND_72;
  wire  _T_70; // @[DCache.scala 316:29]
  wire  _s2_pma_T_cacheable; // @[DCache.scala 320:18]
  reg [39:0] s2_vaddr_r; // @[Reg.scala 15:16]
  reg [63:0] _RAND_73;
  wire [27:0] s2_vaddr_hi; // @[DCache.scala 322:81]
  wire [11:0] s2_vaddr_lo; // @[DCache.scala 322:103]
  wire [39:0] s2_vaddr; // @[Cat.scala 30:58]
  reg  s2_flush_valid_pre_tag_ecc; // @[DCache.scala 326:43]
  reg [31:0] _RAND_74;
  wire  s1_meta_clk_en; // @[DCache.scala 328:62]
  reg [21:0] s2_meta_corrected_r; // @[Reg.scala 15:16]
  reg [31:0] _RAND_75;
  wire [19:0] s2_meta_corrected_0_tag; // @[DCache.scala 332:99]
  wire [1:0] s2_meta_corrected_0_coh_state; // @[DCache.scala 332:99]
  reg [21:0] s2_meta_corrected_r_1; // @[Reg.scala 15:16]
  reg [31:0] _RAND_76;
  wire [19:0] s2_meta_corrected_1_tag; // @[DCache.scala 332:99]
  wire [1:0] s2_meta_corrected_1_coh_state; // @[DCache.scala 332:99]
  reg [21:0] s2_meta_corrected_r_2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_77;
  wire [19:0] s2_meta_corrected_2_tag; // @[DCache.scala 332:99]
  wire [1:0] s2_meta_corrected_2_coh_state; // @[DCache.scala 332:99]
  reg [21:0] s2_meta_corrected_r_3; // @[Reg.scala 15:16]
  reg [31:0] _RAND_78;
  wire [19:0] s2_meta_corrected_3_tag; // @[DCache.scala 332:99]
  wire [1:0] s2_meta_corrected_3_coh_state; // @[DCache.scala 332:99]
  wire  s2_flush_valid; // @[DCache.scala 334:51]
  wire  _s2_data_en_T; // @[DCache.scala 337:23]
  wire  en; // @[DCache.scala 337:38]
  wire  _s2_data_word_en_T; // @[DCache.scala 338:63]
  wire  word_en; // @[DCache.scala 338:22]
  wire [63:0] s1_all_data_ways_0; // @[DCache.scala 296:29 DCache.scala 296:29]
  wire [63:0] s1_all_data_ways_1; // @[DCache.scala 296:29 DCache.scala 296:29]
  wire [63:0] s1_all_data_ways_2; // @[DCache.scala 296:29 DCache.scala 296:29]
  wire [63:0] s1_all_data_ways_3; // @[DCache.scala 296:29 DCache.scala 296:29]
  wire  s1_word_en; // @[DCache.scala 348:27]
  wire  grantIsUncachedData; // @[package.scala 15:47]
  reg  blockUncachedGrant; // @[DCache.scala 721:33]
  reg [31:0] _RAND_79;
  wire  _T_293; // @[DCache.scala 723:54]
  wire  _T_294; // @[DCache.scala 723:31]
  wire  grantIsRefill; // @[DCache.scala 637:29]
  wire  _T_292; // @[DCache.scala 693:23]
  wire  _grantIsCached_T; // @[package.scala 15:47]
  wire  grantIsCached; // @[package.scala 72:59]
  reg [8:0] counter; // @[Edges.scala 228:27]
  reg [31:0] _RAND_80;
  wire  d_first; // @[Edges.scala 230:25]
  wire  _bundleOut_0_d_ready_T_1; // @[DCache.scala 642:50]
  wire  canAcceptCachedGrant; // @[DCache.scala 641:30]
  wire  _bundleOut_0_d_ready_T_2; // @[DCache.scala 642:69]
  wire  _bundleOut_0_d_ready_T_3; // @[DCache.scala 642:24]
  wire  _GEN_233; // @[DCache.scala 693:51]
  wire  tl_out__d_ready; // @[DCache.scala 723:68]
  wire  _T_271; // @[Decoupled.scala 40:37]
  wire  _T_267; // @[package.scala 15:47]
  wire  _T_269; // @[package.scala 72:59]
  wire  _T_268; // @[package.scala 15:47]
  wire  grantIsUncached; // @[package.scala 72:59]
  wire [4:0] _GEN_189; // @[DCache.scala 662:34]
  wire [4:0] _GEN_198; // @[DCache.scala 655:35]
  wire [4:0] _GEN_211; // @[DCache.scala 646:26]
  wire [4:0] s1_data_way; // @[DCache.scala 645:26]
  wire [4:0] _s2_data_T_1; // @[DCache.scala 350:28]
  wire [63:0] _s2_data_T_7; // @[Mux.scala 27:72]
  wire [63:0] _s2_data_T_8; // @[Mux.scala 27:72]
  wire [63:0] _s2_data_T_9; // @[Mux.scala 27:72]
  wire [63:0] _s2_data_T_10; // @[Mux.scala 27:72]
  wire [63:0] _s2_data_T_11; // @[Mux.scala 27:72]
  wire [63:0] _s2_data_T_12; // @[Mux.scala 27:72]
  wire [63:0] _s2_data_T_13; // @[Mux.scala 27:72]
  wire [63:0] _s2_data_T_14; // @[Mux.scala 27:72]
  wire [63:0] _s2_data_T_15; // @[Mux.scala 27:72]
  reg [63:0] s2_data; // @[Reg.scala 15:16]
  reg [63:0] _RAND_81;
  wire [7:0] s2_data_uncorrected_lo_lo_lo; // @[package.scala 202:50]
  wire [7:0] s2_data_uncorrected_lo_lo_hi; // @[package.scala 202:50]
  wire [7:0] s2_data_uncorrected_lo_hi_lo; // @[package.scala 202:50]
  wire [7:0] s2_data_uncorrected_lo_hi_hi; // @[package.scala 202:50]
  wire [7:0] s2_data_uncorrected_hi_lo_lo; // @[package.scala 202:50]
  wire [7:0] s2_data_uncorrected_hi_lo_hi; // @[package.scala 202:50]
  wire [7:0] s2_data_uncorrected_hi_hi_lo; // @[package.scala 202:50]
  wire [7:0] s2_data_uncorrected_hi_hi_hi; // @[package.scala 202:50]
  wire [31:0] s2_data_corrected_lo; // @[Cat.scala 30:58]
  wire [31:0] s2_data_corrected_hi; // @[Cat.scala 30:58]
  wire [63:0] s2_data_corrected; // @[Cat.scala 30:58]
  wire  s2_valid_flush_line; // @[DCache.scala 390:75]
  wire  _s2_valid_miss_T; // @[DCache.scala 394:39]
  wire  _s2_valid_miss_T_2; // @[DCache.scala 394:55]
  wire  s2_valid_miss; // @[DCache.scala 394:73]
  wire  s2_uncached; // @[DCache.scala 395:21]
  wire  _s2_valid_cached_miss_T_1; // @[DCache.scala 396:44]
  wire  _s2_valid_cached_miss_T_2; // @[DCache.scala 396:88]
  wire  s2_valid_cached_miss; // @[DCache.scala 396:60]
  wire  _s2_want_victimize_T; // @[DCache.scala 398:79]
  wire  s2_want_victimize; // @[DCache.scala 398:125]
  wire  _s2_valid_uncached_pending_T; // @[DCache.scala 401:49]
  wire  _s2_valid_uncached_pending_T_1; // @[DCache.scala 401:92]
  wire  s2_valid_uncached_pending; // @[DCache.scala 401:64]
  wire [1:0] s1_victim_way; // @[package.scala 154:13]
  wire [19:0] _s2_victim_tag_T_6; // @[Mux.scala 27:72]
  wire [19:0] _s2_victim_tag_T_7; // @[Mux.scala 27:72]
  wire [19:0] _s2_victim_tag_T_8; // @[Mux.scala 27:72]
  wire [19:0] _s2_victim_tag_T_9; // @[Mux.scala 27:72]
  wire [19:0] _s2_victim_tag_T_10; // @[Mux.scala 27:72]
  wire [19:0] _s2_victim_tag_T_11; // @[Mux.scala 27:72]
  wire [19:0] _s2_victim_tag_T_12; // @[Mux.scala 27:72]
  wire [1:0] _s2_victim_tag_T_13; // @[Mux.scala 27:72]
  wire [1:0] _s2_victim_tag_T_14; // @[Mux.scala 27:72]
  wire [1:0] _s2_victim_tag_T_15; // @[Mux.scala 27:72]
  wire [1:0] _s2_victim_tag_T_16; // @[Mux.scala 27:72]
  wire [1:0] _s2_victim_tag_T_17; // @[Mux.scala 27:72]
  wire [1:0] _s2_victim_tag_T_18; // @[Mux.scala 27:72]
  wire [1:0] _s2_victim_tag_T_19; // @[Mux.scala 27:72]
  wire [19:0] s2_victim_tag; // @[DCache.scala 404:26]
  wire [1:0] s2_victim_state_state; // @[DCache.scala 405:28]
  wire [2:0] _T_133; // @[Misc.scala 37:36]
  wire [2:0] _T_137; // @[Misc.scala 37:36]
  wire [2:0] _T_141; // @[Misc.scala 37:36]
  wire [2:0] _T_145; // @[Misc.scala 37:36]
  wire [2:0] _T_149; // @[Misc.scala 37:36]
  wire [2:0] _T_153; // @[Misc.scala 37:36]
  wire [1:0] _T_154; // @[Misc.scala 37:63]
  wire [2:0] _T_157; // @[Misc.scala 37:36]
  wire [1:0] _T_158; // @[Misc.scala 37:63]
  wire [2:0] _T_161; // @[Misc.scala 37:36]
  wire [1:0] _T_162; // @[Misc.scala 37:63]
  wire [2:0] _T_165; // @[Misc.scala 37:36]
  wire [1:0] _T_166; // @[Misc.scala 37:63]
  wire [2:0] _T_169; // @[Misc.scala 37:36]
  wire [1:0] _T_170; // @[Misc.scala 37:63]
  wire [2:0] _T_173; // @[Misc.scala 37:36]
  wire [1:0] _T_174; // @[Misc.scala 37:63]
  wire [2:0] s2_report_param; // @[Misc.scala 37:36]
  wire [1:0] probeNewCoh_state; // @[Misc.scala 37:63]
  wire [3:0] _T_182; // @[Cat.scala 30:58]
  wire  _T_195; // @[Misc.scala 55:20]
  wire [2:0] _T_197; // @[Misc.scala 37:36]
  wire  _T_199; // @[Misc.scala 55:20]
  wire [2:0] _T_201; // @[Misc.scala 37:36]
  wire  _T_203; // @[Misc.scala 55:20]
  wire [2:0] _T_205; // @[Misc.scala 37:36]
  wire  _T_207; // @[Misc.scala 55:20]
  wire [2:0] _T_209; // @[Misc.scala 37:36]
  wire  _T_211; // @[Misc.scala 55:20]
  wire  _T_212; // @[Misc.scala 37:9]
  wire [2:0] _T_213; // @[Misc.scala 37:36]
  wire  _T_215; // @[Misc.scala 55:20]
  wire  _T_216; // @[Misc.scala 37:9]
  wire [2:0] _T_217; // @[Misc.scala 37:36]
  wire [1:0] _T_218; // @[Misc.scala 37:63]
  wire  _T_219; // @[Misc.scala 55:20]
  wire  _T_220; // @[Misc.scala 37:9]
  wire [2:0] _T_221; // @[Misc.scala 37:36]
  wire [1:0] _T_222; // @[Misc.scala 37:63]
  wire  _T_223; // @[Misc.scala 55:20]
  wire  _T_224; // @[Misc.scala 37:9]
  wire [2:0] _T_225; // @[Misc.scala 37:36]
  wire [1:0] _T_226; // @[Misc.scala 37:63]
  wire  _T_227; // @[Misc.scala 55:20]
  wire  _T_228; // @[Misc.scala 37:9]
  wire [2:0] _T_229; // @[Misc.scala 37:36]
  wire [1:0] _T_230; // @[Misc.scala 37:63]
  wire  _T_231; // @[Misc.scala 55:20]
  wire  _T_232; // @[Misc.scala 37:9]
  wire [2:0] _T_233; // @[Misc.scala 37:36]
  wire [1:0] _T_234; // @[Misc.scala 37:63]
  wire  _T_235; // @[Misc.scala 55:20]
  wire  _T_236; // @[Misc.scala 37:9]
  wire [2:0] _T_237; // @[Misc.scala 37:36]
  wire [1:0] _T_238; // @[Misc.scala 37:63]
  wire  _T_239; // @[Misc.scala 55:20]
  wire  s2_victim_dirty; // @[Misc.scala 37:9]
  wire [2:0] s2_shrink_param; // @[Misc.scala 37:36]
  wire [1:0] voluntaryNewCoh_state; // @[Misc.scala 37:63]
  wire  s2_dont_nack_uncached; // @[DCache.scala 411:57]
  wire  _s2_dont_nack_misc_T_10; // @[DCache.scala 415:17]
  wire  s2_dont_nack_misc; // @[DCache.scala 412:61]
  wire  _io_cpu_s2_nack_T_1; // @[DCache.scala 416:38]
  wire  _io_cpu_s2_nack_T_3; // @[DCache.scala 416:64]
  wire  _metaArb_io_in_1_valid_T; // @[DCache.scala 421:63]
  wire  _metaArb_io_in_1_valid_T_1; // @[DCache.scala 421:93]
  wire [11:0] metaArb_io_in_1_bits_addr_lo; // @[DCache.scala 425:98]
  wire [1:0] new_meta_coh_state; // @[DCache.scala 428:40]
  wire [11:0] metaArb_io_in_2_bits_addr_lo; // @[DCache.scala 437:80]
  wire [19:0] metaArb_io_in_2_bits_data_meta_tag; // @[HellaCache.scala 289:20 HellaCache.scala 290:14]
  wire  _lrscBackingOff_T; // @[DCache.scala 445:34]
  wire  lrscBackingOff; // @[DCache.scala 445:38]
  reg [33:0] lrscAddr; // @[DCache.scala 446:21]
  reg [63:0] _RAND_82;
  wire  lrscAddrMatch; // @[DCache.scala 447:32]
  wire  _s2_sc_fail_T; // @[DCache.scala 448:41]
  wire  s2_sc_fail; // @[DCache.scala 448:26]
  wire  _T_243; // @[DCache.scala 449:23]
  wire  _T_245; // @[DCache.scala 449:32]
  wire  _T_246; // @[DCache.scala 449:54]
  wire [6:0] _lrscCount_T_2; // @[DCache.scala 453:49]
  wire  _T_250; // @[DCache.scala 454:29]
  wire  _pstore1_cmd_T; // @[DCache.scala 463:63]
  reg [4:0] pstore1_cmd; // @[Reg.scala 15:16]
  reg [31:0] _RAND_83;
  reg [63:0] pstore1_data; // @[Reg.scala 15:16]
  reg [63:0] _RAND_84;
  reg [3:0] pstore1_way; // @[Reg.scala 15:16]
  reg [31:0] _RAND_85;
  wire  _pstore1_rmw_T_49; // @[DCache.scala 1159:23]
  wire  _pstore1_rmw_T_50; // @[DCache.scala 1158:21]
  reg  pstore1_rmw_r; // @[Reg.scala 15:16]
  reg [31:0] _RAND_86;
  wire  _pstore1_merge_T; // @[DCache.scala 461:46]
  wire  _pstore1_merge_T_2; // @[DCache.scala 461:58]
  wire  pstore_drain_opportunistic; // @[DCache.scala 473:36]
  reg  pstore_drain_on_miss_REG; // @[DCache.scala 474:56]
  reg [31:0] _RAND_87;
  wire  pstore_drain_on_miss; // @[DCache.scala 474:46]
  wire  pstore1_valid; // @[DCache.scala 478:38]
  wire  _pstore_drain_structural_T; // @[DCache.scala 480:54]
  wire  _pstore_drain_structural_T_1; // @[DCache.scala 480:85]
  wire  _pstore_drain_structural_T_2; // @[DCache.scala 480:98]
  wire  pstore_drain_structural; // @[DCache.scala 480:71]
  wire  _T_254; // @[DCache.scala 477:96]
  wire  _T_255; // @[DCache.scala 481:63]
  wire  _T_256; // @[DCache.scala 481:22]
  wire  _T_258; // @[DCache.scala 481:9]
  wire  _pstore_drain_T_7; // @[DCache.scala 489:41]
  wire  _pstore_drain_T_8; // @[DCache.scala 489:58]
  wire  _pstore_drain_T_9; // @[DCache.scala 489:107]
  wire  _pstore_drain_T_10; // @[DCache.scala 489:76]
  wire  pstore_drain; // @[DCache.scala 488:48]
  wire  _pstore1_held_T_8; // @[DCache.scala 492:71]
  wire  _pstore1_held_T_10; // @[DCache.scala 492:88]
  wire  _advance_pstore1_T_1; // @[DCache.scala 493:79]
  wire  advance_pstore1; // @[DCache.scala 493:61]
  wire  _pstore2_valid_T_1; // @[DCache.scala 494:34]
  wire  _pstore2_valid_T_2; // @[DCache.scala 494:51]
  reg [3:0] pstore2_way; // @[Reg.scala 15:16]
  reg [31:0] _RAND_88;
  wire [63:0] pstore1_storegen_data; // @[DCache.scala 957:27]
  reg [7:0] pstore2_storegen_data_lo_lo_lo; // @[Reg.scala 15:16]
  reg [31:0] _RAND_89;
  reg [7:0] pstore2_storegen_data_lo_lo_hi; // @[Reg.scala 15:16]
  reg [31:0] _RAND_90;
  reg [7:0] pstore2_storegen_data_lo_hi_lo; // @[Reg.scala 15:16]
  reg [31:0] _RAND_91;
  reg [7:0] pstore2_storegen_data_lo_hi_hi; // @[Reg.scala 15:16]
  reg [31:0] _RAND_92;
  reg [7:0] pstore2_storegen_data_hi_lo_lo; // @[Reg.scala 15:16]
  reg [31:0] _RAND_93;
  reg [7:0] pstore2_storegen_data_hi_lo_hi; // @[Reg.scala 15:16]
  reg [31:0] _RAND_94;
  reg [7:0] pstore2_storegen_data_hi_hi_lo; // @[Reg.scala 15:16]
  reg [31:0] _RAND_95;
  reg [7:0] pstore2_storegen_data_hi_hi_hi; // @[Reg.scala 15:16]
  reg [31:0] _RAND_96;
  wire [63:0] pstore2_storegen_data; // @[Cat.scala 30:58]
  wire [39:0] _dataArb_io_in_0_bits_addr_T; // @[DCache.scala 520:36]
  wire [63:0] _dataArb_io_in_0_bits_wdata_T; // @[DCache.scala 522:63]
  wire [7:0] dataArb_io_in_0_bits_wdata_lo_lo_lo; // @[package.scala 202:50]
  wire [7:0] dataArb_io_in_0_bits_wdata_lo_lo_hi; // @[package.scala 202:50]
  wire [7:0] dataArb_io_in_0_bits_wdata_lo_hi_lo; // @[package.scala 202:50]
  wire [7:0] dataArb_io_in_0_bits_wdata_lo_hi_hi; // @[package.scala 202:50]
  wire [7:0] dataArb_io_in_0_bits_wdata_hi_lo_lo; // @[package.scala 202:50]
  wire [7:0] dataArb_io_in_0_bits_wdata_hi_lo_hi; // @[package.scala 202:50]
  wire [7:0] dataArb_io_in_0_bits_wdata_hi_hi_lo; // @[package.scala 202:50]
  wire [7:0] dataArb_io_in_0_bits_wdata_hi_hi_hi; // @[package.scala 202:50]
  wire [31:0] dataArb_io_in_0_bits_wdata_lo; // @[Cat.scala 30:58]
  wire [31:0] dataArb_io_in_0_bits_wdata_hi; // @[Cat.scala 30:58]
  wire [7:0] _dataArb_io_in_0_bits_eccMask_T; // @[DCache.scala 528:47]
  wire  dataArb_io_in_0_bits_eccMask_lo_lo_lo; // @[DCache.scala 1149:66]
  wire  dataArb_io_in_0_bits_eccMask_lo_lo_hi; // @[DCache.scala 1149:66]
  wire  dataArb_io_in_0_bits_eccMask_lo_hi_lo; // @[DCache.scala 1149:66]
  wire  dataArb_io_in_0_bits_eccMask_lo_hi_hi; // @[DCache.scala 1149:66]
  wire  dataArb_io_in_0_bits_eccMask_hi_lo_lo; // @[DCache.scala 1149:66]
  wire  dataArb_io_in_0_bits_eccMask_hi_lo_hi; // @[DCache.scala 1149:66]
  wire  dataArb_io_in_0_bits_eccMask_hi_hi_lo; // @[DCache.scala 1149:66]
  wire  dataArb_io_in_0_bits_eccMask_hi_hi_hi; // @[DCache.scala 1149:66]
  wire [3:0] dataArb_io_in_0_bits_eccMask_lo; // @[Cat.scala 30:58]
  wire [3:0] dataArb_io_in_0_bits_eccMask_hi; // @[Cat.scala 30:58]
  wire [1:0] _a_source_T_1; // @[DCache.scala 548:59]
  wire  a_source; // @[Mux.scala 47:69]
  wire [39:0] acquire_address; // @[DCache.scala 549:49]
  wire [22:0] a_mask; // @[DCache.scala 553:29]
  wire [2:0] _get_a_mask_sizeOH_T; // @[Misc.scala 201:34]
  wire [1:0] get_a_mask_sizeOH_shiftAmount; // @[OneHot.scala 64:49]
  wire [3:0] _get_a_mask_sizeOH_T_1; // @[OneHot.scala 65:12]
  wire [2:0] get_a_mask_sizeOH; // @[Misc.scala 201:81]
  wire  _get_a_mask_T; // @[Misc.scala 205:21]
  wire  get_a_mask_size; // @[Misc.scala 208:26]
  wire  get_a_mask_bit; // @[Misc.scala 209:26]
  wire  get_a_mask_nbit; // @[Misc.scala 210:20]
  wire  _get_a_mask_acc_T; // @[Misc.scala 214:38]
  wire  get_a_mask_acc; // @[Misc.scala 214:29]
  wire  _get_a_mask_acc_T_1; // @[Misc.scala 214:38]
  wire  get_a_mask_acc_1; // @[Misc.scala 214:29]
  wire  get_a_mask_size_1; // @[Misc.scala 208:26]
  wire  get_a_mask_bit_1; // @[Misc.scala 209:26]
  wire  get_a_mask_nbit_1; // @[Misc.scala 210:20]
  wire  get_a_mask_eq_2; // @[Misc.scala 213:27]
  wire  _get_a_mask_acc_T_2; // @[Misc.scala 214:38]
  wire  get_a_mask_acc_2; // @[Misc.scala 214:29]
  wire  get_a_mask_eq_3; // @[Misc.scala 213:27]
  wire  _get_a_mask_acc_T_3; // @[Misc.scala 214:38]
  wire  get_a_mask_acc_3; // @[Misc.scala 214:29]
  wire  get_a_mask_eq_4; // @[Misc.scala 213:27]
  wire  _get_a_mask_acc_T_4; // @[Misc.scala 214:38]
  wire  get_a_mask_acc_4; // @[Misc.scala 214:29]
  wire  get_a_mask_eq_5; // @[Misc.scala 213:27]
  wire  _get_a_mask_acc_T_5; // @[Misc.scala 214:38]
  wire  get_a_mask_acc_5; // @[Misc.scala 214:29]
  wire  get_a_mask_size_2; // @[Misc.scala 208:26]
  wire  get_a_mask_bit_2; // @[Misc.scala 209:26]
  wire  get_a_mask_nbit_2; // @[Misc.scala 210:20]
  wire  get_a_mask_eq_6; // @[Misc.scala 213:27]
  wire  _get_a_mask_acc_T_6; // @[Misc.scala 214:38]
  wire  get_a_mask_lo_lo_lo; // @[Misc.scala 214:29]
  wire  get_a_mask_eq_7; // @[Misc.scala 213:27]
  wire  _get_a_mask_acc_T_7; // @[Misc.scala 214:38]
  wire  get_a_mask_lo_lo_hi; // @[Misc.scala 214:29]
  wire  get_a_mask_eq_8; // @[Misc.scala 213:27]
  wire  _get_a_mask_acc_T_8; // @[Misc.scala 214:38]
  wire  get_a_mask_lo_hi_lo; // @[Misc.scala 214:29]
  wire  get_a_mask_eq_9; // @[Misc.scala 213:27]
  wire  _get_a_mask_acc_T_9; // @[Misc.scala 214:38]
  wire  get_a_mask_lo_hi_hi; // @[Misc.scala 214:29]
  wire  get_a_mask_eq_10; // @[Misc.scala 213:27]
  wire  _get_a_mask_acc_T_10; // @[Misc.scala 214:38]
  wire  get_a_mask_hi_lo_lo; // @[Misc.scala 214:29]
  wire  get_a_mask_eq_11; // @[Misc.scala 213:27]
  wire  _get_a_mask_acc_T_11; // @[Misc.scala 214:38]
  wire  get_a_mask_hi_lo_hi; // @[Misc.scala 214:29]
  wire  get_a_mask_eq_12; // @[Misc.scala 213:27]
  wire  _get_a_mask_acc_T_12; // @[Misc.scala 214:38]
  wire  get_a_mask_hi_hi_lo; // @[Misc.scala 214:29]
  wire  get_a_mask_eq_13; // @[Misc.scala 213:27]
  wire  _get_a_mask_acc_T_13; // @[Misc.scala 214:38]
  wire  get_a_mask_hi_hi_hi; // @[Misc.scala 214:29]
  wire [7:0] get_mask; // @[Cat.scala 30:58]
  wire  _atomics_T; // @[Mux.scala 80:60]
  wire [2:0] _atomics_T_1_opcode; // @[Mux.scala 80:57]
  wire [3:0] atomics_a_size; // @[Edges.scala 513:17 Edges.scala 516:15]
  wire [3:0] _atomics_T_1_size; // @[Mux.scala 80:57]
  wire  _atomics_T_1_source; // @[Mux.scala 80:57]
  wire [31:0] atomics_a_address; // @[Edges.scala 513:17 Edges.scala 518:15]
  wire [31:0] _atomics_T_1_address; // @[Mux.scala 80:57]
  wire [7:0] _atomics_T_1_mask; // @[Mux.scala 80:57]
  wire [63:0] _atomics_T_1_data; // @[Mux.scala 80:57]
  wire  _atomics_T_2; // @[Mux.scala 80:60]
  wire [2:0] _atomics_T_3_opcode; // @[Mux.scala 80:57]
  wire [2:0] _atomics_T_3_param; // @[Mux.scala 80:57]
  wire [3:0] _atomics_T_3_size; // @[Mux.scala 80:57]
  wire  _atomics_T_3_source; // @[Mux.scala 80:57]
  wire [31:0] _atomics_T_3_address; // @[Mux.scala 80:57]
  wire [7:0] _atomics_T_3_mask; // @[Mux.scala 80:57]
  wire [63:0] _atomics_T_3_data; // @[Mux.scala 80:57]
  wire  _atomics_T_4; // @[Mux.scala 80:60]
  wire [2:0] _atomics_T_5_opcode; // @[Mux.scala 80:57]
  wire [2:0] _atomics_T_5_param; // @[Mux.scala 80:57]
  wire [3:0] _atomics_T_5_size; // @[Mux.scala 80:57]
  wire  _atomics_T_5_source; // @[Mux.scala 80:57]
  wire [31:0] _atomics_T_5_address; // @[Mux.scala 80:57]
  wire [7:0] _atomics_T_5_mask; // @[Mux.scala 80:57]
  wire [63:0] _atomics_T_5_data; // @[Mux.scala 80:57]
  wire  _atomics_T_6; // @[Mux.scala 80:60]
  wire [2:0] _atomics_T_7_opcode; // @[Mux.scala 80:57]
  wire [2:0] _atomics_T_7_param; // @[Mux.scala 80:57]
  wire [3:0] _atomics_T_7_size; // @[Mux.scala 80:57]
  wire  _atomics_T_7_source; // @[Mux.scala 80:57]
  wire [31:0] _atomics_T_7_address; // @[Mux.scala 80:57]
  wire [7:0] _atomics_T_7_mask; // @[Mux.scala 80:57]
  wire [63:0] _atomics_T_7_data; // @[Mux.scala 80:57]
  wire  _atomics_T_8; // @[Mux.scala 80:60]
  wire [2:0] _atomics_T_9_opcode; // @[Mux.scala 80:57]
  wire [2:0] _atomics_T_9_param; // @[Mux.scala 80:57]
  wire [3:0] _atomics_T_9_size; // @[Mux.scala 80:57]
  wire  _atomics_T_9_source; // @[Mux.scala 80:57]
  wire [31:0] _atomics_T_9_address; // @[Mux.scala 80:57]
  wire [7:0] _atomics_T_9_mask; // @[Mux.scala 80:57]
  wire [63:0] _atomics_T_9_data; // @[Mux.scala 80:57]
  wire  _atomics_T_10; // @[Mux.scala 80:60]
  wire [2:0] _atomics_T_11_opcode; // @[Mux.scala 80:57]
  wire [2:0] _atomics_T_11_param; // @[Mux.scala 80:57]
  wire [3:0] _atomics_T_11_size; // @[Mux.scala 80:57]
  wire  _atomics_T_11_source; // @[Mux.scala 80:57]
  wire [31:0] _atomics_T_11_address; // @[Mux.scala 80:57]
  wire [7:0] _atomics_T_11_mask; // @[Mux.scala 80:57]
  wire [63:0] _atomics_T_11_data; // @[Mux.scala 80:57]
  wire  _atomics_T_12; // @[Mux.scala 80:60]
  wire [2:0] _atomics_T_13_opcode; // @[Mux.scala 80:57]
  wire [2:0] _atomics_T_13_param; // @[Mux.scala 80:57]
  wire [3:0] _atomics_T_13_size; // @[Mux.scala 80:57]
  wire  _atomics_T_13_source; // @[Mux.scala 80:57]
  wire [31:0] _atomics_T_13_address; // @[Mux.scala 80:57]
  wire [7:0] _atomics_T_13_mask; // @[Mux.scala 80:57]
  wire [63:0] _atomics_T_13_data; // @[Mux.scala 80:57]
  wire  _atomics_T_14; // @[Mux.scala 80:60]
  wire [2:0] _atomics_T_15_opcode; // @[Mux.scala 80:57]
  wire [2:0] _atomics_T_15_param; // @[Mux.scala 80:57]
  wire [3:0] _atomics_T_15_size; // @[Mux.scala 80:57]
  wire  _atomics_T_15_source; // @[Mux.scala 80:57]
  wire [31:0] _atomics_T_15_address; // @[Mux.scala 80:57]
  wire [7:0] _atomics_T_15_mask; // @[Mux.scala 80:57]
  wire [63:0] _atomics_T_15_data; // @[Mux.scala 80:57]
  wire  _atomics_T_16; // @[Mux.scala 80:60]
  wire [2:0] atomics_opcode; // @[Mux.scala 80:57]
  wire [2:0] atomics_param; // @[Mux.scala 80:57]
  wire [3:0] atomics_size; // @[Mux.scala 80:57]
  wire  atomics_source; // @[Mux.scala 80:57]
  wire [31:0] atomics_address; // @[Mux.scala 80:57]
  wire [7:0] atomics_mask; // @[Mux.scala 80:57]
  wire [63:0] atomics_data; // @[Mux.scala 80:57]
  wire [39:0] _GEN_356; // @[DCache.scala 577:43]
  wire [39:0] _tl_out_a_valid_T_1; // @[DCache.scala 577:43]
  wire  _tl_out_a_valid_T_3; // @[DCache.scala 577:118]
  wire  _tl_out_a_valid_T_4; // @[DCache.scala 577:27]
  wire  _tl_out_a_valid_T_6; // @[DCache.scala 576:29]
  wire  _tl_out_a_valid_T_12; // @[DCache.scala 577:125]
  wire  tl_out_a_valid; // @[DCache.scala 575:32]
  wire [2:0] _tl_out_a_bits_T_6_opcode; // @[DCache.scala 582:8]
  wire [2:0] _tl_out_a_bits_T_6_param; // @[DCache.scala 582:8]
  wire [3:0] _tl_out_a_bits_T_6_size; // @[DCache.scala 582:8]
  wire  _tl_out_a_bits_T_6_source; // @[DCache.scala 582:8]
  wire [31:0] _tl_out_a_bits_T_6_address; // @[DCache.scala 582:8]
  wire [7:0] _tl_out_a_bits_T_6_mask; // @[DCache.scala 582:8]
  wire [63:0] _tl_out_a_bits_T_6_data; // @[DCache.scala 582:8]
  wire [2:0] _tl_out_a_bits_T_7_opcode; // @[DCache.scala 581:8]
  wire [2:0] _tl_out_a_bits_T_7_param; // @[DCache.scala 581:8]
  wire [3:0] _tl_out_a_bits_T_7_size; // @[DCache.scala 581:8]
  wire  _tl_out_a_bits_T_7_source; // @[DCache.scala 581:8]
  wire [31:0] _tl_out_a_bits_T_7_address; // @[DCache.scala 581:8]
  wire [7:0] putpartial_mask; // @[Edges.scala 483:17 Edges.scala 489:15]
  wire [7:0] _tl_out_a_bits_T_7_mask; // @[DCache.scala 581:8]
  wire [63:0] _tl_out_a_bits_T_7_data; // @[DCache.scala 581:8]
  wire [2:0] _tl_out_a_bits_T_8_opcode; // @[DCache.scala 580:8]
  wire [2:0] _tl_out_a_bits_T_8_param; // @[DCache.scala 580:8]
  wire [3:0] _tl_out_a_bits_T_8_size; // @[DCache.scala 580:8]
  wire  _tl_out_a_bits_T_8_source; // @[DCache.scala 580:8]
  wire [31:0] _tl_out_a_bits_T_8_address; // @[DCache.scala 580:8]
  wire [7:0] _tl_out_a_bits_T_8_mask; // @[DCache.scala 580:8]
  wire [63:0] _tl_out_a_bits_T_8_data; // @[DCache.scala 580:8]
  wire [2:0] tl_out_a_bits_a_param; // @[Edges.scala 345:17 Edges.scala 347:15]
  wire [31:0] tl_out_a_bits_a_address; // @[Edges.scala 345:17 Edges.scala 350:15]
  wire [1:0] _a_sel_T; // @[OneHot.scala 65:12]
  wire  a_sel; // @[DCache.scala 601:66]
  wire  _T_263; // @[Decoupled.scala 40:37]
  wire  _GEN_142; // @[DCache.scala 605:18]
  wire [26:0] _beats1_decode_T_1; // @[package.scala 234:77]
  wire [8:0] beats1_decode; // @[Edges.scala 219:59]
  wire  beats1_opdata; // @[Edges.scala 105:36]
  wire [8:0] beats1; // @[Edges.scala 220:14]
  wire [8:0] counter1; // @[Edges.scala 229:28]
  wire  _last_T; // @[Edges.scala 231:25]
  wire  _last_T_1; // @[Edges.scala 231:47]
  wire  d_last; // @[Edges.scala 231:37]
  wire  d_done; // @[Edges.scala 232:22]
  wire [8:0] count; // @[Edges.scala 233:25]
  wire [11:0] d_address_inc; // @[Edges.scala 268:29]
  wire  grantIsVoluntary; // @[DCache.scala 636:32]
  wire [2:0] _blockProbeAfterGrantCount_T_1; // @[DCache.scala 640:97]
  wire [1:0] _uncachedRespIdxOH_T; // @[OneHot.scala 65:12]
  wire  uncachedRespIdxOH; // @[DCache.scala 643:90]
  wire  _T_273; // @[DCache.scala 648:13]
  wire  _T_276; // @[DCache.scala 657:17]
  wire  _T_278; // @[DCache.scala 658:17]
  wire [31:0] dontCareBits; // @[DCache.scala 672:55]
  wire [31:0] _GEN_357; // @[DCache.scala 673:26]
  wire [31:0] _s2_req_addr_T_1; // @[DCache.scala 673:26]
  wire  _T_281; // @[DCache.scala 679:13]
  wire  _GEN_196; // @[DCache.scala 678:36]
  wire  _GEN_205; // @[DCache.scala 655:35]
  wire  _GEN_209; // @[DCache.scala 646:26]
  wire  _GEN_218; // @[DCache.scala 646:26]
  wire  _GEN_231; // @[DCache.scala 645:26]
  wire  _bundleOut_0_e_valid_T; // @[DCache.scala 685:36]
  wire  _bundleOut_0_e_valid_T_1; // @[DCache.scala 685:47]
  wire  _bundleOut_0_e_valid_T_2; // @[DCache.scala 685:64]
  wire  tl_out__e_valid; // @[DCache.scala 693:51]
  wire  _T_283; // @[Decoupled.scala 40:37]
  wire  _T_285; // @[DCache.scala 687:47]
  wire  _T_286; // @[DCache.scala 687:58]
  wire  _T_287; // @[DCache.scala 687:26]
  wire  _T_289; // @[DCache.scala 687:9]
  wire  _dataArb_io_in_1_valid_T; // @[DCache.scala 692:44]
  wire  _dataArb_io_in_1_valid_T_1; // @[DCache.scala 692:61]
  wire [39:0] _dataArb_io_in_1_bits_addr_T_1; // @[DCache.scala 699:57]
  wire [39:0] _GEN_358; // @[DCache.scala 699:67]
  wire [39:0] _dataArb_io_in_1_bits_addr_T_2; // @[DCache.scala 699:67]
  wire  _metaArb_io_in_3_valid_T; // @[DCache.scala 712:43]
  wire [3:0] _metaArb_io_in_3_bits_data_T_1; // @[Cat.scala 30:58]
  wire  _metaArb_io_in_3_bits_data_T_6; // @[Mux.scala 80:60]
  wire [1:0] _metaArb_io_in_3_bits_data_T_7; // @[Mux.scala 80:57]
  wire  _metaArb_io_in_3_bits_data_T_8; // @[Mux.scala 80:60]
  wire [1:0] _metaArb_io_in_3_bits_data_T_9; // @[Mux.scala 80:57]
  wire  _metaArb_io_in_3_bits_data_T_10; // @[Mux.scala 80:60]
  wire [1:0] _metaArb_io_in_3_bits_data_T_11; // @[Mux.scala 80:57]
  wire  _metaArb_io_in_3_bits_data_T_12; // @[Mux.scala 80:60]
  wire [1:0] metaArb_io_in_3_bits_data_meta_state; // @[Mux.scala 80:57]
  wire  _GEN_234; // @[DCache.scala 726:29]
  wire  _GEN_235; // @[DCache.scala 726:29]
  wire  _GEN_236; // @[DCache.scala 726:29]
  wire  _metaArb_io_in_6_valid_T_1; // @[DCache.scala 740:79]
  wire  _metaArb_io_in_6_valid_T_2; // @[DCache.scala 740:44]
  wire [7:0] metaArb_io_in_6_bits_addr_hi; // @[DCache.scala 744:58]
  wire [39:0] _metaArb_io_in_6_bits_addr_T; // @[Cat.scala 30:58]
  wire [8:0] counter1_1; // @[Edges.scala 229:28]
  wire [8:0] c_count; // @[Edges.scala 233:25]
  reg  s1_release_data_valid; // @[DCache.scala 772:34]
  reg [31:0] _RAND_97;
  wire  releaseRejected; // @[DCache.scala 774:44]
  wire [9:0] _releaseDataBeat_T; // @[Cat.scala 30:58]
  wire [1:0] _releaseDataBeat_T_1; // @[Cat.scala 30:58]
  wire [1:0] _GEN_359; // @[DCache.scala 775:101]
  wire [1:0] _releaseDataBeat_T_3; // @[DCache.scala 775:101]
  wire [1:0] _releaseDataBeat_T_4; // @[DCache.scala 775:52]
  wire [9:0] _GEN_360; // @[DCache.scala 775:47]
  wire [9:0] releaseDataBeat; // @[DCache.scala 775:47]
  wire  _T_298; // @[DCache.scala 788:34]
  wire  _T_299; // @[DCache.scala 788:52]
  wire  _T_301; // @[DCache.scala 788:13]
  wire  discard_line; // @[DCache.scala 789:46]
  wire  _release_state_T_1; // @[DCache.scala 790:44]
  wire [3:0] _release_state_T_13; // @[DCache.scala 790:27]
  wire [5:0] probe_bits_lo; // @[DCache.scala 793:76]
  wire [25:0] _probe_bits_T_1; // @[Cat.scala 30:58]
  wire [31:0] res_2_address; // @[DCache.scala 793:96]
  wire [3:0] _GEN_244; // @[DCache.scala 787:25]
  wire [3:0] _release_state_T_14; // @[DCache.scala 804:29]
  wire [3:0] _release_state_T_15; // @[DCache.scala 808:29]
  wire [2:0] _GEN_255; // @[DCache.scala 801:45]
  wire [3:0] _GEN_261; // @[DCache.scala 801:45]
  wire [3:0] _GEN_263; // @[DCache.scala 799:36]
  wire [2:0] _GEN_266; // @[DCache.scala 799:36]
  wire [3:0] _GEN_273; // @[DCache.scala 797:28]
  wire [2:0] _GEN_276; // @[DCache.scala 797:28]
  wire [3:0] _GEN_284; // @[DCache.scala 795:21]
  wire [2:0] _GEN_287; // @[DCache.scala 795:21]
  wire  _T_304; // @[DCache.scala 812:25]
  wire [39:0] _metaArb_io_in_6_bits_addr_T_1; // @[Cat.scala 30:58]
  wire [3:0] _GEN_294; // @[DCache.scala 816:37]
  wire  _GEN_295; // @[DCache.scala 816:37]
  wire [3:0] _GEN_299; // @[DCache.scala 812:44]
  wire [3:0] _GEN_301; // @[DCache.scala 823:26]
  wire [3:0] _GEN_303; // @[DCache.scala 821:47]
  wire [2:0] _GEN_307; // @[DCache.scala 825:48]
  wire [2:0] _GEN_316; // @[DCache.scala 830:48]
  wire  _T_315; // @[DCache.scala 850:29]
  wire  _GEN_331; // @[DCache.scala 850:41]
  wire [1:0] newCoh_state; // @[DCache.scala 834:102]
  wire  _dataArb_io_in_2_valid_T; // @[DCache.scala 871:60]
  wire [11:0] _dataArb_io_in_2_bits_addr_T_1; // @[DCache.scala 874:55]
  wire [5:0] _dataArb_io_in_2_bits_addr_T_3; // @[DCache.scala 874:117]
  wire [11:0] _GEN_363; // @[DCache.scala 874:72]
  wire  _metaArb_io_in_4_valid_T_1; // @[package.scala 15:47]
  wire [11:0] metaArb_io_in_4_bits_addr_lo; // @[DCache.scala 883:90]
  wire [19:0] metaArb_io_in_4_bits_data_meta_tag; // @[DCache.scala 884:78]
  wire  _T_316; // @[Decoupled.scala 40:37]
  wire  _io_cpu_ordered_T_4; // @[DCache.scala 898:57]
  wire  _io_cpu_ordered_T_5; // @[DCache.scala 898:94]
  wire  _io_cpu_ordered_T_7; // @[DCache.scala 898:115]
  wire  _s1_xcpt_valid_T_1; // @[DCache.scala 900:40]
  reg  io_cpu_s2_xcpt_REG; // @[DCache.scala 901:32]
  reg [31:0] _RAND_98;
  reg  doUncachedResp; // @[DCache.scala 916:27]
  reg [31:0] _RAND_99;
  wire  _T_321; // @[DCache.scala 920:11]
  wire [31:0] io_cpu_resp_bits_data_shifted; // @[AMOALU.scala 39:24]
  wire  _io_cpu_resp_bits_data_T; // @[AMOALU.scala 42:26]
  wire  _io_cpu_resp_bits_data_T_3; // @[AMOALU.scala 42:76]
  wire [31:0] _io_cpu_resp_bits_data_T_5; // @[Bitwise.scala 72:12]
  wire [31:0] io_cpu_resp_bits_data_hi; // @[AMOALU.scala 42:20]
  wire [63:0] _io_cpu_resp_bits_data_T_7; // @[Cat.scala 30:58]
  wire [15:0] io_cpu_resp_bits_data_shifted_1; // @[AMOALU.scala 39:24]
  wire  _io_cpu_resp_bits_data_T_8; // @[AMOALU.scala 42:26]
  wire  _io_cpu_resp_bits_data_T_11; // @[AMOALU.scala 42:76]
  wire [47:0] _io_cpu_resp_bits_data_T_13; // @[Bitwise.scala 72:12]
  wire [47:0] io_cpu_resp_bits_data_hi_1; // @[AMOALU.scala 42:20]
  wire [63:0] _io_cpu_resp_bits_data_T_15; // @[Cat.scala 30:58]
  wire [7:0] io_cpu_resp_bits_data_shifted_2; // @[AMOALU.scala 39:24]
  wire [7:0] io_cpu_resp_bits_data_lo_2; // @[AMOALU.scala 41:23]
  wire  _io_cpu_resp_bits_data_T_16; // @[AMOALU.scala 42:26]
  wire  _io_cpu_resp_bits_data_T_17; // @[AMOALU.scala 42:38]
  wire  _io_cpu_resp_bits_data_T_19; // @[AMOALU.scala 42:76]
  wire [55:0] _io_cpu_resp_bits_data_T_21; // @[Bitwise.scala 72:12]
  wire [55:0] io_cpu_resp_bits_data_hi_2; // @[AMOALU.scala 42:20]
  wire [63:0] _io_cpu_resp_bits_data_T_23; // @[Cat.scala 30:58]
  wire [63:0] _GEN_364; // @[DCache.scala 942:41]
  reg  REG; // @[DCache.scala 976:18]
  reg [31:0] _RAND_100;
  wire  _GEN_349; // @[DCache.scala 976:27]
  wire [8:0] flushCounterNext; // @[DCache.scala 977:39]
  wire  flushDone; // @[DCache.scala 978:57]
  wire  _s1_flush_valid_T; // @[Decoupled.scala 40:37]
  wire  _s1_flush_valid_T_2; // @[DCache.scala 982:45]
  wire  _s1_flush_valid_T_4; // @[DCache.scala 982:64]
  wire  _s1_flush_valid_T_6; // @[DCache.scala 982:95]
  wire [11:0] metaArb_io_in_5_bits_addr_lo; // @[DCache.scala 986:98]
  wire [8:0] _GEN_351; // @[DCache.scala 1019:20]
  reg [8:0] io_cpu_perf_release_counter; // @[Edges.scala 228:27]
  reg [31:0] _RAND_101;
  wire [8:0] io_cpu_perf_release_counter1; // @[Edges.scala 229:28]
  wire  io_cpu_perf_release_first; // @[Edges.scala 230:25]
  wire  _io_cpu_perf_release_last_T; // @[Edges.scala 231:25]
  wire  io_cpu_perf_release_last; // @[Edges.scala 231:37]
  wire  _GEN_367; // @[DCache.scala 648:13]
  wire  _GEN_370; // @[DCache.scala 658:17]
  wire  _GEN_371; // @[DCache.scala 658:17]
  wire  _GEN_372; // @[DCache.scala 658:17]
  wire  _GEN_380; // @[DCache.scala 679:13]
  wire  _GEN_381; // @[DCache.scala 679:13]
  reg [19:0] DCache_state; // @[Register tracking DCache state]
  reg [31:0] _RAND_102;
  reg  DCache_cov [0:1048575]; // @[Coverage map for DCache]
  reg [31:0] _RAND_103;
  wire  DCache_cov_read_data; // @[Coverage map for DCache]
  wire [19:0] DCache_cov_read_addr; // @[Coverage map for DCache]
  wire  DCache_cov_write_data; // @[Coverage map for DCache]
  wire [19:0] DCache_cov_write_addr; // @[Coverage map for DCache]
  wire  DCache_cov_write_mask; // @[Coverage map for DCache]
  wire  DCache_cov_write_en; // @[Coverage map for DCache]
  reg [29:0] DCache_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_104;
  wire  mux_cond_0;
  wire  mux_cond_1;
  wire  mux_cond_2;
  wire  mux_cond_3;
  wire  mux_cond_4;
  wire  mux_cond_5;
  wire [4:0] s2_req_size_shl;
  wire [19:0] s2_req_size_pad;
  wire [9:0] pstore1_held_shl;
  wire [19:0] pstore1_held_pad;
  wire [5:0] s2_req_signed_shl;
  wire [19:0] s2_req_signed_pad;
  wire [10:0] pstore2_valid_shl;
  wire [19:0] pstore2_valid_pad;
  wire [17:0] s1_flush_valid_shl;
  wire [19:0] s1_flush_valid_pad;
  wire [8:0] uncachedInFlight_0_shl;
  wire [19:0] uncachedInFlight_0_pad;
  wire [18:0] blockUncachedGrant_shl;
  wire [19:0] blockUncachedGrant_pad;
  wire [13:0] probe_bits_param_shl;
  wire [19:0] probe_bits_param_pad;
  wire [16:0] s2_flush_valid_pre_tag_ecc_shl;
  wire [19:0] s2_flush_valid_pre_tag_ecc_pad;
  wire [10:0] s1_read_mask_shl;
  wire [19:0] s1_read_mask_pad;
  wire [13:0] s2_victim_way_r_shl;
  wire [19:0] s2_victim_way_r_pad;
  wire [13:0] s1_probe_shl;
  wire [19:0] s1_probe_pad;
  wire [2:0] release_ack_wait_shl;
  wire [19:0] release_ack_wait_pad;
  wire [12:0] s2_hit_state_state_shl;
  wire [19:0] s2_hit_state_state_pad;
  wire [15:0] cached_grant_wait_shl;
  wire [19:0] cached_grant_wait_pad;
  wire [19:0] s1_valid_shl;
  wire [19:0] s1_valid_pad;
  wire [18:0] s2_pma_cacheable_shl;
  wire [19:0] s2_pma_cacheable_pad;
  wire [17:0] s1_did_read_shl;
  wire [19:0] s1_did_read_pad;
  wire [19:0] s2_probe_shl;
  wire [19:0] s2_probe_pad;
  wire [6:0] s2_hit_way_shl;
  wire [19:0] s2_hit_way_pad;
  wire [9:0] s2_not_nacked_in_s1_shl;
  wire [19:0] s2_not_nacked_in_s1_pad;
  wire [18:0] s2_probe_state_state_shl;
  wire [19:0] s2_probe_state_state_pad;
  wire [4:0] s1_req_size_shl;
  wire [19:0] s1_req_size_pad;
  wire [14:0] pstore1_rmw_r_shl;
  wire [19:0] pstore1_rmw_r_pad;
  wire [7:0] s2_release_data_valid_shl;
  wire [19:0] s2_release_data_valid_pad;
  wire [8:0] s2_valid_shl;
  wire [19:0] s2_valid_pad;
  wire [19:0] pstore_drain_on_miss_REG_shl;
  wire [19:0] pstore_drain_on_miss_REG_pad;
  wire [15:0] resetting_shl;
  wire [19:0] resetting_pad;
  wire [19:0] grantInProgress_shl;
  wire [19:0] grantInProgress_pad;
  wire [12:0] s2_probe_way_shl;
  wire [19:0] s2_probe_way_pad;
  wire [11:0] mux_cond_0_shl;
  wire [19:0] mux_cond_0_pad;
  wire [1:0] mux_cond_1_shl;
  wire [19:0] mux_cond_1_pad;
  wire [15:0] mux_cond_2_shl;
  wire [19:0] mux_cond_2_pad;
  wire [6:0] mux_cond_3_shl;
  wire [19:0] mux_cond_3_pad;
  wire [7:0] mux_cond_4_shl;
  wire [19:0] mux_cond_4_pad;
  wire [7:0] mux_cond_5_shl;
  wire [19:0] mux_cond_5_pad;
  wire [19:0] DCache_xor15;
  wire [19:0] DCache_xor16;
  wire [19:0] DCache_xor7;
  wire [19:0] DCache_xor17;
  wire [19:0] DCache_xor38;
  wire [19:0] DCache_xor18;
  wire [19:0] DCache_xor8;
  wire [19:0] DCache_xor3;
  wire [19:0] DCache_xor19;
  wire [19:0] DCache_xor20;
  wire [19:0] DCache_xor9;
  wire [19:0] DCache_xor21;
  wire [19:0] DCache_xor46;
  wire [19:0] DCache_xor22;
  wire [19:0] DCache_xor10;
  wire [19:0] DCache_xor4;
  wire [19:0] DCache_xor1;
  wire [19:0] DCache_xor23;
  wire [19:0] DCache_xor24;
  wire [19:0] DCache_xor11;
  wire [19:0] DCache_xor25;
  wire [19:0] DCache_xor54;
  wire [19:0] DCache_xor26;
  wire [19:0] DCache_xor12;
  wire [19:0] DCache_xor5;
  wire [19:0] DCache_xor27;
  wire [19:0] DCache_xor28;
  wire [19:0] DCache_xor13;
  wire [19:0] DCache_xor29;
  wire [19:0] DCache_xor62;
  wire [19:0] DCache_xor30;
  wire [19:0] DCache_xor14;
  wire [19:0] DCache_xor6;
  wire [19:0] DCache_xor2;
  wire [19:0] DCache_xor0;
  wire [29:0] data_sum;
  wire [29:0] tlb_sum;
  wire [29:0] pma_checker_sum;
  wire [29:0] metaArb_sum;
  wire [29:0] lfsr_prng_sum;
  wire [29:0] amoalu_sum;
  wire [29:0] dataArb_sum;
  wire  stopEn0;
  wire  stopEn1;
  wire  stopEn2;
  wire  stopEn3;
  wire  stopEn4;
  wire  stopEn5;
  wire  stopEn6;
  wire  stopEn7;
  wire  stopEn8;
  wire  stopEn9;
  wire  dataArb_metaAssert_wire;
  wire  metaArb_metaAssert_wire;
  wire  lfsr_prng_metaAssert_wire;
  wire  tlb_metaAssert_wire;
  wire  pma_checker_metaAssert_wire;
  wire  data_metaAssert_wire;
  wire  amoalu_metaAssert_wire;
  wire  DCache_or7;
  wire  DCache_or8;
  wire  DCache_or3;
  wire  DCache_or9;
  wire  DCache_or10;
  wire  DCache_or4;
  wire  DCache_or1;
  wire  DCache_or11;
  wire  DCache_or12;
  wire  DCache_or5;
  wire  DCache_or13;
  wire  DCache_or30;
  wire  DCache_or14;
  wire  DCache_or6;
  wire  DCache_or2;
  wire  DCache_or0;
  TLB tlb ( // @[DCache.scala 117:19]
    .clock(tlb_clock),
    .reset(tlb_reset),
    .io_req_ready(tlb_io_req_ready),
    .io_req_valid(tlb_io_req_valid),
    .io_req_bits_vaddr(tlb_io_req_bits_vaddr),
    .io_req_bits_passthrough(tlb_io_req_bits_passthrough),
    .io_req_bits_size(tlb_io_req_bits_size),
    .io_req_bits_cmd(tlb_io_req_bits_cmd),
    .io_resp_miss(tlb_io_resp_miss),
    .io_resp_paddr(tlb_io_resp_paddr),
    .io_resp_pf_ld(tlb_io_resp_pf_ld),
    .io_resp_pf_st(tlb_io_resp_pf_st),
    .io_resp_ae_ld(tlb_io_resp_ae_ld),
    .io_resp_ae_st(tlb_io_resp_ae_st),
    .io_resp_ma_ld(tlb_io_resp_ma_ld),
    .io_resp_ma_st(tlb_io_resp_ma_st),
    .io_resp_cacheable(tlb_io_resp_cacheable),
    .io_sfence_valid(tlb_io_sfence_valid),
    .io_sfence_bits_rs1(tlb_io_sfence_bits_rs1),
    .io_sfence_bits_rs2(tlb_io_sfence_bits_rs2),
    .io_sfence_bits_addr(tlb_io_sfence_bits_addr),
    .io_ptw_req_ready(tlb_io_ptw_req_ready),
    .io_ptw_req_valid(tlb_io_ptw_req_valid),
    .io_ptw_req_bits_bits_addr(tlb_io_ptw_req_bits_bits_addr),
    .io_ptw_resp_valid(tlb_io_ptw_resp_valid),
    .io_ptw_resp_bits_ae(tlb_io_ptw_resp_bits_ae),
    .io_ptw_resp_bits_pte_ppn(tlb_io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_d(tlb_io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_a(tlb_io_ptw_resp_bits_pte_a),
    .io_ptw_resp_bits_pte_g(tlb_io_ptw_resp_bits_pte_g),
    .io_ptw_resp_bits_pte_u(tlb_io_ptw_resp_bits_pte_u),
    .io_ptw_resp_bits_pte_x(tlb_io_ptw_resp_bits_pte_x),
    .io_ptw_resp_bits_pte_w(tlb_io_ptw_resp_bits_pte_w),
    .io_ptw_resp_bits_pte_r(tlb_io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_v(tlb_io_ptw_resp_bits_pte_v),
    .io_ptw_resp_bits_level(tlb_io_ptw_resp_bits_level),
    .io_ptw_resp_bits_homogeneous(tlb_io_ptw_resp_bits_homogeneous),
    .io_ptw_ptbr_mode(tlb_io_ptw_ptbr_mode),
    .io_ptw_status_debug(tlb_io_ptw_status_debug),
    .io_ptw_status_dprv(tlb_io_ptw_status_dprv),
    .io_ptw_status_mxr(tlb_io_ptw_status_mxr),
    .io_ptw_status_sum(tlb_io_ptw_status_sum),
    .io_ptw_pmp_0_cfg_l(tlb_io_ptw_pmp_0_cfg_l),
    .io_ptw_pmp_0_cfg_a(tlb_io_ptw_pmp_0_cfg_a),
    .io_ptw_pmp_0_cfg_x(tlb_io_ptw_pmp_0_cfg_x),
    .io_ptw_pmp_0_cfg_w(tlb_io_ptw_pmp_0_cfg_w),
    .io_ptw_pmp_0_cfg_r(tlb_io_ptw_pmp_0_cfg_r),
    .io_ptw_pmp_0_addr(tlb_io_ptw_pmp_0_addr),
    .io_ptw_pmp_0_mask(tlb_io_ptw_pmp_0_mask),
    .io_ptw_pmp_1_cfg_l(tlb_io_ptw_pmp_1_cfg_l),
    .io_ptw_pmp_1_cfg_a(tlb_io_ptw_pmp_1_cfg_a),
    .io_ptw_pmp_1_cfg_x(tlb_io_ptw_pmp_1_cfg_x),
    .io_ptw_pmp_1_cfg_w(tlb_io_ptw_pmp_1_cfg_w),
    .io_ptw_pmp_1_cfg_r(tlb_io_ptw_pmp_1_cfg_r),
    .io_ptw_pmp_1_addr(tlb_io_ptw_pmp_1_addr),
    .io_ptw_pmp_1_mask(tlb_io_ptw_pmp_1_mask),
    .io_ptw_pmp_2_cfg_l(tlb_io_ptw_pmp_2_cfg_l),
    .io_ptw_pmp_2_cfg_a(tlb_io_ptw_pmp_2_cfg_a),
    .io_ptw_pmp_2_cfg_x(tlb_io_ptw_pmp_2_cfg_x),
    .io_ptw_pmp_2_cfg_w(tlb_io_ptw_pmp_2_cfg_w),
    .io_ptw_pmp_2_cfg_r(tlb_io_ptw_pmp_2_cfg_r),
    .io_ptw_pmp_2_addr(tlb_io_ptw_pmp_2_addr),
    .io_ptw_pmp_2_mask(tlb_io_ptw_pmp_2_mask),
    .io_ptw_pmp_3_cfg_l(tlb_io_ptw_pmp_3_cfg_l),
    .io_ptw_pmp_3_cfg_a(tlb_io_ptw_pmp_3_cfg_a),
    .io_ptw_pmp_3_cfg_x(tlb_io_ptw_pmp_3_cfg_x),
    .io_ptw_pmp_3_cfg_w(tlb_io_ptw_pmp_3_cfg_w),
    .io_ptw_pmp_3_cfg_r(tlb_io_ptw_pmp_3_cfg_r),
    .io_ptw_pmp_3_addr(tlb_io_ptw_pmp_3_addr),
    .io_ptw_pmp_3_mask(tlb_io_ptw_pmp_3_mask),
    .io_ptw_pmp_4_cfg_l(tlb_io_ptw_pmp_4_cfg_l),
    .io_ptw_pmp_4_cfg_a(tlb_io_ptw_pmp_4_cfg_a),
    .io_ptw_pmp_4_cfg_x(tlb_io_ptw_pmp_4_cfg_x),
    .io_ptw_pmp_4_cfg_w(tlb_io_ptw_pmp_4_cfg_w),
    .io_ptw_pmp_4_cfg_r(tlb_io_ptw_pmp_4_cfg_r),
    .io_ptw_pmp_4_addr(tlb_io_ptw_pmp_4_addr),
    .io_ptw_pmp_4_mask(tlb_io_ptw_pmp_4_mask),
    .io_ptw_pmp_5_cfg_l(tlb_io_ptw_pmp_5_cfg_l),
    .io_ptw_pmp_5_cfg_a(tlb_io_ptw_pmp_5_cfg_a),
    .io_ptw_pmp_5_cfg_x(tlb_io_ptw_pmp_5_cfg_x),
    .io_ptw_pmp_5_cfg_w(tlb_io_ptw_pmp_5_cfg_w),
    .io_ptw_pmp_5_cfg_r(tlb_io_ptw_pmp_5_cfg_r),
    .io_ptw_pmp_5_addr(tlb_io_ptw_pmp_5_addr),
    .io_ptw_pmp_5_mask(tlb_io_ptw_pmp_5_mask),
    .io_ptw_pmp_6_cfg_l(tlb_io_ptw_pmp_6_cfg_l),
    .io_ptw_pmp_6_cfg_a(tlb_io_ptw_pmp_6_cfg_a),
    .io_ptw_pmp_6_cfg_x(tlb_io_ptw_pmp_6_cfg_x),
    .io_ptw_pmp_6_cfg_w(tlb_io_ptw_pmp_6_cfg_w),
    .io_ptw_pmp_6_cfg_r(tlb_io_ptw_pmp_6_cfg_r),
    .io_ptw_pmp_6_addr(tlb_io_ptw_pmp_6_addr),
    .io_ptw_pmp_6_mask(tlb_io_ptw_pmp_6_mask),
    .io_ptw_pmp_7_cfg_l(tlb_io_ptw_pmp_7_cfg_l),
    .io_ptw_pmp_7_cfg_a(tlb_io_ptw_pmp_7_cfg_a),
    .io_ptw_pmp_7_cfg_x(tlb_io_ptw_pmp_7_cfg_x),
    .io_ptw_pmp_7_cfg_w(tlb_io_ptw_pmp_7_cfg_w),
    .io_ptw_pmp_7_cfg_r(tlb_io_ptw_pmp_7_cfg_r),
    .io_ptw_pmp_7_addr(tlb_io_ptw_pmp_7_addr),
    .io_ptw_pmp_7_mask(tlb_io_ptw_pmp_7_mask),
    .io_covSum(tlb_io_covSum),
    .metaAssert(tlb_metaAssert),
    .metaReset(tlb_metaReset)
  );
  TLB pma_checker ( // @[DCache.scala 118:27]
    .clock(pma_checker_clock),
    .reset(pma_checker_reset),
    .io_req_ready(pma_checker_io_req_ready),
    .io_req_valid(pma_checker_io_req_valid),
    .io_req_bits_vaddr(pma_checker_io_req_bits_vaddr),
    .io_req_bits_passthrough(pma_checker_io_req_bits_passthrough),
    .io_req_bits_size(pma_checker_io_req_bits_size),
    .io_req_bits_cmd(pma_checker_io_req_bits_cmd),
    .io_resp_miss(pma_checker_io_resp_miss),
    .io_resp_paddr(pma_checker_io_resp_paddr),
    .io_resp_pf_ld(pma_checker_io_resp_pf_ld),
    .io_resp_pf_st(pma_checker_io_resp_pf_st),
    .io_resp_ae_ld(pma_checker_io_resp_ae_ld),
    .io_resp_ae_st(pma_checker_io_resp_ae_st),
    .io_resp_ma_ld(pma_checker_io_resp_ma_ld),
    .io_resp_ma_st(pma_checker_io_resp_ma_st),
    .io_resp_cacheable(pma_checker_io_resp_cacheable),
    .io_sfence_valid(pma_checker_io_sfence_valid),
    .io_sfence_bits_rs1(pma_checker_io_sfence_bits_rs1),
    .io_sfence_bits_rs2(pma_checker_io_sfence_bits_rs2),
    .io_sfence_bits_addr(pma_checker_io_sfence_bits_addr),
    .io_ptw_req_ready(pma_checker_io_ptw_req_ready),
    .io_ptw_req_valid(pma_checker_io_ptw_req_valid),
    .io_ptw_req_bits_bits_addr(pma_checker_io_ptw_req_bits_bits_addr),
    .io_ptw_resp_valid(pma_checker_io_ptw_resp_valid),
    .io_ptw_resp_bits_ae(pma_checker_io_ptw_resp_bits_ae),
    .io_ptw_resp_bits_pte_ppn(pma_checker_io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_d(pma_checker_io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_a(pma_checker_io_ptw_resp_bits_pte_a),
    .io_ptw_resp_bits_pte_g(pma_checker_io_ptw_resp_bits_pte_g),
    .io_ptw_resp_bits_pte_u(pma_checker_io_ptw_resp_bits_pte_u),
    .io_ptw_resp_bits_pte_x(pma_checker_io_ptw_resp_bits_pte_x),
    .io_ptw_resp_bits_pte_w(pma_checker_io_ptw_resp_bits_pte_w),
    .io_ptw_resp_bits_pte_r(pma_checker_io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_v(pma_checker_io_ptw_resp_bits_pte_v),
    .io_ptw_resp_bits_level(pma_checker_io_ptw_resp_bits_level),
    .io_ptw_resp_bits_homogeneous(pma_checker_io_ptw_resp_bits_homogeneous),
    .io_ptw_ptbr_mode(pma_checker_io_ptw_ptbr_mode),
    .io_ptw_status_debug(pma_checker_io_ptw_status_debug),
    .io_ptw_status_dprv(pma_checker_io_ptw_status_dprv),
    .io_ptw_status_mxr(pma_checker_io_ptw_status_mxr),
    .io_ptw_status_sum(pma_checker_io_ptw_status_sum),
    .io_ptw_pmp_0_cfg_l(pma_checker_io_ptw_pmp_0_cfg_l),
    .io_ptw_pmp_0_cfg_a(pma_checker_io_ptw_pmp_0_cfg_a),
    .io_ptw_pmp_0_cfg_x(pma_checker_io_ptw_pmp_0_cfg_x),
    .io_ptw_pmp_0_cfg_w(pma_checker_io_ptw_pmp_0_cfg_w),
    .io_ptw_pmp_0_cfg_r(pma_checker_io_ptw_pmp_0_cfg_r),
    .io_ptw_pmp_0_addr(pma_checker_io_ptw_pmp_0_addr),
    .io_ptw_pmp_0_mask(pma_checker_io_ptw_pmp_0_mask),
    .io_ptw_pmp_1_cfg_l(pma_checker_io_ptw_pmp_1_cfg_l),
    .io_ptw_pmp_1_cfg_a(pma_checker_io_ptw_pmp_1_cfg_a),
    .io_ptw_pmp_1_cfg_x(pma_checker_io_ptw_pmp_1_cfg_x),
    .io_ptw_pmp_1_cfg_w(pma_checker_io_ptw_pmp_1_cfg_w),
    .io_ptw_pmp_1_cfg_r(pma_checker_io_ptw_pmp_1_cfg_r),
    .io_ptw_pmp_1_addr(pma_checker_io_ptw_pmp_1_addr),
    .io_ptw_pmp_1_mask(pma_checker_io_ptw_pmp_1_mask),
    .io_ptw_pmp_2_cfg_l(pma_checker_io_ptw_pmp_2_cfg_l),
    .io_ptw_pmp_2_cfg_a(pma_checker_io_ptw_pmp_2_cfg_a),
    .io_ptw_pmp_2_cfg_x(pma_checker_io_ptw_pmp_2_cfg_x),
    .io_ptw_pmp_2_cfg_w(pma_checker_io_ptw_pmp_2_cfg_w),
    .io_ptw_pmp_2_cfg_r(pma_checker_io_ptw_pmp_2_cfg_r),
    .io_ptw_pmp_2_addr(pma_checker_io_ptw_pmp_2_addr),
    .io_ptw_pmp_2_mask(pma_checker_io_ptw_pmp_2_mask),
    .io_ptw_pmp_3_cfg_l(pma_checker_io_ptw_pmp_3_cfg_l),
    .io_ptw_pmp_3_cfg_a(pma_checker_io_ptw_pmp_3_cfg_a),
    .io_ptw_pmp_3_cfg_x(pma_checker_io_ptw_pmp_3_cfg_x),
    .io_ptw_pmp_3_cfg_w(pma_checker_io_ptw_pmp_3_cfg_w),
    .io_ptw_pmp_3_cfg_r(pma_checker_io_ptw_pmp_3_cfg_r),
    .io_ptw_pmp_3_addr(pma_checker_io_ptw_pmp_3_addr),
    .io_ptw_pmp_3_mask(pma_checker_io_ptw_pmp_3_mask),
    .io_ptw_pmp_4_cfg_l(pma_checker_io_ptw_pmp_4_cfg_l),
    .io_ptw_pmp_4_cfg_a(pma_checker_io_ptw_pmp_4_cfg_a),
    .io_ptw_pmp_4_cfg_x(pma_checker_io_ptw_pmp_4_cfg_x),
    .io_ptw_pmp_4_cfg_w(pma_checker_io_ptw_pmp_4_cfg_w),
    .io_ptw_pmp_4_cfg_r(pma_checker_io_ptw_pmp_4_cfg_r),
    .io_ptw_pmp_4_addr(pma_checker_io_ptw_pmp_4_addr),
    .io_ptw_pmp_4_mask(pma_checker_io_ptw_pmp_4_mask),
    .io_ptw_pmp_5_cfg_l(pma_checker_io_ptw_pmp_5_cfg_l),
    .io_ptw_pmp_5_cfg_a(pma_checker_io_ptw_pmp_5_cfg_a),
    .io_ptw_pmp_5_cfg_x(pma_checker_io_ptw_pmp_5_cfg_x),
    .io_ptw_pmp_5_cfg_w(pma_checker_io_ptw_pmp_5_cfg_w),
    .io_ptw_pmp_5_cfg_r(pma_checker_io_ptw_pmp_5_cfg_r),
    .io_ptw_pmp_5_addr(pma_checker_io_ptw_pmp_5_addr),
    .io_ptw_pmp_5_mask(pma_checker_io_ptw_pmp_5_mask),
    .io_ptw_pmp_6_cfg_l(pma_checker_io_ptw_pmp_6_cfg_l),
    .io_ptw_pmp_6_cfg_a(pma_checker_io_ptw_pmp_6_cfg_a),
    .io_ptw_pmp_6_cfg_x(pma_checker_io_ptw_pmp_6_cfg_x),
    .io_ptw_pmp_6_cfg_w(pma_checker_io_ptw_pmp_6_cfg_w),
    .io_ptw_pmp_6_cfg_r(pma_checker_io_ptw_pmp_6_cfg_r),
    .io_ptw_pmp_6_addr(pma_checker_io_ptw_pmp_6_addr),
    .io_ptw_pmp_6_mask(pma_checker_io_ptw_pmp_6_mask),
    .io_ptw_pmp_7_cfg_l(pma_checker_io_ptw_pmp_7_cfg_l),
    .io_ptw_pmp_7_cfg_a(pma_checker_io_ptw_pmp_7_cfg_a),
    .io_ptw_pmp_7_cfg_x(pma_checker_io_ptw_pmp_7_cfg_x),
    .io_ptw_pmp_7_cfg_w(pma_checker_io_ptw_pmp_7_cfg_w),
    .io_ptw_pmp_7_cfg_r(pma_checker_io_ptw_pmp_7_cfg_r),
    .io_ptw_pmp_7_addr(pma_checker_io_ptw_pmp_7_addr),
    .io_ptw_pmp_7_mask(pma_checker_io_ptw_pmp_7_mask),
    .io_covSum(pma_checker_io_covSum),
    .metaAssert(pma_checker_metaAssert),
    .metaReset(pma_checker_metaReset)
  );
  MaxPeriodFibonacciLFSR lfsr_prng ( // @[PRNG.scala 82:22]
    .clock(lfsr_prng_clock),
    .reset(lfsr_prng_reset),
    .io_increment(lfsr_prng_io_increment),
    .io_out_0(lfsr_prng_io_out_0),
    .io_out_1(lfsr_prng_io_out_1),
    .io_out_2(lfsr_prng_io_out_2),
    .io_out_3(lfsr_prng_io_out_3),
    .io_out_4(lfsr_prng_io_out_4),
    .io_out_5(lfsr_prng_io_out_5),
    .io_out_6(lfsr_prng_io_out_6),
    .io_out_7(lfsr_prng_io_out_7),
    .io_out_8(lfsr_prng_io_out_8),
    .io_out_9(lfsr_prng_io_out_9),
    .io_out_10(lfsr_prng_io_out_10),
    .io_out_11(lfsr_prng_io_out_11),
    .io_out_12(lfsr_prng_io_out_12),
    .io_out_13(lfsr_prng_io_out_13),
    .io_out_14(lfsr_prng_io_out_14),
    .io_out_15(lfsr_prng_io_out_15),
    .io_covSum(lfsr_prng_io_covSum),
    .metaAssert(lfsr_prng_metaAssert),
    .metaReset(lfsr_prng_metaReset)
  );
  DCacheModuleImpl_Anon_1 metaArb ( // @[DCache.scala 122:23]
    .io_in_0_valid(metaArb_io_in_0_valid),
    .io_in_0_bits_addr(metaArb_io_in_0_bits_addr),
    .io_in_0_bits_idx(metaArb_io_in_0_bits_idx),
    .io_in_1_valid(metaArb_io_in_1_valid),
    .io_in_1_bits_addr(metaArb_io_in_1_bits_addr),
    .io_in_1_bits_idx(metaArb_io_in_1_bits_idx),
    .io_in_1_bits_data(metaArb_io_in_1_bits_data),
    .io_in_2_valid(metaArb_io_in_2_valid),
    .io_in_2_bits_addr(metaArb_io_in_2_bits_addr),
    .io_in_2_bits_idx(metaArb_io_in_2_bits_idx),
    .io_in_2_bits_way_en(metaArb_io_in_2_bits_way_en),
    .io_in_2_bits_data(metaArb_io_in_2_bits_data),
    .io_in_3_valid(metaArb_io_in_3_valid),
    .io_in_3_bits_addr(metaArb_io_in_3_bits_addr),
    .io_in_3_bits_idx(metaArb_io_in_3_bits_idx),
    .io_in_3_bits_way_en(metaArb_io_in_3_bits_way_en),
    .io_in_3_bits_data(metaArb_io_in_3_bits_data),
    .io_in_4_ready(metaArb_io_in_4_ready),
    .io_in_4_valid(metaArb_io_in_4_valid),
    .io_in_4_bits_addr(metaArb_io_in_4_bits_addr),
    .io_in_4_bits_idx(metaArb_io_in_4_bits_idx),
    .io_in_4_bits_way_en(metaArb_io_in_4_bits_way_en),
    .io_in_4_bits_data(metaArb_io_in_4_bits_data),
    .io_in_5_ready(metaArb_io_in_5_ready),
    .io_in_5_valid(metaArb_io_in_5_valid),
    .io_in_5_bits_addr(metaArb_io_in_5_bits_addr),
    .io_in_5_bits_idx(metaArb_io_in_5_bits_idx),
    .io_in_6_ready(metaArb_io_in_6_ready),
    .io_in_6_valid(metaArb_io_in_6_valid),
    .io_in_6_bits_addr(metaArb_io_in_6_bits_addr),
    .io_in_6_bits_idx(metaArb_io_in_6_bits_idx),
    .io_in_6_bits_way_en(metaArb_io_in_6_bits_way_en),
    .io_in_6_bits_data(metaArb_io_in_6_bits_data),
    .io_in_7_ready(metaArb_io_in_7_ready),
    .io_in_7_valid(metaArb_io_in_7_valid),
    .io_in_7_bits_addr(metaArb_io_in_7_bits_addr),
    .io_in_7_bits_idx(metaArb_io_in_7_bits_idx),
    .io_in_7_bits_way_en(metaArb_io_in_7_bits_way_en),
    .io_in_7_bits_data(metaArb_io_in_7_bits_data),
    .io_out_valid(metaArb_io_out_valid),
    .io_out_bits_write(metaArb_io_out_bits_write),
    .io_out_bits_addr(metaArb_io_out_bits_addr),
    .io_out_bits_idx(metaArb_io_out_bits_idx),
    .io_out_bits_way_en(metaArb_io_out_bits_way_en),
    .io_out_bits_data(metaArb_io_out_bits_data),
    .io_covSum(metaArb_io_covSum),
    .metaAssert(metaArb_metaAssert)
  );
  DCacheDataArray data ( // @[DCache.scala 132:20]
    .clock(data_clock),
    .io_req_valid(data_io_req_valid),
    .io_req_bits_addr(data_io_req_bits_addr),
    .io_req_bits_write(data_io_req_bits_write),
    .io_req_bits_wdata(data_io_req_bits_wdata),
    .io_req_bits_eccMask(data_io_req_bits_eccMask),
    .io_req_bits_way_en(data_io_req_bits_way_en),
    .io_resp_0(data_io_resp_0),
    .io_resp_1(data_io_resp_1),
    .io_resp_2(data_io_resp_2),
    .io_resp_3(data_io_resp_3),
    .io_covSum(data_io_covSum),
    .metaAssert(data_metaAssert),
    .metaReset(data_metaReset)
  );
  DCacheModuleImpl_Anon_2 dataArb ( // @[DCache.scala 133:23]
    .io_in_0_valid(dataArb_io_in_0_valid),
    .io_in_0_bits_addr(dataArb_io_in_0_bits_addr),
    .io_in_0_bits_write(dataArb_io_in_0_bits_write),
    .io_in_0_bits_wdata(dataArb_io_in_0_bits_wdata),
    .io_in_0_bits_eccMask(dataArb_io_in_0_bits_eccMask),
    .io_in_0_bits_way_en(dataArb_io_in_0_bits_way_en),
    .io_in_1_ready(dataArb_io_in_1_ready),
    .io_in_1_valid(dataArb_io_in_1_valid),
    .io_in_1_bits_addr(dataArb_io_in_1_bits_addr),
    .io_in_1_bits_write(dataArb_io_in_1_bits_write),
    .io_in_1_bits_wdata(dataArb_io_in_1_bits_wdata),
    .io_in_1_bits_way_en(dataArb_io_in_1_bits_way_en),
    .io_in_2_ready(dataArb_io_in_2_ready),
    .io_in_2_valid(dataArb_io_in_2_valid),
    .io_in_2_bits_addr(dataArb_io_in_2_bits_addr),
    .io_in_2_bits_wdata(dataArb_io_in_2_bits_wdata),
    .io_in_3_ready(dataArb_io_in_3_ready),
    .io_in_3_valid(dataArb_io_in_3_valid),
    .io_in_3_bits_addr(dataArb_io_in_3_bits_addr),
    .io_in_3_bits_wdata(dataArb_io_in_3_bits_wdata),
    .io_in_3_bits_wordMask(dataArb_io_in_3_bits_wordMask),
    .io_out_valid(dataArb_io_out_valid),
    .io_out_bits_addr(dataArb_io_out_bits_addr),
    .io_out_bits_write(dataArb_io_out_bits_write),
    .io_out_bits_wdata(dataArb_io_out_bits_wdata),
    .io_out_bits_eccMask(dataArb_io_out_bits_eccMask),
    .io_out_bits_way_en(dataArb_io_out_bits_way_en),
    .io_covSum(dataArb_io_covSum),
    .metaAssert(dataArb_metaAssert)
  );
  AMOALU amoalu ( // @[DCache.scala 950:26]
    .io_mask(amoalu_io_mask),
    .io_cmd(amoalu_io_cmd),
    .io_lhs(amoalu_io_lhs),
    .io_rhs(amoalu_io_rhs),
    .io_out(amoalu_io_out),
    .io_covSum(amoalu_io_covSum),
    .metaAssert(amoalu_metaAssert)
  );
  assign tag_array_0_s1_meta_addr = tag_array_0_s1_meta_addr_pipe_0;
  assign tag_array_0_s1_meta_data = tag_array_0[tag_array_0_s1_meta_addr]; // @[DescribedSRAM.scala 19:26]
  assign tag_array_0_MPORT_data = metaArb_io_out_bits_data;
  assign tag_array_0_MPORT_addr = metaArb_io_out_bits_idx;
  assign tag_array_0_MPORT_mask = metaArb_io_out_bits_way_en[0];
  assign tag_array_0_MPORT_en = metaArb_io_out_valid & metaArb_io_out_bits_write;
  assign tag_array_1_s1_meta_addr = tag_array_1_s1_meta_addr_pipe_0;
  assign tag_array_1_s1_meta_data = tag_array_1[tag_array_1_s1_meta_addr]; // @[DescribedSRAM.scala 19:26]
  assign tag_array_1_MPORT_data = metaArb_io_out_bits_data;
  assign tag_array_1_MPORT_addr = metaArb_io_out_bits_idx;
  assign tag_array_1_MPORT_mask = metaArb_io_out_bits_way_en[1];
  assign tag_array_1_MPORT_en = metaArb_io_out_valid & metaArb_io_out_bits_write;
  assign tag_array_2_s1_meta_addr = tag_array_2_s1_meta_addr_pipe_0;
  assign tag_array_2_s1_meta_data = tag_array_2[tag_array_2_s1_meta_addr]; // @[DescribedSRAM.scala 19:26]
  assign tag_array_2_MPORT_data = metaArb_io_out_bits_data;
  assign tag_array_2_MPORT_addr = metaArb_io_out_bits_idx;
  assign tag_array_2_MPORT_mask = metaArb_io_out_bits_way_en[2];
  assign tag_array_2_MPORT_en = metaArb_io_out_valid & metaArb_io_out_bits_write;
  assign tag_array_3_s1_meta_addr = tag_array_3_s1_meta_addr_pipe_0;
  assign tag_array_3_s1_meta_data = tag_array_3[tag_array_3_s1_meta_addr]; // @[DescribedSRAM.scala 19:26]
  assign tag_array_3_MPORT_data = metaArb_io_out_bits_data;
  assign tag_array_3_MPORT_addr = metaArb_io_out_bits_idx;
  assign tag_array_3_MPORT_mask = metaArb_io_out_bits_way_en[3];
  assign tag_array_3_MPORT_en = metaArb_io_out_valid & metaArb_io_out_bits_write;
  assign lfsr_lo = {lfsr_prng_io_out_7,lfsr_prng_io_out_6,lfsr_prng_io_out_5,lfsr_prng_io_out_4,lfsr_prng_io_out_3,lfsr_prng_io_out_2,lfsr_prng_io_out_1,lfsr_prng_io_out_0}; // @[PRNG.scala 86:17]
  assign lfsr = {lfsr_prng_io_out_15,lfsr_prng_io_out_14,lfsr_prng_io_out_13,lfsr_prng_io_out_12,lfsr_prng_io_out_11,lfsr_prng_io_out_10,lfsr_prng_io_out_9,lfsr_prng_io_out_8,lfsr_lo}; // @[PRNG.scala 86:17]
  assign s1_valid_x9 = io_cpu_req_ready & io_cpu_req_valid; // @[Decoupled.scala 40:37]
  assign _block_probe_for_core_progress_T = blockProbeAfterGrantCount > 3'h0; // @[DCache.scala 737:65]
  assign lrscValid = lrscCount > 7'h3; // @[DCache.scala 444:29]
  assign block_probe_for_core_progress = _block_probe_for_core_progress_T | lrscValid; // @[DCache.scala 737:69]
  assign _releaseInFlight_T = s1_probe | s2_probe; // @[DCache.scala 305:34]
  assign _releaseInFlight_T_1 = release_state != 4'h0; // @[DCache.scala 305:63]
  assign releaseInFlight = _releaseInFlight_T | _releaseInFlight_T_1; // @[DCache.scala 305:46]
  assign _block_probe_for_pending_release_ack_T = auto_out_b_bits_address ^ release_ack_addr; // @[DCache.scala 738:88]
  assign _block_probe_for_pending_release_ack_T_2 = _block_probe_for_pending_release_ack_T[20:6] == 15'h0; // @[DCache.scala 738:163]
  assign block_probe_for_pending_release_ack = release_ack_wait & _block_probe_for_pending_release_ack_T_2; // @[DCache.scala 738:62]
  assign _block_probe_for_ordering_T = releaseInFlight | block_probe_for_pending_release_ack; // @[DCache.scala 739:50]
  assign block_probe_for_ordering = _block_probe_for_ordering_T | grantInProgress; // @[DCache.scala 739:89]
  assign _bundleOut_0_b_ready_T = block_probe_for_core_progress | block_probe_for_ordering; // @[DCache.scala 741:79]
  assign _bundleOut_0_b_ready_T_1 = _bundleOut_0_b_ready_T | s1_valid; // @[DCache.scala 741:107]
  assign _bundleOut_0_b_ready_T_2 = _bundleOut_0_b_ready_T_1 | s2_valid; // @[DCache.scala 741:119]
  assign tl_out__b_ready = metaArb_io_in_6_ready & ~_bundleOut_0_b_ready_T_2; // @[DCache.scala 741:44]
  assign s1_probe_x12 = tl_out__b_ready & auto_out_b_valid; // @[Decoupled.scala 40:37]
  assign s1_valid_masked = s1_valid & ~io_cpu_s1_kill; // @[DCache.scala 166:34]
  assign s2_meta_error = |4'h0; // @[DCache.scala 333:83]
  assign _T_118 = {probe_bits_param,s2_probe_state_state}; // @[Cat.scala 30:58]
  assign _T_175 = 4'h3 == _T_118; // @[Misc.scala 55:20]
  assign _T_171 = 4'h2 == _T_118; // @[Misc.scala 55:20]
  assign _T_167 = 4'h1 == _T_118; // @[Misc.scala 55:20]
  assign _T_163 = 4'h0 == _T_118; // @[Misc.scala 55:20]
  assign _T_159 = 4'h7 == _T_118; // @[Misc.scala 55:20]
  assign _T_155 = 4'h6 == _T_118; // @[Misc.scala 55:20]
  assign _T_151 = 4'h5 == _T_118; // @[Misc.scala 55:20]
  assign _T_147 = 4'h4 == _T_118; // @[Misc.scala 55:20]
  assign _T_143 = 4'hb == _T_118; // @[Misc.scala 55:20]
  assign _T_139 = 4'ha == _T_118; // @[Misc.scala 55:20]
  assign _T_135 = 4'h9 == _T_118; // @[Misc.scala 55:20]
  assign _T_131 = 4'h8 == _T_118; // @[Misc.scala 55:20]
  assign _T_148 = _T_147 ? 1'h0 : _T_143; // @[Misc.scala 37:9]
  assign _T_152 = _T_151 ? 1'h0 : _T_148; // @[Misc.scala 37:9]
  assign _T_156 = _T_155 ? 1'h0 : _T_152; // @[Misc.scala 37:9]
  assign _T_160 = _T_159 | _T_156; // @[Misc.scala 37:9]
  assign _T_164 = _T_163 ? 1'h0 : _T_160; // @[Misc.scala 37:9]
  assign _T_168 = _T_167 ? 1'h0 : _T_164; // @[Misc.scala 37:9]
  assign _T_172 = _T_171 ? 1'h0 : _T_168; // @[Misc.scala 37:9]
  assign s2_prb_ack_data = _T_175 | _T_172; // @[Misc.scala 37:9]
  assign _T_303 = s2_probe_state_state > 2'h0; // @[Metadata.scala 49:45]
  assign _last_T_2 = counter_1 == 9'h1; // @[Edges.scala 231:25]
  assign _T_308 = release_state == 4'h1; // @[package.scala 15:47]
  assign _T_309 = release_state == 4'h6; // @[package.scala 15:47]
  assign _T_311 = _T_308 | _T_309; // @[package.scala 72:59]
  assign _T_310 = release_state == 4'h9; // @[package.scala 15:47]
  assign _T_312 = _T_311 | _T_310; // @[package.scala 72:59]
  assign _GEN_323 = _T_310 ? 3'h6 : 3'h7; // @[DCache.scala 835:52]
  assign _T_307 = release_state == 4'h2; // @[DCache.scala 830:25]
  assign _T_306 = release_state == 4'h3; // @[DCache.scala 825:25]
  assign _GEN_315 = _T_307 ? 3'h5 : 3'h4; // @[DCache.scala 830:48]
  assign tl_out__c_bits_opcode = _T_312 ? _GEN_323 : _GEN_315; // @[DCache.scala 834:102]
  assign beats1_opdata_1 = tl_out__c_bits_opcode[0]; // @[Edges.scala 101:36]
  assign tl_out__c_bits_size = _T_312 ? 4'h6 : probe_bits_size; // @[DCache.scala 834:102]
  assign _beats1_decode_T_5 = 27'hfff << tl_out__c_bits_size; // @[package.scala 234:77]
  assign beats1_decode_1 = ~_beats1_decode_T_5[11:3]; // @[Edges.scala 219:59]
  assign beats1_1 = beats1_opdata_1 ? beats1_decode_1 : 9'h0; // @[Edges.scala 220:14]
  assign _last_T_3 = beats1_1 == 9'h0; // @[Edges.scala 231:47]
  assign c_last = _last_T_2 | _last_T_3; // @[Edges.scala 231:37]
  assign _T_305 = release_state == 4'h5; // @[DCache.scala 821:25]
  assign c_first = counter_1 == 9'h0; // @[Edges.scala 230:25]
  assign _bundleOut_0_c_valid_T_3 = c_first & release_ack_wait; // @[DCache.scala 781:128]
  assign _bundleOut_0_c_valid_T_5 = s2_release_data_valid & ~_bundleOut_0_c_valid_T_3; // @[DCache.scala 781:115]
  assign _GEN_264 = s2_prb_ack_data ? _bundleOut_0_c_valid_T_5 : 1'h1; // @[DCache.scala 799:36]
  assign _GEN_274 = s2_meta_error ? _bundleOut_0_c_valid_T_5 : _GEN_264; // @[DCache.scala 797:28]
  assign _GEN_285 = s2_probe ? _GEN_274 : _bundleOut_0_c_valid_T_5; // @[DCache.scala 795:21]
  assign _GEN_302 = _T_305 | _GEN_285; // @[DCache.scala 821:47]
  assign tl_out__c_valid = _T_306 | _GEN_302; // @[DCache.scala 825:48]
  assign _T_297 = auto_out_c_ready & tl_out__c_valid; // @[Decoupled.scala 40:37]
  assign releaseDone = c_last & _T_297; // @[Edges.scala 232:22]
  assign _GEN_262 = _T_303 | ~releaseDone; // @[DCache.scala 801:45]
  assign _GEN_272 = s2_prb_ack_data | _GEN_262; // @[DCache.scala 799:36]
  assign probeNack = s2_meta_error | _GEN_272; // @[DCache.scala 797:28]
  assign _s1_read_T = s1_req_cmd == 5'h0; // @[Consts.scala 81:31]
  assign _s1_read_T_1 = s1_req_cmd == 5'h6; // @[Consts.scala 81:48]
  assign _s1_read_T_2 = _s1_read_T | _s1_read_T_1; // @[Consts.scala 81:41]
  assign _s1_read_T_3 = s1_req_cmd == 5'h7; // @[Consts.scala 81:65]
  assign _s1_read_T_4 = _s1_read_T_2 | _s1_read_T_3; // @[Consts.scala 81:58]
  assign _s1_read_T_5 = s1_req_cmd == 5'h4; // @[package.scala 15:47]
  assign _s1_read_T_6 = s1_req_cmd == 5'h9; // @[package.scala 15:47]
  assign _s1_read_T_9 = _s1_read_T_5 | _s1_read_T_6; // @[package.scala 72:59]
  assign _s1_read_T_7 = s1_req_cmd == 5'ha; // @[package.scala 15:47]
  assign _s1_read_T_10 = _s1_read_T_9 | _s1_read_T_7; // @[package.scala 72:59]
  assign _s1_read_T_8 = s1_req_cmd == 5'hb; // @[package.scala 15:47]
  assign _s1_read_T_11 = _s1_read_T_10 | _s1_read_T_8; // @[package.scala 72:59]
  assign _s1_read_T_12 = s1_req_cmd == 5'h8; // @[package.scala 15:47]
  assign _s1_read_T_13 = s1_req_cmd == 5'hc; // @[package.scala 15:47]
  assign _s1_read_T_17 = _s1_read_T_12 | _s1_read_T_13; // @[package.scala 72:59]
  assign _s1_read_T_14 = s1_req_cmd == 5'hd; // @[package.scala 15:47]
  assign _s1_read_T_18 = _s1_read_T_17 | _s1_read_T_14; // @[package.scala 72:59]
  assign _s1_read_T_15 = s1_req_cmd == 5'he; // @[package.scala 15:47]
  assign _s1_read_T_19 = _s1_read_T_18 | _s1_read_T_15; // @[package.scala 72:59]
  assign _s1_read_T_16 = s1_req_cmd == 5'hf; // @[package.scala 15:47]
  assign _s1_read_T_20 = _s1_read_T_19 | _s1_read_T_16; // @[package.scala 72:59]
  assign _s1_read_T_21 = _s1_read_T_11 | _s1_read_T_20; // @[Consts.scala 79:44]
  assign s1_read = _s1_read_T_4 | _s1_read_T_21; // @[Consts.scala 81:75]
  assign _s2_write_T = s2_req_cmd == 5'h1; // @[Consts.scala 82:32]
  assign _s2_write_T_1 = s2_req_cmd == 5'h11; // @[Consts.scala 82:49]
  assign _s2_write_T_2 = _s2_write_T | _s2_write_T_1; // @[Consts.scala 82:42]
  assign _s2_write_T_3 = s2_req_cmd == 5'h7; // @[Consts.scala 82:66]
  assign _s2_write_T_4 = _s2_write_T_2 | _s2_write_T_3; // @[Consts.scala 82:59]
  assign _s2_write_T_5 = s2_req_cmd == 5'h4; // @[package.scala 15:47]
  assign _s2_write_T_6 = s2_req_cmd == 5'h9; // @[package.scala 15:47]
  assign _s2_write_T_9 = _s2_write_T_5 | _s2_write_T_6; // @[package.scala 72:59]
  assign _s2_write_T_7 = s2_req_cmd == 5'ha; // @[package.scala 15:47]
  assign _s2_write_T_10 = _s2_write_T_9 | _s2_write_T_7; // @[package.scala 72:59]
  assign _s2_write_T_8 = s2_req_cmd == 5'hb; // @[package.scala 15:47]
  assign _s2_write_T_11 = _s2_write_T_10 | _s2_write_T_8; // @[package.scala 72:59]
  assign _s2_write_T_12 = s2_req_cmd == 5'h8; // @[package.scala 15:47]
  assign _s2_write_T_13 = s2_req_cmd == 5'hc; // @[package.scala 15:47]
  assign _s2_write_T_17 = _s2_write_T_12 | _s2_write_T_13; // @[package.scala 72:59]
  assign _s2_write_T_14 = s2_req_cmd == 5'hd; // @[package.scala 15:47]
  assign _s2_write_T_18 = _s2_write_T_17 | _s2_write_T_14; // @[package.scala 72:59]
  assign _s2_write_T_15 = s2_req_cmd == 5'he; // @[package.scala 15:47]
  assign _s2_write_T_19 = _s2_write_T_18 | _s2_write_T_15; // @[package.scala 72:59]
  assign _s2_write_T_16 = s2_req_cmd == 5'hf; // @[package.scala 15:47]
  assign _s2_write_T_20 = _s2_write_T_19 | _s2_write_T_16; // @[package.scala 72:59]
  assign _s2_write_T_21 = _s2_write_T_11 | _s2_write_T_20; // @[Consts.scala 79:44]
  assign s2_write = _s2_write_T_4 | _s2_write_T_21; // @[Consts.scala 82:76]
  assign _pstore1_valid_likely_T = s2_valid & s2_write; // @[DCache.scala 476:39]
  assign pstore1_valid_likely = _pstore1_valid_likely_T | pstore1_held; // @[DCache.scala 476:51]
  assign s1_vaddr_hi = s1_req_addr[39:12]; // @[DCache.scala 177:56]
  assign s1_vaddr_lo = s1_req_addr[11:0]; // @[DCache.scala 177:78]
  assign s1_vaddr = {s1_vaddr_hi,s1_vaddr_lo}; // @[Cat.scala 30:58]
  assign _s1_hazard_T_2 = pstore1_addr[11:3] == s1_vaddr[11:3]; // @[DCache.scala 532:31]
  assign _s1_write_T = s1_req_cmd == 5'h1; // @[Consts.scala 82:32]
  assign _s1_write_T_1 = s1_req_cmd == 5'h11; // @[Consts.scala 82:49]
  assign _s1_write_T_2 = _s1_write_T | _s1_write_T_1; // @[Consts.scala 82:42]
  assign _s1_write_T_4 = _s1_write_T_2 | _s1_read_T_3; // @[Consts.scala 82:59]
  assign s1_write = _s1_write_T_4 | _s1_read_T_21; // @[Consts.scala 82:76]
  assign s1_hazard_hi_hi_hi = |pstore1_mask[7]; // @[DCache.scala 1149:66]
  assign s1_hazard_hi_hi_lo = |pstore1_mask[6]; // @[DCache.scala 1149:66]
  assign s1_hazard_hi_lo_hi = |pstore1_mask[5]; // @[DCache.scala 1149:66]
  assign s1_hazard_hi_lo_lo = |pstore1_mask[4]; // @[DCache.scala 1149:66]
  assign s1_hazard_lo_hi_hi = |pstore1_mask[3]; // @[DCache.scala 1149:66]
  assign s1_hazard_lo_hi_lo = |pstore1_mask[2]; // @[DCache.scala 1149:66]
  assign s1_hazard_lo_lo_hi = |pstore1_mask[1]; // @[DCache.scala 1149:66]
  assign s1_hazard_lo_lo_lo = |pstore1_mask[0]; // @[DCache.scala 1149:66]
  assign _s1_hazard_T_11 = {s1_hazard_hi_hi_hi,s1_hazard_hi_hi_lo,s1_hazard_hi_lo_hi,s1_hazard_hi_lo_lo,s1_hazard_lo_hi_hi,s1_hazard_lo_hi_lo,s1_hazard_lo_lo_hi,s1_hazard_lo_lo_lo}; // @[Cat.scala 30:58]
  assign s1_hazard_hi_hi_hi_1 = _s1_hazard_T_11[7]; // @[Bitwise.scala 26:51]
  assign s1_hazard_hi_hi_lo_1 = _s1_hazard_T_11[6]; // @[Bitwise.scala 26:51]
  assign s1_hazard_hi_lo_hi_1 = _s1_hazard_T_11[5]; // @[Bitwise.scala 26:51]
  assign s1_hazard_hi_lo_lo_1 = _s1_hazard_T_11[4]; // @[Bitwise.scala 26:51]
  assign s1_hazard_lo_hi_hi_1 = _s1_hazard_T_11[3]; // @[Bitwise.scala 26:51]
  assign s1_hazard_lo_hi_lo_1 = _s1_hazard_T_11[2]; // @[Bitwise.scala 26:51]
  assign s1_hazard_lo_lo_hi_1 = _s1_hazard_T_11[1]; // @[Bitwise.scala 26:51]
  assign s1_hazard_lo_lo_lo_1 = _s1_hazard_T_11[0]; // @[Bitwise.scala 26:51]
  assign _s1_hazard_T_12 = {s1_hazard_hi_hi_hi_1,s1_hazard_hi_hi_lo_1,s1_hazard_hi_lo_hi_1,s1_hazard_hi_lo_lo_1,s1_hazard_lo_hi_hi_1,s1_hazard_lo_hi_lo_1,s1_hazard_lo_lo_hi_1,s1_hazard_lo_lo_lo_1}; // @[Cat.scala 30:58]
  assign _s1_mask_xwr_upper_T_2 = s1_req_size >= 2'h1; // @[AMOALU.scala 17:57]
  assign s1_mask_xwr_hi = s1_req_addr[0] | _s1_mask_xwr_upper_T_2; // @[AMOALU.scala 17:46]
  assign s1_mask_xwr_lo = s1_req_addr[0] ? 1'h0 : 1'h1; // @[AMOALU.scala 18:22]
  assign _s1_mask_xwr_T = {s1_mask_xwr_hi,s1_mask_xwr_lo}; // @[Cat.scala 30:58]
  assign _s1_mask_xwr_upper_T_5 = s1_req_addr[1] ? _s1_mask_xwr_T : 2'h0; // @[AMOALU.scala 17:22]
  assign _s1_mask_xwr_upper_T_6 = s1_req_size >= 2'h2; // @[AMOALU.scala 17:57]
  assign _s1_mask_xwr_upper_T_7 = _s1_mask_xwr_upper_T_6 ? 2'h3 : 2'h0; // @[AMOALU.scala 17:51]
  assign s1_mask_xwr_hi_1 = _s1_mask_xwr_upper_T_5 | _s1_mask_xwr_upper_T_7; // @[AMOALU.scala 17:46]
  assign s1_mask_xwr_lo_1 = s1_req_addr[1] ? 2'h0 : _s1_mask_xwr_T; // @[AMOALU.scala 18:22]
  assign _s1_mask_xwr_T_1 = {s1_mask_xwr_hi_1,s1_mask_xwr_lo_1}; // @[Cat.scala 30:58]
  assign _s1_mask_xwr_upper_T_9 = s1_req_addr[2] ? _s1_mask_xwr_T_1 : 4'h0; // @[AMOALU.scala 17:22]
  assign _s1_mask_xwr_upper_T_10 = s1_req_size >= 2'h3; // @[AMOALU.scala 17:57]
  assign _s1_mask_xwr_upper_T_11 = _s1_mask_xwr_upper_T_10 ? 4'hf : 4'h0; // @[AMOALU.scala 17:51]
  assign s1_mask_xwr_hi_2 = _s1_mask_xwr_upper_T_9 | _s1_mask_xwr_upper_T_11; // @[AMOALU.scala 17:46]
  assign s1_mask_xwr_lo_2 = s1_req_addr[2] ? 4'h0 : _s1_mask_xwr_T_1; // @[AMOALU.scala 18:22]
  assign s1_mask_xwr = {s1_mask_xwr_hi_2,s1_mask_xwr_lo_2}; // @[Cat.scala 30:58]
  assign s1_hazard_hi_hi_hi_2 = |s1_mask_xwr[7]; // @[DCache.scala 1149:66]
  assign s1_hazard_hi_hi_lo_2 = |s1_mask_xwr[6]; // @[DCache.scala 1149:66]
  assign s1_hazard_hi_lo_hi_2 = |s1_mask_xwr[5]; // @[DCache.scala 1149:66]
  assign s1_hazard_hi_lo_lo_2 = |s1_mask_xwr[4]; // @[DCache.scala 1149:66]
  assign s1_hazard_lo_hi_hi_2 = |s1_mask_xwr[3]; // @[DCache.scala 1149:66]
  assign s1_hazard_lo_hi_lo_2 = |s1_mask_xwr[2]; // @[DCache.scala 1149:66]
  assign s1_hazard_lo_lo_hi_2 = |s1_mask_xwr[1]; // @[DCache.scala 1149:66]
  assign s1_hazard_lo_lo_lo_2 = |s1_mask_xwr[0]; // @[DCache.scala 1149:66]
  assign _s1_hazard_T_21 = {s1_hazard_hi_hi_hi_2,s1_hazard_hi_hi_lo_2,s1_hazard_hi_lo_hi_2,s1_hazard_hi_lo_lo_2,s1_hazard_lo_hi_hi_2,s1_hazard_lo_hi_lo_2,s1_hazard_lo_lo_hi_2,s1_hazard_lo_lo_lo_2}; // @[Cat.scala 30:58]
  assign s1_hazard_hi_hi_hi_3 = _s1_hazard_T_21[7]; // @[Bitwise.scala 26:51]
  assign s1_hazard_hi_hi_lo_3 = _s1_hazard_T_21[6]; // @[Bitwise.scala 26:51]
  assign s1_hazard_hi_lo_hi_3 = _s1_hazard_T_21[5]; // @[Bitwise.scala 26:51]
  assign s1_hazard_hi_lo_lo_3 = _s1_hazard_T_21[4]; // @[Bitwise.scala 26:51]
  assign s1_hazard_lo_hi_hi_3 = _s1_hazard_T_21[3]; // @[Bitwise.scala 26:51]
  assign s1_hazard_lo_hi_lo_3 = _s1_hazard_T_21[2]; // @[Bitwise.scala 26:51]
  assign s1_hazard_lo_lo_hi_3 = _s1_hazard_T_21[1]; // @[Bitwise.scala 26:51]
  assign s1_hazard_lo_lo_lo_3 = _s1_hazard_T_21[0]; // @[Bitwise.scala 26:51]
  assign _s1_hazard_T_22 = {s1_hazard_hi_hi_hi_3,s1_hazard_hi_hi_lo_3,s1_hazard_hi_lo_hi_3,s1_hazard_hi_lo_lo_3,s1_hazard_lo_hi_hi_3,s1_hazard_lo_hi_lo_3,s1_hazard_lo_lo_hi_3,s1_hazard_lo_lo_lo_3}; // @[Cat.scala 30:58]
  assign _s1_hazard_T_23 = _s1_hazard_T_12 & _s1_hazard_T_22; // @[DCache.scala 533:38]
  assign _s1_hazard_T_24 = |_s1_hazard_T_23; // @[DCache.scala 533:66]
  assign _s1_hazard_T_25 = pstore1_mask & s1_mask_xwr; // @[DCache.scala 533:77]
  assign _s1_hazard_T_26 = |_s1_hazard_T_25; // @[DCache.scala 533:92]
  assign _s1_hazard_T_27 = s1_write ? _s1_hazard_T_24 : _s1_hazard_T_26; // @[DCache.scala 533:8]
  assign _s1_hazard_T_28 = _s1_hazard_T_2 & _s1_hazard_T_27; // @[DCache.scala 532:65]
  assign _s1_hazard_T_29 = pstore1_valid_likely & _s1_hazard_T_28; // @[DCache.scala 535:27]
  assign _s1_hazard_T_32 = pstore2_addr[11:3] == s1_vaddr[11:3]; // @[DCache.scala 532:31]
  assign s1_hazard_hi_hi_hi_4 = |mask[7]; // @[DCache.scala 1149:66]
  assign s1_hazard_hi_hi_lo_4 = |mask[6]; // @[DCache.scala 1149:66]
  assign s1_hazard_hi_lo_hi_4 = |mask[5]; // @[DCache.scala 1149:66]
  assign s1_hazard_hi_lo_lo_4 = |mask[4]; // @[DCache.scala 1149:66]
  assign s1_hazard_lo_hi_hi_4 = |mask[3]; // @[DCache.scala 1149:66]
  assign s1_hazard_lo_hi_lo_4 = |mask[2]; // @[DCache.scala 1149:66]
  assign s1_hazard_lo_lo_hi_4 = |mask[1]; // @[DCache.scala 1149:66]
  assign s1_hazard_lo_lo_lo_4 = |mask[0]; // @[DCache.scala 1149:66]
  assign _s1_hazard_T_41 = {s1_hazard_hi_hi_hi_4,s1_hazard_hi_hi_lo_4,s1_hazard_hi_lo_hi_4,s1_hazard_hi_lo_lo_4,s1_hazard_lo_hi_hi_4,s1_hazard_lo_hi_lo_4,s1_hazard_lo_lo_hi_4,s1_hazard_lo_lo_lo_4}; // @[Cat.scala 30:58]
  assign s1_hazard_hi_hi_hi_5 = _s1_hazard_T_41[7]; // @[Bitwise.scala 26:51]
  assign s1_hazard_hi_hi_lo_5 = _s1_hazard_T_41[6]; // @[Bitwise.scala 26:51]
  assign s1_hazard_hi_lo_hi_5 = _s1_hazard_T_41[5]; // @[Bitwise.scala 26:51]
  assign s1_hazard_hi_lo_lo_5 = _s1_hazard_T_41[4]; // @[Bitwise.scala 26:51]
  assign s1_hazard_lo_hi_hi_5 = _s1_hazard_T_41[3]; // @[Bitwise.scala 26:51]
  assign s1_hazard_lo_hi_lo_5 = _s1_hazard_T_41[2]; // @[Bitwise.scala 26:51]
  assign s1_hazard_lo_lo_hi_5 = _s1_hazard_T_41[1]; // @[Bitwise.scala 26:51]
  assign s1_hazard_lo_lo_lo_5 = _s1_hazard_T_41[0]; // @[Bitwise.scala 26:51]
  assign _s1_hazard_T_42 = {s1_hazard_hi_hi_hi_5,s1_hazard_hi_hi_lo_5,s1_hazard_hi_lo_hi_5,s1_hazard_hi_lo_lo_5,s1_hazard_lo_hi_hi_5,s1_hazard_lo_hi_lo_5,s1_hazard_lo_lo_hi_5,s1_hazard_lo_lo_lo_5}; // @[Cat.scala 30:58]
  assign _s1_hazard_T_53 = _s1_hazard_T_42 & _s1_hazard_T_22; // @[DCache.scala 533:38]
  assign _s1_hazard_T_54 = |_s1_hazard_T_53; // @[DCache.scala 533:66]
  assign _s1_hazard_T_55 = mask & s1_mask_xwr; // @[DCache.scala 533:77]
  assign _s1_hazard_T_56 = |_s1_hazard_T_55; // @[DCache.scala 533:92]
  assign _s1_hazard_T_57 = s1_write ? _s1_hazard_T_54 : _s1_hazard_T_56; // @[DCache.scala 533:8]
  assign _s1_hazard_T_58 = _s1_hazard_T_32 & _s1_hazard_T_57; // @[DCache.scala 532:65]
  assign _s1_hazard_T_59 = pstore2_valid & _s1_hazard_T_58; // @[DCache.scala 536:21]
  assign s1_hazard = _s1_hazard_T_29 | _s1_hazard_T_59; // @[DCache.scala 535:69]
  assign s1_raw_hazard = s1_read & s1_hazard; // @[DCache.scala 537:31]
  assign _T_262 = s1_valid & s1_raw_hazard; // @[DCache.scala 542:18]
  assign _s2_valid_no_xcpt_T = {io_cpu_s2_xcpt_ma_ld,io_cpu_s2_xcpt_ma_st,io_cpu_s2_xcpt_pf_ld,io_cpu_s2_xcpt_pf_st,io_cpu_s2_xcpt_ae_ld,io_cpu_s2_xcpt_ae_st}; // @[DCache.scala 303:54]
  assign _s2_valid_no_xcpt_T_1 = |_s2_valid_no_xcpt_T; // @[DCache.scala 303:61]
  assign s2_valid_no_xcpt = s2_valid & ~_s2_valid_no_xcpt_T_1; // @[DCache.scala 303:35]
  assign s2_valid_masked = s2_valid_no_xcpt & s2_not_nacked_in_s1; // @[DCache.scala 308:42]
  assign _s2_valid_hit_maybe_flush_pre_data_ecc_and_waw_T_1 = s2_valid_masked & ~s2_meta_error; // @[DCache.scala 368:71]
  assign _c_cat_T_45 = s2_req_cmd == 5'h3; // @[Consts.scala 83:54]
  assign _c_cat_T_46 = s2_write | _c_cat_T_45; // @[Consts.scala 83:47]
  assign _c_cat_T_47 = s2_req_cmd == 5'h6; // @[Consts.scala 83:71]
  assign c_cat_lo = _c_cat_T_46 | _c_cat_T_47; // @[Consts.scala 83:64]
  assign _T_71 = {s2_write,c_cat_lo,s2_hit_state_state}; // @[Cat.scala 30:58]
  assign _T_117 = 4'h3 == _T_71; // @[Misc.scala 48:20]
  assign _T_114 = 4'h2 == _T_71; // @[Misc.scala 48:20]
  assign _T_111 = 4'h1 == _T_71; // @[Misc.scala 48:20]
  assign _T_108 = 4'h7 == _T_71; // @[Misc.scala 48:20]
  assign _T_105 = 4'h6 == _T_71; // @[Misc.scala 48:20]
  assign _T_102 = 4'hf == _T_71; // @[Misc.scala 48:20]
  assign _T_99 = 4'he == _T_71; // @[Misc.scala 48:20]
  assign _T_96 = 4'h0 == _T_71; // @[Misc.scala 48:20]
  assign _T_93 = 4'h5 == _T_71; // @[Misc.scala 48:20]
  assign _T_90 = 4'h4 == _T_71; // @[Misc.scala 48:20]
  assign _T_87 = 4'hd == _T_71; // @[Misc.scala 48:20]
  assign _T_84 = 4'hc == _T_71; // @[Misc.scala 48:20]
  assign _T_103 = _T_102 | _T_99; // @[Misc.scala 34:9]
  assign _T_106 = _T_105 | _T_103; // @[Misc.scala 34:9]
  assign _T_109 = _T_108 | _T_106; // @[Misc.scala 34:9]
  assign _T_112 = _T_111 | _T_109; // @[Misc.scala 34:9]
  assign _T_115 = _T_114 | _T_112; // @[Misc.scala 34:9]
  assign s2_hit = _T_117 | _T_115; // @[Misc.scala 34:9]
  assign s2_valid_hit_maybe_flush_pre_data_ecc_and_waw = _s2_valid_hit_maybe_flush_pre_data_ecc_and_waw_T_1 & s2_hit; // @[DCache.scala 368:89]
  assign _s2_read_T = s2_req_cmd == 5'h0; // @[Consts.scala 81:31]
  assign _s2_read_T_2 = _s2_read_T | _c_cat_T_47; // @[Consts.scala 81:41]
  assign _s2_read_T_4 = _s2_read_T_2 | _s2_write_T_3; // @[Consts.scala 81:58]
  assign s2_read = _s2_read_T_4 | _s2_write_T_21; // @[Consts.scala 81:75]
  assign s2_readwrite = s2_read | s2_write; // @[DCache.scala 325:30]
  assign s2_valid_hit_pre_data_ecc_and_waw = s2_valid_hit_maybe_flush_pre_data_ecc_and_waw & s2_readwrite; // @[DCache.scala 389:89]
  assign _T_86 = _T_84 ? 2'h1 : 2'h0; // @[Misc.scala 34:36]
  assign _T_89 = _T_87 ? 2'h2 : _T_86; // @[Misc.scala 34:36]
  assign _T_92 = _T_90 ? 2'h1 : _T_89; // @[Misc.scala 34:36]
  assign _T_95 = _T_93 ? 2'h2 : _T_92; // @[Misc.scala 34:36]
  assign _T_98 = _T_96 ? 2'h0 : _T_95; // @[Misc.scala 34:36]
  assign _T_101 = _T_99 ? 2'h3 : _T_98; // @[Misc.scala 34:36]
  assign _T_104 = _T_102 ? 2'h3 : _T_101; // @[Misc.scala 34:36]
  assign _T_107 = _T_105 ? 2'h2 : _T_104; // @[Misc.scala 34:36]
  assign _T_110 = _T_108 ? 2'h3 : _T_107; // @[Misc.scala 34:36]
  assign _T_113 = _T_111 ? 2'h1 : _T_110; // @[Misc.scala 34:36]
  assign _T_116 = _T_114 ? 2'h2 : _T_113; // @[Misc.scala 34:36]
  assign s2_grow_param = _T_117 ? 2'h3 : _T_116; // @[Misc.scala 34:36]
  assign _s2_update_meta_T = s2_hit_state_state == s2_grow_param; // @[Metadata.scala 45:46]
  assign s2_update_meta = ~_s2_update_meta_T; // @[Metadata.scala 46:40]
  assign _T_241 = s2_valid_hit_pre_data_ecc_and_waw & s2_update_meta; // @[DCache.scala 417:62]
  assign _T_242 = io_cpu_s2_nack | _T_241; // @[DCache.scala 417:24]
  assign s1_readwrite = s1_read | s1_write; // @[DCache.scala 190:30]
  assign _s1_flush_line_T = s1_req_cmd == 5'h5; // @[DCache.scala 192:34]
  assign s1_flush_line = _s1_flush_line_T & s1_req_size[0]; // @[DCache.scala 192:50]
  assign _s1_cmd_uses_tlb_T = s1_readwrite | s1_flush_line; // @[DCache.scala 248:38]
  assign _s1_cmd_uses_tlb_T_1 = s1_req_cmd == 5'h17; // @[DCache.scala 248:69]
  assign s1_cmd_uses_tlb = _s1_cmd_uses_tlb_T | _s1_cmd_uses_tlb_T_1; // @[DCache.scala 248:55]
  assign _T_13 = s1_valid & s1_cmd_uses_tlb; // @[DCache.scala 254:39]
  assign _T_14 = _T_13 & tlb_io_resp_miss; // @[DCache.scala 254:58]
  assign _GEN_117 = _T_242 | _T_14; // @[DCache.scala 417:82]
  assign _GEN_141 = _T_262 | _GEN_117; // @[DCache.scala 542:36]
  assign _GEN_283 = probeNack | _GEN_141; // @[DCache.scala 810:24]
  assign s1_nack = s2_probe ? _GEN_283 : _GEN_141; // @[DCache.scala 795:21]
  assign s1_valid_not_nacked = s1_valid & ~s1_nack; // @[DCache.scala 167:38]
  assign s0_clk_en = metaArb_io_out_valid & ~metaArb_io_out_bits_write; // @[DCache.scala 170:40]
  assign s0_req_addr_hi = metaArb_io_out_bits_addr[39:6]; // @[DCache.scala 173:47]
  assign s0_req_addr_lo = io_cpu_req_bits_addr[5:0]; // @[DCache.scala 173:84]
  assign s0_req_addr = {s0_req_addr_hi,s0_req_addr_lo}; // @[Cat.scala 30:58]
  assign s0_req_phys = ~metaArb_io_in_7_ready | io_cpu_req_bits_phys; // @[DCache.scala 175:34]
  assign s1_sfence = s1_req_cmd == 5'h14; // @[DCache.scala 191:30]
  assign inWriteback = _T_308 | _T_307; // @[package.scala 72:59]
  assign _io_cpu_req_ready_T = release_state == 4'h0; // @[DCache.scala 211:38]
  assign _io_cpu_req_ready_T_2 = _io_cpu_req_ready_T & ~cached_grant_wait; // @[DCache.scala 211:51]
  assign _io_cpu_req_ready_T_4 = _io_cpu_req_ready_T_2 & ~s1_nack; // @[DCache.scala 211:73]
  assign _s0_read_T = io_cpu_req_bits_cmd == 5'h0; // @[Consts.scala 81:31]
  assign _s0_read_T_1 = io_cpu_req_bits_cmd == 5'h6; // @[Consts.scala 81:48]
  assign _s0_read_T_2 = _s0_read_T | _s0_read_T_1; // @[Consts.scala 81:41]
  assign _s0_read_T_3 = io_cpu_req_bits_cmd == 5'h7; // @[Consts.scala 81:65]
  assign _s0_read_T_4 = _s0_read_T_2 | _s0_read_T_3; // @[Consts.scala 81:58]
  assign _s0_read_T_5 = io_cpu_req_bits_cmd == 5'h4; // @[package.scala 15:47]
  assign _s0_read_T_6 = io_cpu_req_bits_cmd == 5'h9; // @[package.scala 15:47]
  assign _s0_read_T_7 = io_cpu_req_bits_cmd == 5'ha; // @[package.scala 15:47]
  assign _s0_read_T_8 = io_cpu_req_bits_cmd == 5'hb; // @[package.scala 15:47]
  assign _s0_read_T_9 = _s0_read_T_5 | _s0_read_T_6; // @[package.scala 72:59]
  assign _s0_read_T_10 = _s0_read_T_9 | _s0_read_T_7; // @[package.scala 72:59]
  assign _s0_read_T_11 = _s0_read_T_10 | _s0_read_T_8; // @[package.scala 72:59]
  assign _s0_read_T_12 = io_cpu_req_bits_cmd == 5'h8; // @[package.scala 15:47]
  assign _s0_read_T_13 = io_cpu_req_bits_cmd == 5'hc; // @[package.scala 15:47]
  assign _s0_read_T_14 = io_cpu_req_bits_cmd == 5'hd; // @[package.scala 15:47]
  assign _s0_read_T_15 = io_cpu_req_bits_cmd == 5'he; // @[package.scala 15:47]
  assign _s0_read_T_16 = io_cpu_req_bits_cmd == 5'hf; // @[package.scala 15:47]
  assign _s0_read_T_17 = _s0_read_T_12 | _s0_read_T_13; // @[package.scala 72:59]
  assign _s0_read_T_18 = _s0_read_T_17 | _s0_read_T_14; // @[package.scala 72:59]
  assign _s0_read_T_19 = _s0_read_T_18 | _s0_read_T_15; // @[package.scala 72:59]
  assign _s0_read_T_20 = _s0_read_T_19 | _s0_read_T_16; // @[package.scala 72:59]
  assign _s0_read_T_21 = _s0_read_T_11 | _s0_read_T_20; // @[Consts.scala 79:44]
  assign s0_read = _s0_read_T_4 | _s0_read_T_21; // @[Consts.scala 81:75]
  assign _dataArb_io_in_3_valid_res_T = io_cpu_req_bits_cmd == 5'h1; // @[package.scala 15:47]
  assign _dataArb_io_in_3_valid_res_T_1 = io_cpu_req_bits_cmd == 5'h3; // @[package.scala 15:47]
  assign _dataArb_io_in_3_valid_res_T_2 = _dataArb_io_in_3_valid_res_T | _dataArb_io_in_3_valid_res_T_1; // @[package.scala 72:59]
  assign res = ~_dataArb_io_in_3_valid_res_T_2; // @[DCache.scala 1153:15]
  assign _dataArb_io_in_3_valid_T_24 = io_cpu_req_bits_cmd == 5'h11; // @[Consts.scala 82:49]
  assign _dataArb_io_in_3_valid_T_25 = _dataArb_io_in_3_valid_res_T | _dataArb_io_in_3_valid_T_24; // @[Consts.scala 82:42]
  assign _dataArb_io_in_3_valid_T_27 = _dataArb_io_in_3_valid_T_25 | _s0_read_T_3; // @[Consts.scala 82:59]
  assign _dataArb_io_in_3_valid_T_45 = _dataArb_io_in_3_valid_T_27 | _s0_read_T_21; // @[Consts.scala 82:76]
  assign _dataArb_io_in_3_valid_T_49 = _dataArb_io_in_3_valid_T_45 & _dataArb_io_in_3_valid_T_24; // @[DCache.scala 1159:23]
  assign _dataArb_io_in_3_valid_T_50 = s0_read | _dataArb_io_in_3_valid_T_49; // @[DCache.scala 1158:21]
  assign _dataArb_io_in_3_valid_T_52 = ~_dataArb_io_in_3_valid_T_50 | res; // @[DCache.scala 1154:28]
  assign _dataArb_io_in_3_valid_T_54 = _dataArb_io_in_3_valid_T_52 | reset; // @[DCache.scala 1154:11]
  assign _dataArb_io_in_3_valid_T_56 = io_cpu_req_valid & res; // @[DCache.scala 220:46]
  assign dataArb_io_in_3_bits_addr_hi = io_cpu_req_bits_addr[39:12]; // @[DCache.scala 223:89]
  assign dataArb_io_in_3_bits_addr_lo = io_cpu_req_bits_addr[11:0]; // @[DCache.scala 223:120]
  assign _dataArb_io_in_3_bits_addr_T = {dataArb_io_in_3_bits_addr_hi,dataArb_io_in_3_bits_addr_lo}; // @[Cat.scala 30:58]
  assign _T_4 = ~dataArb_io_in_3_ready & s0_read; // @[DCache.scala 236:33]
  assign _GEN_28 = _T_4 ? 1'h0 : _io_cpu_req_ready_T_4; // @[DCache.scala 236:45]
  assign _s1_did_read_T_51 = io_cpu_req_valid & _dataArb_io_in_3_valid_T_50; // @[DCache.scala 237:75]
  assign _s1_did_read_T_52 = dataArb_io_in_3_ready & _s1_did_read_T_51; // @[DCache.scala 237:54]
  assign _GEN_31 = metaArb_io_in_7_ready ? _GEN_28 : 1'h0; // @[DCache.scala 245:34]
  assign _T_8 = ~tlb_io_req_ready & ~tlb_io_ptw_resp_valid; // @[DCache.scala 253:27]
  assign _T_10 = _T_8 & ~io_cpu_req_bits_phys; // @[DCache.scala 253:53]
  assign _GEN_32 = _T_10 ? 1'h0 : _GEN_31; // @[DCache.scala 253:79]
  assign s1_paddr_hi = tlb_io_resp_paddr[31:12]; // @[DCache.scala 269:99]
  assign s1_paddr = {s1_paddr_hi,s1_vaddr_lo}; // @[Cat.scala 30:58]
  assign _WIRE_2 = tag_array_0_s1_meta_data;
  assign s1_meta_uncorrected_0_tag = _WIRE_2[19:0]; // @[DCache.scala 286:80]
  assign s1_meta_uncorrected_0_coh_state = _WIRE_2[21:20]; // @[DCache.scala 286:80]
  assign _WIRE_3 = tag_array_1_s1_meta_data;
  assign s1_meta_uncorrected_1_tag = _WIRE_3[19:0]; // @[DCache.scala 286:80]
  assign s1_meta_uncorrected_1_coh_state = _WIRE_3[21:20]; // @[DCache.scala 286:80]
  assign _WIRE_4 = tag_array_2_s1_meta_data;
  assign s1_meta_uncorrected_2_tag = _WIRE_4[19:0]; // @[DCache.scala 286:80]
  assign s1_meta_uncorrected_2_coh_state = _WIRE_4[21:20]; // @[DCache.scala 286:80]
  assign _WIRE_5 = tag_array_3_s1_meta_data;
  assign s1_meta_uncorrected_3_tag = _WIRE_5[19:0]; // @[DCache.scala 286:80]
  assign s1_meta_uncorrected_3_coh_state = _WIRE_5[21:20]; // @[DCache.scala 286:80]
  assign s1_tag = s1_paddr[31:12]; // @[DCache.scala 287:29]
  assign _T_32 = s1_meta_uncorrected_0_coh_state > 2'h0; // @[Metadata.scala 49:45]
  assign _T_33 = s1_meta_uncorrected_0_tag == s1_tag; // @[DCache.scala 288:83]
  assign lo_lo = _T_32 & _T_33; // @[DCache.scala 288:74]
  assign _T_34 = s1_meta_uncorrected_1_coh_state > 2'h0; // @[Metadata.scala 49:45]
  assign _T_35 = s1_meta_uncorrected_1_tag == s1_tag; // @[DCache.scala 288:83]
  assign lo_hi = _T_34 & _T_35; // @[DCache.scala 288:74]
  assign _T_36 = s1_meta_uncorrected_2_coh_state > 2'h0; // @[Metadata.scala 49:45]
  assign _T_37 = s1_meta_uncorrected_2_tag == s1_tag; // @[DCache.scala 288:83]
  assign hi_lo = _T_36 & _T_37; // @[DCache.scala 288:74]
  assign _T_38 = s1_meta_uncorrected_3_coh_state > 2'h0; // @[Metadata.scala 49:45]
  assign _T_39 = s1_meta_uncorrected_3_tag == s1_tag; // @[DCache.scala 288:83]
  assign hi_hi = _T_38 & _T_39; // @[DCache.scala 288:74]
  assign s1_meta_hit_way = {hi_hi,hi_lo,lo_hi,lo_lo}; // @[Cat.scala 30:58]
  assign _T_42 = _T_33 & ~s1_flush_valid; // @[DCache.scala 290:59]
  assign _T_43 = _T_42 ? s1_meta_uncorrected_0_coh_state : 2'h0; // @[DCache.scala 290:41]
  assign _T_46 = _T_35 & ~s1_flush_valid; // @[DCache.scala 290:59]
  assign _T_47 = _T_46 ? s1_meta_uncorrected_1_coh_state : 2'h0; // @[DCache.scala 290:41]
  assign _T_50 = _T_37 & ~s1_flush_valid; // @[DCache.scala 290:59]
  assign _T_51 = _T_50 ? s1_meta_uncorrected_2_coh_state : 2'h0; // @[DCache.scala 290:41]
  assign _T_54 = _T_39 & ~s1_flush_valid; // @[DCache.scala 290:59]
  assign _T_55 = _T_54 ? s1_meta_uncorrected_3_coh_state : 2'h0; // @[DCache.scala 290:41]
  assign _T_56 = _T_43 | _T_47; // @[DCache.scala 291:19]
  assign _T_57 = _T_56 | _T_51; // @[DCache.scala 291:19]
  assign s1_meta_hit_state_state = _T_57 | _T_55; // @[DCache.scala 291:19]
  assign s2_hit_valid = s2_hit_state_state > 2'h0; // @[Metadata.scala 49:45]
  assign s2_victim_way = 4'h1 << s2_victim_way_r; // @[OneHot.scala 58:35]
  assign s2_victim_or_hit_way = s2_hit_valid ? s2_hit_way : s2_victim_way; // @[DCache.scala 403:33]
  assign releaseWay = _T_312 ? s2_victim_or_hit_way : s2_probe_way; // @[DCache.scala 834:102]
  assign s1_data_way_x35 = inWriteback ? releaseWay : s1_meta_hit_way; // @[DCache.scala 294:61]
  assign tl_d_data_encoded_lo_lo_lo = auto_out_d_bits_data[7:0]; // @[package.scala 202:50]
  assign tl_d_data_encoded_lo_lo_hi = auto_out_d_bits_data[15:8]; // @[package.scala 202:50]
  assign tl_d_data_encoded_lo_hi_lo = auto_out_d_bits_data[23:16]; // @[package.scala 202:50]
  assign tl_d_data_encoded_lo_hi_hi = auto_out_d_bits_data[31:24]; // @[package.scala 202:50]
  assign tl_d_data_encoded_hi_lo_lo = auto_out_d_bits_data[39:32]; // @[package.scala 202:50]
  assign tl_d_data_encoded_hi_lo_hi = auto_out_d_bits_data[47:40]; // @[package.scala 202:50]
  assign tl_d_data_encoded_hi_hi_lo = auto_out_d_bits_data[55:48]; // @[package.scala 202:50]
  assign tl_d_data_encoded_hi_hi_hi = auto_out_d_bits_data[63:56]; // @[package.scala 202:50]
  assign tl_d_data_encoded_lo = {tl_d_data_encoded_lo_hi_hi,tl_d_data_encoded_lo_hi_lo,tl_d_data_encoded_lo_lo_hi,tl_d_data_encoded_lo_lo_lo}; // @[Cat.scala 30:58]
  assign tl_d_data_encoded_hi = {tl_d_data_encoded_hi_hi_hi,tl_d_data_encoded_hi_hi_lo,tl_d_data_encoded_hi_lo_hi,tl_d_data_encoded_hi_lo_lo}; // @[Cat.scala 30:58]
  assign _tl_d_data_encoded_T = {tl_d_data_encoded_hi_hi_hi,tl_d_data_encoded_hi_hi_lo,tl_d_data_encoded_hi_lo_hi,tl_d_data_encoded_hi_lo_lo,tl_d_data_encoded_lo_hi_hi,tl_d_data_encoded_lo_hi_lo,tl_d_data_encoded_lo_lo_hi,tl_d_data_encoded_lo_lo_lo}; // @[Cat.scala 30:58]
  assign _T_61 = s1_valid_masked & _s1_write_T_1; // @[DCache.scala 300:28]
  assign _T_65 = &8'hff; // @[DCache.scala 300:93]
  assign _T_66 = ~_T_61 | _T_65; // @[DCache.scala 300:53]
  assign _T_68 = _T_66 | reset; // @[DCache.scala 300:9]
  assign s2_valid_x37 = s1_valid_masked & ~s1_sfence; // @[DCache.scala 302:43]
  assign _s2_cmd_flush_all_T = s2_req_cmd == 5'h5; // @[DCache.scala 311:37]
  assign s2_cmd_flush_line = _s2_cmd_flush_all_T & s2_req_size[0]; // @[DCache.scala 312:54]
  assign _T_70 = s1_valid_not_nacked | s1_flush_valid; // @[DCache.scala 316:29]
  assign _s2_pma_T_cacheable = tlb_io_resp_cacheable; // @[DCache.scala 320:18]
  assign s2_vaddr_hi = s2_vaddr_r[39:12]; // @[DCache.scala 322:81]
  assign s2_vaddr_lo = s2_req_addr[11:0]; // @[DCache.scala 322:103]
  assign s2_vaddr = {s2_vaddr_hi,s2_vaddr_lo}; // @[Cat.scala 30:58]
  assign s1_meta_clk_en = _T_70 | s1_probe; // @[DCache.scala 328:62]
  assign s2_meta_corrected_0_tag = s2_meta_corrected_r[19:0]; // @[DCache.scala 332:99]
  assign s2_meta_corrected_0_coh_state = s2_meta_corrected_r[21:20]; // @[DCache.scala 332:99]
  assign s2_meta_corrected_1_tag = s2_meta_corrected_r_1[19:0]; // @[DCache.scala 332:99]
  assign s2_meta_corrected_1_coh_state = s2_meta_corrected_r_1[21:20]; // @[DCache.scala 332:99]
  assign s2_meta_corrected_2_tag = s2_meta_corrected_r_2[19:0]; // @[DCache.scala 332:99]
  assign s2_meta_corrected_2_coh_state = s2_meta_corrected_r_2[21:20]; // @[DCache.scala 332:99]
  assign s2_meta_corrected_3_tag = s2_meta_corrected_r_3[19:0]; // @[DCache.scala 332:99]
  assign s2_meta_corrected_3_coh_state = s2_meta_corrected_r_3[21:20]; // @[DCache.scala 332:99]
  assign s2_flush_valid = s2_flush_valid_pre_tag_ecc & ~s2_meta_error; // @[DCache.scala 334:51]
  assign _s2_data_en_T = s1_valid | inWriteback; // @[DCache.scala 337:23]
  assign en = _s2_data_en_T | io_cpu_replay_next; // @[DCache.scala 337:38]
  assign _s2_data_word_en_T = s1_did_read & s1_read_mask; // @[DCache.scala 338:63]
  assign word_en = inWriteback | _s2_data_word_en_T; // @[DCache.scala 338:22]
  assign s1_all_data_ways_0 = data_io_resp_0; // @[DCache.scala 296:29 DCache.scala 296:29]
  assign s1_all_data_ways_1 = data_io_resp_1; // @[DCache.scala 296:29 DCache.scala 296:29]
  assign s1_all_data_ways_2 = data_io_resp_2; // @[DCache.scala 296:29 DCache.scala 296:29]
  assign s1_all_data_ways_3 = data_io_resp_3; // @[DCache.scala 296:29 DCache.scala 296:29]
  assign s1_word_en = io_cpu_replay_next ? 1'h1 : word_en; // @[DCache.scala 348:27]
  assign grantIsUncachedData = auto_out_d_bits_opcode == 3'h1; // @[package.scala 15:47]
  assign _T_293 = blockUncachedGrant | s1_valid; // @[DCache.scala 723:54]
  assign _T_294 = grantIsUncachedData & _T_293; // @[DCache.scala 723:31]
  assign grantIsRefill = auto_out_d_bits_opcode == 3'h5; // @[DCache.scala 637:29]
  assign _T_292 = grantIsRefill & ~dataArb_io_in_1_ready; // @[DCache.scala 693:23]
  assign _grantIsCached_T = auto_out_d_bits_opcode == 3'h4; // @[package.scala 15:47]
  assign grantIsCached = _grantIsCached_T | grantIsRefill; // @[package.scala 72:59]
  assign d_first = counter == 9'h0; // @[Edges.scala 230:25]
  assign _bundleOut_0_d_ready_T_1 = ~d_first | auto_out_e_ready; // @[DCache.scala 642:50]
  assign canAcceptCachedGrant = ~_T_312; // @[DCache.scala 641:30]
  assign _bundleOut_0_d_ready_T_2 = _bundleOut_0_d_ready_T_1 & canAcceptCachedGrant; // @[DCache.scala 642:69]
  assign _bundleOut_0_d_ready_T_3 = grantIsCached ? _bundleOut_0_d_ready_T_2 : 1'h1; // @[DCache.scala 642:24]
  assign _GEN_233 = _T_292 ? 1'h0 : _bundleOut_0_d_ready_T_3; // @[DCache.scala 693:51]
  assign tl_out__d_ready = _T_294 ? 1'h0 : _GEN_233; // @[DCache.scala 723:68]
  assign _T_271 = tl_out__d_ready & auto_out_d_valid; // @[Decoupled.scala 40:37]
  assign _T_267 = auto_out_d_bits_opcode == 3'h0; // @[package.scala 15:47]
  assign _T_269 = grantIsUncachedData | _T_267; // @[package.scala 72:59]
  assign _T_268 = auto_out_d_bits_opcode == 3'h2; // @[package.scala 15:47]
  assign grantIsUncached = _T_269 | _T_268; // @[package.scala 72:59]
  assign _GEN_189 = grantIsUncachedData ? 5'h10 : {{1'd0}, s1_data_way_x35}; // @[DCache.scala 662:34]
  assign _GEN_198 = grantIsUncached ? _GEN_189 : {{1'd0}, s1_data_way_x35}; // @[DCache.scala 655:35]
  assign _GEN_211 = grantIsCached ? {{1'd0}, s1_data_way_x35} : _GEN_198; // @[DCache.scala 646:26]
  assign s1_data_way = _T_271 ? _GEN_211 : {{1'd0}, s1_data_way_x35}; // @[DCache.scala 645:26]
  assign _s2_data_T_1 = s1_word_en ? s1_data_way : 5'h0; // @[DCache.scala 350:28]
  assign _s2_data_T_7 = _s2_data_T_1[0] ? s1_all_data_ways_0 : 64'h0; // @[Mux.scala 27:72]
  assign _s2_data_T_8 = _s2_data_T_1[1] ? s1_all_data_ways_1 : 64'h0; // @[Mux.scala 27:72]
  assign _s2_data_T_9 = _s2_data_T_1[2] ? s1_all_data_ways_2 : 64'h0; // @[Mux.scala 27:72]
  assign _s2_data_T_10 = _s2_data_T_1[3] ? s1_all_data_ways_3 : 64'h0; // @[Mux.scala 27:72]
  assign _s2_data_T_11 = _s2_data_T_1[4] ? _tl_d_data_encoded_T : 64'h0; // @[Mux.scala 27:72]
  assign _s2_data_T_12 = _s2_data_T_7 | _s2_data_T_8; // @[Mux.scala 27:72]
  assign _s2_data_T_13 = _s2_data_T_12 | _s2_data_T_9; // @[Mux.scala 27:72]
  assign _s2_data_T_14 = _s2_data_T_13 | _s2_data_T_10; // @[Mux.scala 27:72]
  assign _s2_data_T_15 = _s2_data_T_14 | _s2_data_T_11; // @[Mux.scala 27:72]
  assign s2_data_uncorrected_lo_lo_lo = s2_data[7:0]; // @[package.scala 202:50]
  assign s2_data_uncorrected_lo_lo_hi = s2_data[15:8]; // @[package.scala 202:50]
  assign s2_data_uncorrected_lo_hi_lo = s2_data[23:16]; // @[package.scala 202:50]
  assign s2_data_uncorrected_lo_hi_hi = s2_data[31:24]; // @[package.scala 202:50]
  assign s2_data_uncorrected_hi_lo_lo = s2_data[39:32]; // @[package.scala 202:50]
  assign s2_data_uncorrected_hi_lo_hi = s2_data[47:40]; // @[package.scala 202:50]
  assign s2_data_uncorrected_hi_hi_lo = s2_data[55:48]; // @[package.scala 202:50]
  assign s2_data_uncorrected_hi_hi_hi = s2_data[63:56]; // @[package.scala 202:50]
  assign s2_data_corrected_lo = {s2_data_uncorrected_lo_hi_hi,s2_data_uncorrected_lo_hi_lo,s2_data_uncorrected_lo_lo_hi,s2_data_uncorrected_lo_lo_lo}; // @[Cat.scala 30:58]
  assign s2_data_corrected_hi = {s2_data_uncorrected_hi_hi_hi,s2_data_uncorrected_hi_hi_lo,s2_data_uncorrected_hi_lo_hi,s2_data_uncorrected_hi_lo_lo}; // @[Cat.scala 30:58]
  assign s2_data_corrected = {s2_data_uncorrected_hi_hi_hi,s2_data_uncorrected_hi_hi_lo,s2_data_uncorrected_hi_lo_hi,s2_data_uncorrected_hi_lo_lo,s2_data_uncorrected_lo_hi_hi,s2_data_uncorrected_lo_hi_lo,s2_data_uncorrected_lo_lo_hi,s2_data_uncorrected_lo_lo_lo}; // @[Cat.scala 30:58]
  assign s2_valid_flush_line = s2_valid_hit_maybe_flush_pre_data_ecc_and_waw & s2_cmd_flush_line; // @[DCache.scala 390:75]
  assign _s2_valid_miss_T = s2_valid_masked & s2_readwrite; // @[DCache.scala 394:39]
  assign _s2_valid_miss_T_2 = _s2_valid_miss_T & ~s2_meta_error; // @[DCache.scala 394:55]
  assign s2_valid_miss = _s2_valid_miss_T_2 & ~s2_hit; // @[DCache.scala 394:73]
  assign s2_uncached = ~s2_pma_cacheable; // @[DCache.scala 395:21]
  assign _s2_valid_cached_miss_T_1 = s2_valid_miss & ~s2_uncached; // @[DCache.scala 396:44]
  assign _s2_valid_cached_miss_T_2 = |uncachedInFlight_0; // @[DCache.scala 396:88]
  assign s2_valid_cached_miss = _s2_valid_cached_miss_T_1 & ~_s2_valid_cached_miss_T_2; // @[DCache.scala 396:60]
  assign _s2_want_victimize_T = s2_valid_cached_miss | s2_valid_flush_line; // @[DCache.scala 398:79]
  assign s2_want_victimize = _s2_want_victimize_T | s2_flush_valid; // @[DCache.scala 398:125]
  assign _s2_valid_uncached_pending_T = s2_valid_miss & s2_uncached; // @[DCache.scala 401:49]
  assign _s2_valid_uncached_pending_T_1 = &uncachedInFlight_0; // @[DCache.scala 401:92]
  assign s2_valid_uncached_pending = _s2_valid_uncached_pending_T & ~_s2_valid_uncached_pending_T_1; // @[DCache.scala 401:64]
  assign s1_victim_way = lfsr[1:0]; // @[package.scala 154:13]
  assign _s2_victim_tag_T_6 = s2_victim_way[0] ? s2_meta_corrected_0_tag : 20'h0; // @[Mux.scala 27:72]
  assign _s2_victim_tag_T_7 = s2_victim_way[1] ? s2_meta_corrected_1_tag : 20'h0; // @[Mux.scala 27:72]
  assign _s2_victim_tag_T_8 = s2_victim_way[2] ? s2_meta_corrected_2_tag : 20'h0; // @[Mux.scala 27:72]
  assign _s2_victim_tag_T_9 = s2_victim_way[3] ? s2_meta_corrected_3_tag : 20'h0; // @[Mux.scala 27:72]
  assign _s2_victim_tag_T_10 = _s2_victim_tag_T_6 | _s2_victim_tag_T_7; // @[Mux.scala 27:72]
  assign _s2_victim_tag_T_11 = _s2_victim_tag_T_10 | _s2_victim_tag_T_8; // @[Mux.scala 27:72]
  assign _s2_victim_tag_T_12 = _s2_victim_tag_T_11 | _s2_victim_tag_T_9; // @[Mux.scala 27:72]
  assign _s2_victim_tag_T_13 = s2_victim_way[0] ? s2_meta_corrected_0_coh_state : 2'h0; // @[Mux.scala 27:72]
  assign _s2_victim_tag_T_14 = s2_victim_way[1] ? s2_meta_corrected_1_coh_state : 2'h0; // @[Mux.scala 27:72]
  assign _s2_victim_tag_T_15 = s2_victim_way[2] ? s2_meta_corrected_2_coh_state : 2'h0; // @[Mux.scala 27:72]
  assign _s2_victim_tag_T_16 = s2_victim_way[3] ? s2_meta_corrected_3_coh_state : 2'h0; // @[Mux.scala 27:72]
  assign _s2_victim_tag_T_17 = _s2_victim_tag_T_13 | _s2_victim_tag_T_14; // @[Mux.scala 27:72]
  assign _s2_victim_tag_T_18 = _s2_victim_tag_T_17 | _s2_victim_tag_T_15; // @[Mux.scala 27:72]
  assign _s2_victim_tag_T_19 = _s2_victim_tag_T_18 | _s2_victim_tag_T_16; // @[Mux.scala 27:72]
  assign s2_victim_tag = s2_valid_flush_line ? s2_req_addr[31:12] : _s2_victim_tag_T_12; // @[DCache.scala 404:26]
  assign s2_victim_state_state = s2_hit_valid ? s2_hit_state_state : _s2_victim_tag_T_19; // @[DCache.scala 405:28]
  assign _T_133 = _T_131 ? 3'h5 : 3'h0; // @[Misc.scala 37:36]
  assign _T_137 = _T_135 ? 3'h2 : _T_133; // @[Misc.scala 37:36]
  assign _T_141 = _T_139 ? 3'h1 : _T_137; // @[Misc.scala 37:36]
  assign _T_145 = _T_143 ? 3'h1 : _T_141; // @[Misc.scala 37:36]
  assign _T_149 = _T_147 ? 3'h5 : _T_145; // @[Misc.scala 37:36]
  assign _T_153 = _T_151 ? 3'h4 : _T_149; // @[Misc.scala 37:36]
  assign _T_154 = _T_151 ? 2'h1 : 2'h0; // @[Misc.scala 37:63]
  assign _T_157 = _T_155 ? 3'h0 : _T_153; // @[Misc.scala 37:36]
  assign _T_158 = _T_155 ? 2'h1 : _T_154; // @[Misc.scala 37:63]
  assign _T_161 = _T_159 ? 3'h0 : _T_157; // @[Misc.scala 37:36]
  assign _T_162 = _T_159 ? 2'h1 : _T_158; // @[Misc.scala 37:63]
  assign _T_165 = _T_163 ? 3'h5 : _T_161; // @[Misc.scala 37:36]
  assign _T_166 = _T_163 ? 2'h0 : _T_162; // @[Misc.scala 37:63]
  assign _T_169 = _T_167 ? 3'h4 : _T_165; // @[Misc.scala 37:36]
  assign _T_170 = _T_167 ? 2'h1 : _T_166; // @[Misc.scala 37:63]
  assign _T_173 = _T_171 ? 3'h3 : _T_169; // @[Misc.scala 37:36]
  assign _T_174 = _T_171 ? 2'h2 : _T_170; // @[Misc.scala 37:63]
  assign s2_report_param = _T_175 ? 3'h3 : _T_173; // @[Misc.scala 37:36]
  assign probeNewCoh_state = _T_175 ? 2'h2 : _T_174; // @[Misc.scala 37:63]
  assign _T_182 = {2'h2,s2_victim_state_state}; // @[Cat.scala 30:58]
  assign _T_195 = 4'h8 == _T_182; // @[Misc.scala 55:20]
  assign _T_197 = _T_195 ? 3'h5 : 3'h0; // @[Misc.scala 37:36]
  assign _T_199 = 4'h9 == _T_182; // @[Misc.scala 55:20]
  assign _T_201 = _T_199 ? 3'h2 : _T_197; // @[Misc.scala 37:36]
  assign _T_203 = 4'ha == _T_182; // @[Misc.scala 55:20]
  assign _T_205 = _T_203 ? 3'h1 : _T_201; // @[Misc.scala 37:36]
  assign _T_207 = 4'hb == _T_182; // @[Misc.scala 55:20]
  assign _T_209 = _T_207 ? 3'h1 : _T_205; // @[Misc.scala 37:36]
  assign _T_211 = 4'h4 == _T_182; // @[Misc.scala 55:20]
  assign _T_212 = _T_211 ? 1'h0 : _T_207; // @[Misc.scala 37:9]
  assign _T_213 = _T_211 ? 3'h5 : _T_209; // @[Misc.scala 37:36]
  assign _T_215 = 4'h5 == _T_182; // @[Misc.scala 55:20]
  assign _T_216 = _T_215 ? 1'h0 : _T_212; // @[Misc.scala 37:9]
  assign _T_217 = _T_215 ? 3'h4 : _T_213; // @[Misc.scala 37:36]
  assign _T_218 = _T_215 ? 2'h1 : 2'h0; // @[Misc.scala 37:63]
  assign _T_219 = 4'h6 == _T_182; // @[Misc.scala 55:20]
  assign _T_220 = _T_219 ? 1'h0 : _T_216; // @[Misc.scala 37:9]
  assign _T_221 = _T_219 ? 3'h0 : _T_217; // @[Misc.scala 37:36]
  assign _T_222 = _T_219 ? 2'h1 : _T_218; // @[Misc.scala 37:63]
  assign _T_223 = 4'h7 == _T_182; // @[Misc.scala 55:20]
  assign _T_224 = _T_223 | _T_220; // @[Misc.scala 37:9]
  assign _T_225 = _T_223 ? 3'h0 : _T_221; // @[Misc.scala 37:36]
  assign _T_226 = _T_223 ? 2'h1 : _T_222; // @[Misc.scala 37:63]
  assign _T_227 = 4'h0 == _T_182; // @[Misc.scala 55:20]
  assign _T_228 = _T_227 ? 1'h0 : _T_224; // @[Misc.scala 37:9]
  assign _T_229 = _T_227 ? 3'h5 : _T_225; // @[Misc.scala 37:36]
  assign _T_230 = _T_227 ? 2'h0 : _T_226; // @[Misc.scala 37:63]
  assign _T_231 = 4'h1 == _T_182; // @[Misc.scala 55:20]
  assign _T_232 = _T_231 ? 1'h0 : _T_228; // @[Misc.scala 37:9]
  assign _T_233 = _T_231 ? 3'h4 : _T_229; // @[Misc.scala 37:36]
  assign _T_234 = _T_231 ? 2'h1 : _T_230; // @[Misc.scala 37:63]
  assign _T_235 = 4'h2 == _T_182; // @[Misc.scala 55:20]
  assign _T_236 = _T_235 ? 1'h0 : _T_232; // @[Misc.scala 37:9]
  assign _T_237 = _T_235 ? 3'h3 : _T_233; // @[Misc.scala 37:36]
  assign _T_238 = _T_235 ? 2'h2 : _T_234; // @[Misc.scala 37:63]
  assign _T_239 = 4'h3 == _T_182; // @[Misc.scala 55:20]
  assign s2_victim_dirty = _T_239 | _T_236; // @[Misc.scala 37:9]
  assign s2_shrink_param = _T_239 ? 3'h3 : _T_237; // @[Misc.scala 37:36]
  assign voluntaryNewCoh_state = _T_239 ? 2'h2 : _T_238; // @[Misc.scala 37:63]
  assign s2_dont_nack_uncached = s2_valid_uncached_pending & auto_out_a_ready; // @[DCache.scala 411:57]
  assign _s2_dont_nack_misc_T_10 = s2_req_cmd == 5'h17; // @[DCache.scala 415:17]
  assign s2_dont_nack_misc = _s2_valid_hit_maybe_flush_pre_data_ecc_and_waw_T_1 & _s2_dont_nack_misc_T_10; // @[DCache.scala 412:61]
  assign _io_cpu_s2_nack_T_1 = s2_valid_no_xcpt & ~s2_dont_nack_uncached; // @[DCache.scala 416:38]
  assign _io_cpu_s2_nack_T_3 = _io_cpu_s2_nack_T_1 & ~s2_dont_nack_misc; // @[DCache.scala 416:64]
  assign _metaArb_io_in_1_valid_T = s2_valid_masked | s2_flush_valid_pre_tag_ecc; // @[DCache.scala 421:63]
  assign _metaArb_io_in_1_valid_T_1 = _metaArb_io_in_1_valid_T | s2_probe; // @[DCache.scala 421:93]
  assign metaArb_io_in_1_bits_addr_lo = {metaArb_io_in_1_bits_idx, 6'h0}; // @[DCache.scala 425:98]
  assign new_meta_coh_state = s2_meta_error ? 2'h0 : s2_meta_corrected_3_coh_state; // @[DCache.scala 428:40]
  assign metaArb_io_in_2_bits_addr_lo = s2_vaddr[11:0]; // @[DCache.scala 437:80]
  assign metaArb_io_in_2_bits_data_meta_tag = s2_req_addr[31:12]; // @[HellaCache.scala 289:20 HellaCache.scala 290:14]
  assign _lrscBackingOff_T = lrscCount > 7'h0; // @[DCache.scala 445:34]
  assign lrscBackingOff = _lrscBackingOff_T & ~lrscValid; // @[DCache.scala 445:38]
  assign lrscAddrMatch = lrscAddr == s2_req_addr[39:6]; // @[DCache.scala 447:32]
  assign _s2_sc_fail_T = lrscValid & lrscAddrMatch; // @[DCache.scala 448:41]
  assign s2_sc_fail = _s2_write_T_3 & ~_s2_sc_fail_T; // @[DCache.scala 448:26]
  assign _T_243 = s2_valid_hit_pre_data_ecc_and_waw & _c_cat_T_47; // @[DCache.scala 449:23]
  assign _T_245 = _T_243 & ~cached_grant_wait; // @[DCache.scala 449:32]
  assign _T_246 = _T_245 | s2_valid_cached_miss; // @[DCache.scala 449:54]
  assign _lrscCount_T_2 = lrscCount - 7'h1; // @[DCache.scala 453:49]
  assign _T_250 = s2_valid_masked & lrscValid; // @[DCache.scala 454:29]
  assign _pstore1_cmd_T = s1_valid_not_nacked & s1_write; // @[DCache.scala 463:63]
  assign _pstore1_rmw_T_49 = s1_write & _s1_write_T_1; // @[DCache.scala 1159:23]
  assign _pstore1_rmw_T_50 = s1_read | _pstore1_rmw_T_49; // @[DCache.scala 1158:21]
  assign _pstore1_merge_T = s2_valid_hit_pre_data_ecc_and_waw & s2_write; // @[DCache.scala 461:46]
  assign _pstore1_merge_T_2 = _pstore1_merge_T & ~s2_sc_fail; // @[DCache.scala 461:58]
  assign pstore_drain_opportunistic = ~_dataArb_io_in_3_valid_T_56; // @[DCache.scala 473:36]
  assign pstore_drain_on_miss = releaseInFlight | pstore_drain_on_miss_REG; // @[DCache.scala 474:46]
  assign pstore1_valid = _pstore1_merge_T_2 | pstore1_held; // @[DCache.scala 478:38]
  assign _pstore_drain_structural_T = pstore1_valid_likely & pstore2_valid; // @[DCache.scala 480:54]
  assign _pstore_drain_structural_T_1 = s1_valid & s1_write; // @[DCache.scala 480:85]
  assign _pstore_drain_structural_T_2 = _pstore_drain_structural_T_1 | pstore1_rmw_r; // @[DCache.scala 480:98]
  assign pstore_drain_structural = _pstore_drain_structural_T & _pstore_drain_structural_T_2; // @[DCache.scala 480:71]
  assign _T_254 = _pstore1_merge_T | pstore1_held; // @[DCache.scala 477:96]
  assign _T_255 = _T_254 == pstore1_valid; // @[DCache.scala 481:63]
  assign _T_256 = pstore1_rmw_r | _T_255; // @[DCache.scala 481:22]
  assign _T_258 = _T_256 | reset; // @[DCache.scala 481:9]
  assign _pstore_drain_T_7 = _T_254 & ~pstore1_rmw_r; // @[DCache.scala 489:41]
  assign _pstore_drain_T_8 = _pstore_drain_T_7 | pstore2_valid; // @[DCache.scala 489:58]
  assign _pstore_drain_T_9 = pstore_drain_opportunistic | pstore_drain_on_miss; // @[DCache.scala 489:107]
  assign _pstore_drain_T_10 = _pstore_drain_T_8 & _pstore_drain_T_9; // @[DCache.scala 489:76]
  assign pstore_drain = pstore_drain_structural | _pstore_drain_T_10; // @[DCache.scala 488:48]
  assign _pstore1_held_T_8 = pstore1_valid & pstore2_valid; // @[DCache.scala 492:71]
  assign _pstore1_held_T_10 = _pstore1_held_T_8 & ~pstore_drain; // @[DCache.scala 492:88]
  assign _advance_pstore1_T_1 = pstore2_valid == pstore_drain; // @[DCache.scala 493:79]
  assign advance_pstore1 = pstore1_valid & _advance_pstore1_T_1; // @[DCache.scala 493:61]
  assign _pstore2_valid_T_1 = pstore2_valid & ~pstore_drain; // @[DCache.scala 494:34]
  assign _pstore2_valid_T_2 = _pstore2_valid_T_1 | advance_pstore1; // @[DCache.scala 494:51]
  assign pstore1_storegen_data = amoalu_io_out; // @[DCache.scala 957:27]
  assign pstore2_storegen_data = {pstore2_storegen_data_hi_hi_hi,pstore2_storegen_data_hi_hi_lo,pstore2_storegen_data_hi_lo_hi,pstore2_storegen_data_hi_lo_lo,pstore2_storegen_data_lo_hi_hi,pstore2_storegen_data_lo_hi_lo,pstore2_storegen_data_lo_lo_hi,pstore2_storegen_data_lo_lo_lo}; // @[Cat.scala 30:58]
  assign _dataArb_io_in_0_bits_addr_T = pstore2_valid ? pstore2_addr : pstore1_addr; // @[DCache.scala 520:36]
  assign _dataArb_io_in_0_bits_wdata_T = pstore2_valid ? pstore2_storegen_data : pstore1_data; // @[DCache.scala 522:63]
  assign dataArb_io_in_0_bits_wdata_lo_lo_lo = _dataArb_io_in_0_bits_wdata_T[7:0]; // @[package.scala 202:50]
  assign dataArb_io_in_0_bits_wdata_lo_lo_hi = _dataArb_io_in_0_bits_wdata_T[15:8]; // @[package.scala 202:50]
  assign dataArb_io_in_0_bits_wdata_lo_hi_lo = _dataArb_io_in_0_bits_wdata_T[23:16]; // @[package.scala 202:50]
  assign dataArb_io_in_0_bits_wdata_lo_hi_hi = _dataArb_io_in_0_bits_wdata_T[31:24]; // @[package.scala 202:50]
  assign dataArb_io_in_0_bits_wdata_hi_lo_lo = _dataArb_io_in_0_bits_wdata_T[39:32]; // @[package.scala 202:50]
  assign dataArb_io_in_0_bits_wdata_hi_lo_hi = _dataArb_io_in_0_bits_wdata_T[47:40]; // @[package.scala 202:50]
  assign dataArb_io_in_0_bits_wdata_hi_hi_lo = _dataArb_io_in_0_bits_wdata_T[55:48]; // @[package.scala 202:50]
  assign dataArb_io_in_0_bits_wdata_hi_hi_hi = _dataArb_io_in_0_bits_wdata_T[63:56]; // @[package.scala 202:50]
  assign dataArb_io_in_0_bits_wdata_lo = {dataArb_io_in_0_bits_wdata_lo_hi_hi,dataArb_io_in_0_bits_wdata_lo_hi_lo,dataArb_io_in_0_bits_wdata_lo_lo_hi,dataArb_io_in_0_bits_wdata_lo_lo_lo}; // @[Cat.scala 30:58]
  assign dataArb_io_in_0_bits_wdata_hi = {dataArb_io_in_0_bits_wdata_hi_hi_hi,dataArb_io_in_0_bits_wdata_hi_hi_lo,dataArb_io_in_0_bits_wdata_hi_lo_hi,dataArb_io_in_0_bits_wdata_hi_lo_lo}; // @[Cat.scala 30:58]
  assign _dataArb_io_in_0_bits_eccMask_T = pstore2_valid ? mask : pstore1_mask; // @[DCache.scala 528:47]
  assign dataArb_io_in_0_bits_eccMask_lo_lo_lo = |_dataArb_io_in_0_bits_eccMask_T[0]; // @[DCache.scala 1149:66]
  assign dataArb_io_in_0_bits_eccMask_lo_lo_hi = |_dataArb_io_in_0_bits_eccMask_T[1]; // @[DCache.scala 1149:66]
  assign dataArb_io_in_0_bits_eccMask_lo_hi_lo = |_dataArb_io_in_0_bits_eccMask_T[2]; // @[DCache.scala 1149:66]
  assign dataArb_io_in_0_bits_eccMask_lo_hi_hi = |_dataArb_io_in_0_bits_eccMask_T[3]; // @[DCache.scala 1149:66]
  assign dataArb_io_in_0_bits_eccMask_hi_lo_lo = |_dataArb_io_in_0_bits_eccMask_T[4]; // @[DCache.scala 1149:66]
  assign dataArb_io_in_0_bits_eccMask_hi_lo_hi = |_dataArb_io_in_0_bits_eccMask_T[5]; // @[DCache.scala 1149:66]
  assign dataArb_io_in_0_bits_eccMask_hi_hi_lo = |_dataArb_io_in_0_bits_eccMask_T[6]; // @[DCache.scala 1149:66]
  assign dataArb_io_in_0_bits_eccMask_hi_hi_hi = |_dataArb_io_in_0_bits_eccMask_T[7]; // @[DCache.scala 1149:66]
  assign dataArb_io_in_0_bits_eccMask_lo = {dataArb_io_in_0_bits_eccMask_lo_hi_hi,dataArb_io_in_0_bits_eccMask_lo_hi_lo,dataArb_io_in_0_bits_eccMask_lo_lo_hi,dataArb_io_in_0_bits_eccMask_lo_lo_lo}; // @[Cat.scala 30:58]
  assign dataArb_io_in_0_bits_eccMask_hi = {dataArb_io_in_0_bits_eccMask_hi_hi_hi,dataArb_io_in_0_bits_eccMask_hi_hi_lo,dataArb_io_in_0_bits_eccMask_hi_lo_hi,dataArb_io_in_0_bits_eccMask_hi_lo_lo}; // @[Cat.scala 30:58]
  assign _a_source_T_1 = {~uncachedInFlight_0, 1'h0}; // @[DCache.scala 548:59]
  assign a_source = _a_source_T_1[0] ? 1'h0 : 1'h1; // @[Mux.scala 47:69]
  assign acquire_address = {s2_req_addr[39:6], 6'h0}; // @[DCache.scala 549:49]
  assign a_mask = {{15'd0}, pstore1_mask}; // @[DCache.scala 553:29]
  assign _get_a_mask_sizeOH_T = {{1'd0}, s2_req_size}; // @[Misc.scala 201:34]
  assign get_a_mask_sizeOH_shiftAmount = _get_a_mask_sizeOH_T[1:0]; // @[OneHot.scala 64:49]
  assign _get_a_mask_sizeOH_T_1 = 4'h1 << get_a_mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12]
  assign get_a_mask_sizeOH = _get_a_mask_sizeOH_T_1[2:0] | 3'h1; // @[Misc.scala 201:81]
  assign _get_a_mask_T = s2_req_size >= 2'h3; // @[Misc.scala 205:21]
  assign get_a_mask_size = get_a_mask_sizeOH[2]; // @[Misc.scala 208:26]
  assign get_a_mask_bit = s2_req_addr[2]; // @[Misc.scala 209:26]
  assign get_a_mask_nbit = ~get_a_mask_bit; // @[Misc.scala 210:20]
  assign _get_a_mask_acc_T = get_a_mask_size & get_a_mask_nbit; // @[Misc.scala 214:38]
  assign get_a_mask_acc = _get_a_mask_T | _get_a_mask_acc_T; // @[Misc.scala 214:29]
  assign _get_a_mask_acc_T_1 = get_a_mask_size & get_a_mask_bit; // @[Misc.scala 214:38]
  assign get_a_mask_acc_1 = _get_a_mask_T | _get_a_mask_acc_T_1; // @[Misc.scala 214:29]
  assign get_a_mask_size_1 = get_a_mask_sizeOH[1]; // @[Misc.scala 208:26]
  assign get_a_mask_bit_1 = s2_req_addr[1]; // @[Misc.scala 209:26]
  assign get_a_mask_nbit_1 = ~get_a_mask_bit_1; // @[Misc.scala 210:20]
  assign get_a_mask_eq_2 = get_a_mask_nbit & get_a_mask_nbit_1; // @[Misc.scala 213:27]
  assign _get_a_mask_acc_T_2 = get_a_mask_size_1 & get_a_mask_eq_2; // @[Misc.scala 214:38]
  assign get_a_mask_acc_2 = get_a_mask_acc | _get_a_mask_acc_T_2; // @[Misc.scala 214:29]
  assign get_a_mask_eq_3 = get_a_mask_nbit & get_a_mask_bit_1; // @[Misc.scala 213:27]
  assign _get_a_mask_acc_T_3 = get_a_mask_size_1 & get_a_mask_eq_3; // @[Misc.scala 214:38]
  assign get_a_mask_acc_3 = get_a_mask_acc | _get_a_mask_acc_T_3; // @[Misc.scala 214:29]
  assign get_a_mask_eq_4 = get_a_mask_bit & get_a_mask_nbit_1; // @[Misc.scala 213:27]
  assign _get_a_mask_acc_T_4 = get_a_mask_size_1 & get_a_mask_eq_4; // @[Misc.scala 214:38]
  assign get_a_mask_acc_4 = get_a_mask_acc_1 | _get_a_mask_acc_T_4; // @[Misc.scala 214:29]
  assign get_a_mask_eq_5 = get_a_mask_bit & get_a_mask_bit_1; // @[Misc.scala 213:27]
  assign _get_a_mask_acc_T_5 = get_a_mask_size_1 & get_a_mask_eq_5; // @[Misc.scala 214:38]
  assign get_a_mask_acc_5 = get_a_mask_acc_1 | _get_a_mask_acc_T_5; // @[Misc.scala 214:29]
  assign get_a_mask_size_2 = get_a_mask_sizeOH[0]; // @[Misc.scala 208:26]
  assign get_a_mask_bit_2 = s2_req_addr[0]; // @[Misc.scala 209:26]
  assign get_a_mask_nbit_2 = ~get_a_mask_bit_2; // @[Misc.scala 210:20]
  assign get_a_mask_eq_6 = get_a_mask_eq_2 & get_a_mask_nbit_2; // @[Misc.scala 213:27]
  assign _get_a_mask_acc_T_6 = get_a_mask_size_2 & get_a_mask_eq_6; // @[Misc.scala 214:38]
  assign get_a_mask_lo_lo_lo = get_a_mask_acc_2 | _get_a_mask_acc_T_6; // @[Misc.scala 214:29]
  assign get_a_mask_eq_7 = get_a_mask_eq_2 & get_a_mask_bit_2; // @[Misc.scala 213:27]
  assign _get_a_mask_acc_T_7 = get_a_mask_size_2 & get_a_mask_eq_7; // @[Misc.scala 214:38]
  assign get_a_mask_lo_lo_hi = get_a_mask_acc_2 | _get_a_mask_acc_T_7; // @[Misc.scala 214:29]
  assign get_a_mask_eq_8 = get_a_mask_eq_3 & get_a_mask_nbit_2; // @[Misc.scala 213:27]
  assign _get_a_mask_acc_T_8 = get_a_mask_size_2 & get_a_mask_eq_8; // @[Misc.scala 214:38]
  assign get_a_mask_lo_hi_lo = get_a_mask_acc_3 | _get_a_mask_acc_T_8; // @[Misc.scala 214:29]
  assign get_a_mask_eq_9 = get_a_mask_eq_3 & get_a_mask_bit_2; // @[Misc.scala 213:27]
  assign _get_a_mask_acc_T_9 = get_a_mask_size_2 & get_a_mask_eq_9; // @[Misc.scala 214:38]
  assign get_a_mask_lo_hi_hi = get_a_mask_acc_3 | _get_a_mask_acc_T_9; // @[Misc.scala 214:29]
  assign get_a_mask_eq_10 = get_a_mask_eq_4 & get_a_mask_nbit_2; // @[Misc.scala 213:27]
  assign _get_a_mask_acc_T_10 = get_a_mask_size_2 & get_a_mask_eq_10; // @[Misc.scala 214:38]
  assign get_a_mask_hi_lo_lo = get_a_mask_acc_4 | _get_a_mask_acc_T_10; // @[Misc.scala 214:29]
  assign get_a_mask_eq_11 = get_a_mask_eq_4 & get_a_mask_bit_2; // @[Misc.scala 213:27]
  assign _get_a_mask_acc_T_11 = get_a_mask_size_2 & get_a_mask_eq_11; // @[Misc.scala 214:38]
  assign get_a_mask_hi_lo_hi = get_a_mask_acc_4 | _get_a_mask_acc_T_11; // @[Misc.scala 214:29]
  assign get_a_mask_eq_12 = get_a_mask_eq_5 & get_a_mask_nbit_2; // @[Misc.scala 213:27]
  assign _get_a_mask_acc_T_12 = get_a_mask_size_2 & get_a_mask_eq_12; // @[Misc.scala 214:38]
  assign get_a_mask_hi_hi_lo = get_a_mask_acc_5 | _get_a_mask_acc_T_12; // @[Misc.scala 214:29]
  assign get_a_mask_eq_13 = get_a_mask_eq_5 & get_a_mask_bit_2; // @[Misc.scala 213:27]
  assign _get_a_mask_acc_T_13 = get_a_mask_size_2 & get_a_mask_eq_13; // @[Misc.scala 214:38]
  assign get_a_mask_hi_hi_hi = get_a_mask_acc_5 | _get_a_mask_acc_T_13; // @[Misc.scala 214:29]
  assign get_mask = {get_a_mask_hi_hi_hi,get_a_mask_hi_hi_lo,get_a_mask_hi_lo_hi,get_a_mask_hi_lo_lo,get_a_mask_lo_hi_hi,get_a_mask_lo_hi_lo,get_a_mask_lo_lo_hi,get_a_mask_lo_lo_lo}; // @[Cat.scala 30:58]
  assign _atomics_T = 5'h4 == s2_req_cmd; // @[Mux.scala 80:60]
  assign _atomics_T_1_opcode = _atomics_T ? 3'h3 : 3'h0; // @[Mux.scala 80:57]
  assign atomics_a_size = {{2'd0}, s2_req_size}; // @[Edges.scala 513:17 Edges.scala 516:15]
  assign _atomics_T_1_size = _atomics_T ? atomics_a_size : 4'h0; // @[Mux.scala 80:57]
  assign _atomics_T_1_source = _atomics_T & a_source; // @[Mux.scala 80:57]
  assign atomics_a_address = s2_req_addr[31:0]; // @[Edges.scala 513:17 Edges.scala 518:15]
  assign _atomics_T_1_address = _atomics_T ? atomics_a_address : 32'h0; // @[Mux.scala 80:57]
  assign _atomics_T_1_mask = _atomics_T ? get_mask : 8'h0; // @[Mux.scala 80:57]
  assign _atomics_T_1_data = _atomics_T ? pstore1_data : 64'h0; // @[Mux.scala 80:57]
  assign _atomics_T_2 = 5'h9 == s2_req_cmd; // @[Mux.scala 80:60]
  assign _atomics_T_3_opcode = _atomics_T_2 ? 3'h3 : _atomics_T_1_opcode; // @[Mux.scala 80:57]
  assign _atomics_T_3_param = _atomics_T_2 ? 3'h0 : _atomics_T_1_opcode; // @[Mux.scala 80:57]
  assign _atomics_T_3_size = _atomics_T_2 ? atomics_a_size : _atomics_T_1_size; // @[Mux.scala 80:57]
  assign _atomics_T_3_source = _atomics_T_2 ? a_source : _atomics_T_1_source; // @[Mux.scala 80:57]
  assign _atomics_T_3_address = _atomics_T_2 ? atomics_a_address : _atomics_T_1_address; // @[Mux.scala 80:57]
  assign _atomics_T_3_mask = _atomics_T_2 ? get_mask : _atomics_T_1_mask; // @[Mux.scala 80:57]
  assign _atomics_T_3_data = _atomics_T_2 ? pstore1_data : _atomics_T_1_data; // @[Mux.scala 80:57]
  assign _atomics_T_4 = 5'ha == s2_req_cmd; // @[Mux.scala 80:60]
  assign _atomics_T_5_opcode = _atomics_T_4 ? 3'h3 : _atomics_T_3_opcode; // @[Mux.scala 80:57]
  assign _atomics_T_5_param = _atomics_T_4 ? 3'h1 : _atomics_T_3_param; // @[Mux.scala 80:57]
  assign _atomics_T_5_size = _atomics_T_4 ? atomics_a_size : _atomics_T_3_size; // @[Mux.scala 80:57]
  assign _atomics_T_5_source = _atomics_T_4 ? a_source : _atomics_T_3_source; // @[Mux.scala 80:57]
  assign _atomics_T_5_address = _atomics_T_4 ? atomics_a_address : _atomics_T_3_address; // @[Mux.scala 80:57]
  assign _atomics_T_5_mask = _atomics_T_4 ? get_mask : _atomics_T_3_mask; // @[Mux.scala 80:57]
  assign _atomics_T_5_data = _atomics_T_4 ? pstore1_data : _atomics_T_3_data; // @[Mux.scala 80:57]
  assign _atomics_T_6 = 5'hb == s2_req_cmd; // @[Mux.scala 80:60]
  assign _atomics_T_7_opcode = _atomics_T_6 ? 3'h3 : _atomics_T_5_opcode; // @[Mux.scala 80:57]
  assign _atomics_T_7_param = _atomics_T_6 ? 3'h2 : _atomics_T_5_param; // @[Mux.scala 80:57]
  assign _atomics_T_7_size = _atomics_T_6 ? atomics_a_size : _atomics_T_5_size; // @[Mux.scala 80:57]
  assign _atomics_T_7_source = _atomics_T_6 ? a_source : _atomics_T_5_source; // @[Mux.scala 80:57]
  assign _atomics_T_7_address = _atomics_T_6 ? atomics_a_address : _atomics_T_5_address; // @[Mux.scala 80:57]
  assign _atomics_T_7_mask = _atomics_T_6 ? get_mask : _atomics_T_5_mask; // @[Mux.scala 80:57]
  assign _atomics_T_7_data = _atomics_T_6 ? pstore1_data : _atomics_T_5_data; // @[Mux.scala 80:57]
  assign _atomics_T_8 = 5'h8 == s2_req_cmd; // @[Mux.scala 80:60]
  assign _atomics_T_9_opcode = _atomics_T_8 ? 3'h2 : _atomics_T_7_opcode; // @[Mux.scala 80:57]
  assign _atomics_T_9_param = _atomics_T_8 ? 3'h4 : _atomics_T_7_param; // @[Mux.scala 80:57]
  assign _atomics_T_9_size = _atomics_T_8 ? atomics_a_size : _atomics_T_7_size; // @[Mux.scala 80:57]
  assign _atomics_T_9_source = _atomics_T_8 ? a_source : _atomics_T_7_source; // @[Mux.scala 80:57]
  assign _atomics_T_9_address = _atomics_T_8 ? atomics_a_address : _atomics_T_7_address; // @[Mux.scala 80:57]
  assign _atomics_T_9_mask = _atomics_T_8 ? get_mask : _atomics_T_7_mask; // @[Mux.scala 80:57]
  assign _atomics_T_9_data = _atomics_T_8 ? pstore1_data : _atomics_T_7_data; // @[Mux.scala 80:57]
  assign _atomics_T_10 = 5'hc == s2_req_cmd; // @[Mux.scala 80:60]
  assign _atomics_T_11_opcode = _atomics_T_10 ? 3'h2 : _atomics_T_9_opcode; // @[Mux.scala 80:57]
  assign _atomics_T_11_param = _atomics_T_10 ? 3'h0 : _atomics_T_9_param; // @[Mux.scala 80:57]
  assign _atomics_T_11_size = _atomics_T_10 ? atomics_a_size : _atomics_T_9_size; // @[Mux.scala 80:57]
  assign _atomics_T_11_source = _atomics_T_10 ? a_source : _atomics_T_9_source; // @[Mux.scala 80:57]
  assign _atomics_T_11_address = _atomics_T_10 ? atomics_a_address : _atomics_T_9_address; // @[Mux.scala 80:57]
  assign _atomics_T_11_mask = _atomics_T_10 ? get_mask : _atomics_T_9_mask; // @[Mux.scala 80:57]
  assign _atomics_T_11_data = _atomics_T_10 ? pstore1_data : _atomics_T_9_data; // @[Mux.scala 80:57]
  assign _atomics_T_12 = 5'hd == s2_req_cmd; // @[Mux.scala 80:60]
  assign _atomics_T_13_opcode = _atomics_T_12 ? 3'h2 : _atomics_T_11_opcode; // @[Mux.scala 80:57]
  assign _atomics_T_13_param = _atomics_T_12 ? 3'h1 : _atomics_T_11_param; // @[Mux.scala 80:57]
  assign _atomics_T_13_size = _atomics_T_12 ? atomics_a_size : _atomics_T_11_size; // @[Mux.scala 80:57]
  assign _atomics_T_13_source = _atomics_T_12 ? a_source : _atomics_T_11_source; // @[Mux.scala 80:57]
  assign _atomics_T_13_address = _atomics_T_12 ? atomics_a_address : _atomics_T_11_address; // @[Mux.scala 80:57]
  assign _atomics_T_13_mask = _atomics_T_12 ? get_mask : _atomics_T_11_mask; // @[Mux.scala 80:57]
  assign _atomics_T_13_data = _atomics_T_12 ? pstore1_data : _atomics_T_11_data; // @[Mux.scala 80:57]
  assign _atomics_T_14 = 5'he == s2_req_cmd; // @[Mux.scala 80:60]
  assign _atomics_T_15_opcode = _atomics_T_14 ? 3'h2 : _atomics_T_13_opcode; // @[Mux.scala 80:57]
  assign _atomics_T_15_param = _atomics_T_14 ? 3'h2 : _atomics_T_13_param; // @[Mux.scala 80:57]
  assign _atomics_T_15_size = _atomics_T_14 ? atomics_a_size : _atomics_T_13_size; // @[Mux.scala 80:57]
  assign _atomics_T_15_source = _atomics_T_14 ? a_source : _atomics_T_13_source; // @[Mux.scala 80:57]
  assign _atomics_T_15_address = _atomics_T_14 ? atomics_a_address : _atomics_T_13_address; // @[Mux.scala 80:57]
  assign _atomics_T_15_mask = _atomics_T_14 ? get_mask : _atomics_T_13_mask; // @[Mux.scala 80:57]
  assign _atomics_T_15_data = _atomics_T_14 ? pstore1_data : _atomics_T_13_data; // @[Mux.scala 80:57]
  assign _atomics_T_16 = 5'hf == s2_req_cmd; // @[Mux.scala 80:60]
  assign atomics_opcode = _atomics_T_16 ? 3'h2 : _atomics_T_15_opcode; // @[Mux.scala 80:57]
  assign atomics_param = _atomics_T_16 ? 3'h3 : _atomics_T_15_param; // @[Mux.scala 80:57]
  assign atomics_size = _atomics_T_16 ? atomics_a_size : _atomics_T_15_size; // @[Mux.scala 80:57]
  assign atomics_source = _atomics_T_16 ? a_source : _atomics_T_15_source; // @[Mux.scala 80:57]
  assign atomics_address = _atomics_T_16 ? atomics_a_address : _atomics_T_15_address; // @[Mux.scala 80:57]
  assign atomics_mask = _atomics_T_16 ? get_mask : _atomics_T_15_mask; // @[Mux.scala 80:57]
  assign atomics_data = _atomics_T_16 ? pstore1_data : _atomics_T_15_data; // @[Mux.scala 80:57]
  assign _GEN_356 = {{8'd0}, release_ack_addr}; // @[DCache.scala 577:43]
  assign _tl_out_a_valid_T_1 = s2_req_addr ^ _GEN_356; // @[DCache.scala 577:43]
  assign _tl_out_a_valid_T_3 = _tl_out_a_valid_T_1[20:6] == 15'h0; // @[DCache.scala 577:118]
  assign _tl_out_a_valid_T_4 = release_ack_wait & _tl_out_a_valid_T_3; // @[DCache.scala 577:27]
  assign _tl_out_a_valid_T_6 = s2_valid_cached_miss & ~_tl_out_a_valid_T_4; // @[DCache.scala 576:29]
  assign _tl_out_a_valid_T_12 = _tl_out_a_valid_T_6 & ~s2_victim_dirty; // @[DCache.scala 577:125]
  assign tl_out_a_valid = s2_valid_uncached_pending | _tl_out_a_valid_T_12; // @[DCache.scala 575:32]
  assign _tl_out_a_bits_T_6_opcode = s2_read ? atomics_opcode : 3'h0; // @[DCache.scala 582:8]
  assign _tl_out_a_bits_T_6_param = s2_read ? atomics_param : 3'h0; // @[DCache.scala 582:8]
  assign _tl_out_a_bits_T_6_size = s2_read ? atomics_size : atomics_a_size; // @[DCache.scala 582:8]
  assign _tl_out_a_bits_T_6_source = s2_read ? atomics_source : a_source; // @[DCache.scala 582:8]
  assign _tl_out_a_bits_T_6_address = s2_read ? atomics_address : atomics_a_address; // @[DCache.scala 582:8]
  assign _tl_out_a_bits_T_6_mask = s2_read ? atomics_mask : get_mask; // @[DCache.scala 582:8]
  assign _tl_out_a_bits_T_6_data = s2_read ? atomics_data : pstore1_data; // @[DCache.scala 582:8]
  assign _tl_out_a_bits_T_7_opcode = _s2_write_T_1 ? 3'h1 : _tl_out_a_bits_T_6_opcode; // @[DCache.scala 581:8]
  assign _tl_out_a_bits_T_7_param = _s2_write_T_1 ? 3'h0 : _tl_out_a_bits_T_6_param; // @[DCache.scala 581:8]
  assign _tl_out_a_bits_T_7_size = _s2_write_T_1 ? atomics_a_size : _tl_out_a_bits_T_6_size; // @[DCache.scala 581:8]
  assign _tl_out_a_bits_T_7_source = _s2_write_T_1 ? a_source : _tl_out_a_bits_T_6_source; // @[DCache.scala 581:8]
  assign _tl_out_a_bits_T_7_address = _s2_write_T_1 ? atomics_a_address : _tl_out_a_bits_T_6_address; // @[DCache.scala 581:8]
  assign putpartial_mask = a_mask[7:0]; // @[Edges.scala 483:17 Edges.scala 489:15]
  assign _tl_out_a_bits_T_7_mask = _s2_write_T_1 ? putpartial_mask : _tl_out_a_bits_T_6_mask; // @[DCache.scala 581:8]
  assign _tl_out_a_bits_T_7_data = _s2_write_T_1 ? pstore1_data : _tl_out_a_bits_T_6_data; // @[DCache.scala 581:8]
  assign _tl_out_a_bits_T_8_opcode = s2_write ? _tl_out_a_bits_T_7_opcode : 3'h4; // @[DCache.scala 580:8]
  assign _tl_out_a_bits_T_8_param = s2_write ? _tl_out_a_bits_T_7_param : 3'h0; // @[DCache.scala 580:8]
  assign _tl_out_a_bits_T_8_size = s2_write ? _tl_out_a_bits_T_7_size : atomics_a_size; // @[DCache.scala 580:8]
  assign _tl_out_a_bits_T_8_source = s2_write ? _tl_out_a_bits_T_7_source : a_source; // @[DCache.scala 580:8]
  assign _tl_out_a_bits_T_8_address = s2_write ? _tl_out_a_bits_T_7_address : atomics_a_address; // @[DCache.scala 580:8]
  assign _tl_out_a_bits_T_8_mask = s2_write ? _tl_out_a_bits_T_7_mask : get_mask; // @[DCache.scala 580:8]
  assign _tl_out_a_bits_T_8_data = s2_write ? _tl_out_a_bits_T_7_data : 64'h0; // @[DCache.scala 580:8]
  assign tl_out_a_bits_a_param = {{1'd0}, s2_grow_param}; // @[Edges.scala 345:17 Edges.scala 347:15]
  assign tl_out_a_bits_a_address = acquire_address[31:0]; // @[Edges.scala 345:17 Edges.scala 350:15]
  assign _a_sel_T = 2'h1 << a_source; // @[OneHot.scala 65:12]
  assign a_sel = _a_sel_T[1]; // @[DCache.scala 601:66]
  assign _T_263 = auto_out_a_ready & tl_out_a_valid; // @[Decoupled.scala 40:37]
  assign _GEN_142 = a_sel | uncachedInFlight_0; // @[DCache.scala 605:18]
  assign _beats1_decode_T_1 = 27'hfff << auto_out_d_bits_size; // @[package.scala 234:77]
  assign beats1_decode = ~_beats1_decode_T_1[11:3]; // @[Edges.scala 219:59]
  assign beats1_opdata = auto_out_d_bits_opcode[0]; // @[Edges.scala 105:36]
  assign beats1 = beats1_opdata ? beats1_decode : 9'h0; // @[Edges.scala 220:14]
  assign counter1 = counter - 9'h1; // @[Edges.scala 229:28]
  assign _last_T = counter == 9'h1; // @[Edges.scala 231:25]
  assign _last_T_1 = beats1 == 9'h0; // @[Edges.scala 231:47]
  assign d_last = _last_T | _last_T_1; // @[Edges.scala 231:37]
  assign d_done = d_last & _T_271; // @[Edges.scala 232:22]
  assign count = beats1 & ~counter1; // @[Edges.scala 233:25]
  assign d_address_inc = {count, 3'h0}; // @[Edges.scala 268:29]
  assign grantIsVoluntary = auto_out_d_bits_opcode == 3'h6; // @[DCache.scala 636:32]
  assign _blockProbeAfterGrantCount_T_1 = blockProbeAfterGrantCount - 3'h1; // @[DCache.scala 640:97]
  assign _uncachedRespIdxOH_T = 2'h1 << auto_out_d_bits_source; // @[OneHot.scala 65:12]
  assign uncachedRespIdxOH = _uncachedRespIdxOH_T[1]; // @[DCache.scala 643:90]
  assign _T_273 = cached_grant_wait | reset; // @[DCache.scala 648:13]
  assign _T_276 = uncachedRespIdxOH & d_last; // @[DCache.scala 657:17]
  assign _T_278 = uncachedInFlight_0 | reset; // @[DCache.scala 658:17]
  assign dontCareBits = {s1_paddr[31:3], 3'h0}; // @[DCache.scala 672:55]
  assign _GEN_357 = {{29'd0}, uncachedReqs_0_addr[2:0]}; // @[DCache.scala 673:26]
  assign _s2_req_addr_T_1 = dontCareBits | _GEN_357; // @[DCache.scala 673:26]
  assign _T_281 = release_ack_wait | reset; // @[DCache.scala 679:13]
  assign _GEN_196 = grantIsVoluntary ? 1'h0 : release_ack_wait; // @[DCache.scala 678:36]
  assign _GEN_205 = grantIsUncached ? release_ack_wait : _GEN_196; // @[DCache.scala 655:35]
  assign _GEN_209 = grantIsCached & d_last; // @[DCache.scala 646:26]
  assign _GEN_218 = grantIsCached ? release_ack_wait : _GEN_205; // @[DCache.scala 646:26]
  assign _GEN_231 = _T_271 ? _GEN_218 : release_ack_wait; // @[DCache.scala 645:26]
  assign _bundleOut_0_e_valid_T = auto_out_d_valid & d_first; // @[DCache.scala 685:36]
  assign _bundleOut_0_e_valid_T_1 = _bundleOut_0_e_valid_T & grantIsCached; // @[DCache.scala 685:47]
  assign _bundleOut_0_e_valid_T_2 = _bundleOut_0_e_valid_T_1 & canAcceptCachedGrant; // @[DCache.scala 685:64]
  assign tl_out__e_valid = _T_292 ? 1'h0 : _bundleOut_0_e_valid_T_2; // @[DCache.scala 693:51]
  assign _T_283 = auto_out_e_ready & tl_out__e_valid; // @[Decoupled.scala 40:37]
  assign _T_285 = _T_271 & d_first; // @[DCache.scala 687:47]
  assign _T_286 = _T_285 & grantIsCached; // @[DCache.scala 687:58]
  assign _T_287 = _T_283 == _T_286; // @[DCache.scala 687:26]
  assign _T_289 = _T_287 | reset; // @[DCache.scala 687:9]
  assign _dataArb_io_in_1_valid_T = auto_out_d_valid & grantIsRefill; // @[DCache.scala 692:44]
  assign _dataArb_io_in_1_valid_T_1 = _dataArb_io_in_1_valid_T & canAcceptCachedGrant; // @[DCache.scala 692:61]
  assign _dataArb_io_in_1_bits_addr_T_1 = {s2_vaddr[39:6], 6'h0}; // @[DCache.scala 699:57]
  assign _GEN_358 = {{28'd0}, d_address_inc}; // @[DCache.scala 699:67]
  assign _dataArb_io_in_1_bits_addr_T_2 = _dataArb_io_in_1_bits_addr_T_1 | _GEN_358; // @[DCache.scala 699:67]
  assign _metaArb_io_in_3_valid_T = grantIsCached & d_done; // @[DCache.scala 712:43]
  assign _metaArb_io_in_3_bits_data_T_1 = {s2_write,c_cat_lo,auto_out_d_bits_param}; // @[Cat.scala 30:58]
  assign _metaArb_io_in_3_bits_data_T_6 = 4'h1 == _metaArb_io_in_3_bits_data_T_1; // @[Mux.scala 80:60]
  assign _metaArb_io_in_3_bits_data_T_7 = _metaArb_io_in_3_bits_data_T_6 ? 2'h1 : 2'h0; // @[Mux.scala 80:57]
  assign _metaArb_io_in_3_bits_data_T_8 = 4'h0 == _metaArb_io_in_3_bits_data_T_1; // @[Mux.scala 80:60]
  assign _metaArb_io_in_3_bits_data_T_9 = _metaArb_io_in_3_bits_data_T_8 ? 2'h2 : _metaArb_io_in_3_bits_data_T_7; // @[Mux.scala 80:57]
  assign _metaArb_io_in_3_bits_data_T_10 = 4'h4 == _metaArb_io_in_3_bits_data_T_1; // @[Mux.scala 80:60]
  assign _metaArb_io_in_3_bits_data_T_11 = _metaArb_io_in_3_bits_data_T_10 ? 2'h2 : _metaArb_io_in_3_bits_data_T_9; // @[Mux.scala 80:57]
  assign _metaArb_io_in_3_bits_data_T_12 = 4'hc == _metaArb_io_in_3_bits_data_T_1; // @[Mux.scala 80:60]
  assign metaArb_io_in_3_bits_data_meta_state = _metaArb_io_in_3_bits_data_T_12 ? 2'h3 : _metaArb_io_in_3_bits_data_T_11; // @[Mux.scala 80:57]
  assign _GEN_234 = auto_out_d_valid ? 1'h0 : _GEN_32; // @[DCache.scala 726:29]
  assign _GEN_235 = auto_out_d_valid | _dataArb_io_in_1_valid_T_1; // @[DCache.scala 726:29]
  assign _GEN_236 = auto_out_d_valid ? 1'h0 : 1'h1; // @[DCache.scala 726:29]
  assign _metaArb_io_in_6_valid_T_1 = ~block_probe_for_core_progress | lrscBackingOff; // @[DCache.scala 740:79]
  assign _metaArb_io_in_6_valid_T_2 = auto_out_b_valid & _metaArb_io_in_6_valid_T_1; // @[DCache.scala 740:44]
  assign metaArb_io_in_6_bits_addr_hi = io_cpu_req_bits_addr[39:32]; // @[DCache.scala 744:58]
  assign _metaArb_io_in_6_bits_addr_T = {metaArb_io_in_6_bits_addr_hi,auto_out_b_bits_address}; // @[Cat.scala 30:58]
  assign counter1_1 = counter_1 - 9'h1; // @[Edges.scala 229:28]
  assign c_count = beats1_1 & ~counter1_1; // @[Edges.scala 233:25]
  assign releaseRejected = s2_release_data_valid & ~_T_297; // @[DCache.scala 774:44]
  assign _releaseDataBeat_T = {1'h0,c_count}; // @[Cat.scala 30:58]
  assign _releaseDataBeat_T_1 = {1'h0,s2_release_data_valid}; // @[Cat.scala 30:58]
  assign _GEN_359 = {{1'd0}, s1_release_data_valid}; // @[DCache.scala 775:101]
  assign _releaseDataBeat_T_3 = _GEN_359 + _releaseDataBeat_T_1; // @[DCache.scala 775:101]
  assign _releaseDataBeat_T_4 = releaseRejected ? 2'h0 : _releaseDataBeat_T_3; // @[DCache.scala 775:52]
  assign _GEN_360 = {{8'd0}, _releaseDataBeat_T_4}; // @[DCache.scala 775:47]
  assign releaseDataBeat = _releaseDataBeat_T + _GEN_360; // @[DCache.scala 775:47]
  assign _T_298 = s2_valid_flush_line | s2_flush_valid; // @[DCache.scala 788:34]
  assign _T_299 = _T_298 | io_cpu_s2_nack; // @[DCache.scala 788:52]
  assign _T_301 = _T_299 | reset; // @[DCache.scala 788:13]
  assign discard_line = s2_valid_flush_line & s2_req_size[1]; // @[DCache.scala 789:46]
  assign _release_state_T_1 = s2_victim_dirty & ~discard_line; // @[DCache.scala 790:44]
  assign _release_state_T_13 = _release_state_T_1 ? 4'h1 : 4'h6; // @[DCache.scala 790:27]
  assign probe_bits_lo = s2_req_addr[11:6]; // @[DCache.scala 793:76]
  assign _probe_bits_T_1 = {s2_victim_tag,probe_bits_lo}; // @[Cat.scala 30:58]
  assign res_2_address = {_probe_bits_T_1, 6'h0}; // @[DCache.scala 793:96]
  assign _GEN_244 = s2_want_victimize ? _release_state_T_13 : release_state; // @[DCache.scala 787:25]
  assign _release_state_T_14 = releaseDone ? 4'h7 : 4'h3; // @[DCache.scala 804:29]
  assign _release_state_T_15 = releaseDone ? 4'h0 : 4'h5; // @[DCache.scala 808:29]
  assign _GEN_255 = _T_303 ? s2_report_param : 3'h5; // @[DCache.scala 801:45]
  assign _GEN_261 = _T_303 ? _release_state_T_14 : _release_state_T_15; // @[DCache.scala 801:45]
  assign _GEN_263 = s2_prb_ack_data ? 4'h2 : _GEN_261; // @[DCache.scala 799:36]
  assign _GEN_266 = s2_prb_ack_data ? 3'h5 : _GEN_255; // @[DCache.scala 799:36]
  assign _GEN_273 = s2_meta_error ? 4'h4 : _GEN_263; // @[DCache.scala 797:28]
  assign _GEN_276 = s2_meta_error ? 3'h5 : _GEN_266; // @[DCache.scala 797:28]
  assign _GEN_284 = s2_probe ? _GEN_273 : _GEN_244; // @[DCache.scala 795:21]
  assign _GEN_287 = s2_probe ? _GEN_276 : 3'h5; // @[DCache.scala 795:21]
  assign _T_304 = release_state == 4'h4; // @[DCache.scala 812:25]
  assign _metaArb_io_in_6_bits_addr_T_1 = {metaArb_io_in_6_bits_addr_hi,probe_bits_address}; // @[Cat.scala 30:58]
  assign _GEN_294 = metaArb_io_in_6_ready ? 4'h0 : _GEN_284; // @[DCache.scala 816:37]
  assign _GEN_295 = metaArb_io_in_6_ready | s1_probe_x12; // @[DCache.scala 816:37]
  assign _GEN_299 = _T_304 ? _GEN_294 : _GEN_284; // @[DCache.scala 812:44]
  assign _GEN_301 = releaseDone ? 4'h0 : _GEN_299; // @[DCache.scala 823:26]
  assign _GEN_303 = _T_305 ? _GEN_301 : _GEN_299; // @[DCache.scala 821:47]
  assign _GEN_307 = _T_306 ? s2_report_param : _GEN_287; // @[DCache.scala 825:48]
  assign _GEN_316 = _T_307 ? s2_report_param : _GEN_307; // @[DCache.scala 830:48]
  assign _T_315 = _T_297 & c_first; // @[DCache.scala 850:29]
  assign _GEN_331 = _T_315 | _GEN_231; // @[DCache.scala 850:41]
  assign newCoh_state = _T_312 ? voluntaryNewCoh_state : probeNewCoh_state; // @[DCache.scala 834:102]
  assign _dataArb_io_in_2_valid_T = releaseDataBeat < 10'h8; // @[DCache.scala 871:60]
  assign _dataArb_io_in_2_bits_addr_T_1 = {probe_bits_address[11:6], 6'h0}; // @[DCache.scala 874:55]
  assign _dataArb_io_in_2_bits_addr_T_3 = {releaseDataBeat[2:0], 3'h0}; // @[DCache.scala 874:117]
  assign _GEN_363 = {{6'd0}, _dataArb_io_in_2_bits_addr_T_3}; // @[DCache.scala 874:72]
  assign _metaArb_io_in_4_valid_T_1 = release_state == 4'h7; // @[package.scala 15:47]
  assign metaArb_io_in_4_bits_addr_lo = probe_bits_address[11:0]; // @[DCache.scala 883:90]
  assign metaArb_io_in_4_bits_data_meta_tag = probe_bits_address[31:12]; // @[DCache.scala 884:78]
  assign _T_316 = metaArb_io_in_4_ready & metaArb_io_in_4_valid; // @[Decoupled.scala 40:37]
  assign _io_cpu_ordered_T_4 = s1_valid | s2_valid; // @[DCache.scala 898:57]
  assign _io_cpu_ordered_T_5 = _io_cpu_ordered_T_4 | cached_grant_wait; // @[DCache.scala 898:94]
  assign _io_cpu_ordered_T_7 = _io_cpu_ordered_T_5 | _s2_valid_cached_miss_T_2; // @[DCache.scala 898:115]
  assign _s1_xcpt_valid_T_1 = tlb_io_req_valid; // @[DCache.scala 900:40]
  assign _T_321 = ~s2_valid_hit_pre_data_ecc_and_waw | reset; // @[DCache.scala 920:11]
  assign io_cpu_resp_bits_data_shifted = get_a_mask_bit ? s2_data_corrected[63:32] : s2_data_corrected[31:0]; // @[AMOALU.scala 39:24]
  assign _io_cpu_resp_bits_data_T = s2_req_size == 2'h2; // @[AMOALU.scala 42:26]
  assign _io_cpu_resp_bits_data_T_3 = s2_req_signed & io_cpu_resp_bits_data_shifted[31]; // @[AMOALU.scala 42:76]
  assign _io_cpu_resp_bits_data_T_5 = _io_cpu_resp_bits_data_T_3 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  assign io_cpu_resp_bits_data_hi = _io_cpu_resp_bits_data_T ? _io_cpu_resp_bits_data_T_5 : s2_data_corrected[63:32]; // @[AMOALU.scala 42:20]
  assign _io_cpu_resp_bits_data_T_7 = {io_cpu_resp_bits_data_hi,io_cpu_resp_bits_data_shifted}; // @[Cat.scala 30:58]
  assign io_cpu_resp_bits_data_shifted_1 = get_a_mask_bit_1 ? _io_cpu_resp_bits_data_T_7[31:16] : _io_cpu_resp_bits_data_T_7[15:0]; // @[AMOALU.scala 39:24]
  assign _io_cpu_resp_bits_data_T_8 = s2_req_size == 2'h1; // @[AMOALU.scala 42:26]
  assign _io_cpu_resp_bits_data_T_11 = s2_req_signed & io_cpu_resp_bits_data_shifted_1[15]; // @[AMOALU.scala 42:76]
  assign _io_cpu_resp_bits_data_T_13 = _io_cpu_resp_bits_data_T_11 ? 48'hffffffffffff : 48'h0; // @[Bitwise.scala 72:12]
  assign io_cpu_resp_bits_data_hi_1 = _io_cpu_resp_bits_data_T_8 ? _io_cpu_resp_bits_data_T_13 : _io_cpu_resp_bits_data_T_7[63:16]; // @[AMOALU.scala 42:20]
  assign _io_cpu_resp_bits_data_T_15 = {io_cpu_resp_bits_data_hi_1,io_cpu_resp_bits_data_shifted_1}; // @[Cat.scala 30:58]
  assign io_cpu_resp_bits_data_shifted_2 = get_a_mask_bit_2 ? _io_cpu_resp_bits_data_T_15[15:8] : _io_cpu_resp_bits_data_T_15[7:0]; // @[AMOALU.scala 39:24]
  assign io_cpu_resp_bits_data_lo_2 = _s2_write_T_3 ? 8'h0 : io_cpu_resp_bits_data_shifted_2; // @[AMOALU.scala 41:23]
  assign _io_cpu_resp_bits_data_T_16 = s2_req_size == 2'h0; // @[AMOALU.scala 42:26]
  assign _io_cpu_resp_bits_data_T_17 = _io_cpu_resp_bits_data_T_16 | _s2_write_T_3; // @[AMOALU.scala 42:38]
  assign _io_cpu_resp_bits_data_T_19 = s2_req_signed & io_cpu_resp_bits_data_lo_2[7]; // @[AMOALU.scala 42:76]
  assign _io_cpu_resp_bits_data_T_21 = _io_cpu_resp_bits_data_T_19 ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 72:12]
  assign io_cpu_resp_bits_data_hi_2 = _io_cpu_resp_bits_data_T_17 ? _io_cpu_resp_bits_data_T_21 : _io_cpu_resp_bits_data_T_15[63:8]; // @[AMOALU.scala 42:20]
  assign _io_cpu_resp_bits_data_T_23 = {io_cpu_resp_bits_data_hi_2,io_cpu_resp_bits_data_lo_2}; // @[Cat.scala 30:58]
  assign _GEN_364 = {{63'd0}, s2_sc_fail}; // @[DCache.scala 942:41]
  assign _GEN_349 = REG | resetting; // @[DCache.scala 976:27]
  assign flushCounterNext = flushCounter + 8'h1; // @[DCache.scala 977:39]
  assign flushDone = flushCounterNext[8:6] == 3'h4; // @[DCache.scala 978:57]
  assign _s1_flush_valid_T = metaArb_io_in_5_ready & metaArb_io_in_5_valid; // @[Decoupled.scala 40:37]
  assign _s1_flush_valid_T_2 = _s1_flush_valid_T & ~s1_flush_valid; // @[DCache.scala 982:45]
  assign _s1_flush_valid_T_4 = _s1_flush_valid_T_2 & ~s2_flush_valid_pre_tag_ecc; // @[DCache.scala 982:64]
  assign _s1_flush_valid_T_6 = _s1_flush_valid_T_4 & _io_cpu_req_ready_T; // @[DCache.scala 982:95]
  assign metaArb_io_in_5_bits_addr_lo = {metaArb_io_in_5_bits_idx, 6'h0}; // @[DCache.scala 986:98]
  assign _GEN_351 = resetting ? flushCounterNext : {{1'd0}, flushCounter}; // @[DCache.scala 1019:20]
  assign io_cpu_perf_release_counter1 = io_cpu_perf_release_counter - 9'h1; // @[Edges.scala 229:28]
  assign io_cpu_perf_release_first = io_cpu_perf_release_counter == 9'h0; // @[Edges.scala 230:25]
  assign _io_cpu_perf_release_last_T = io_cpu_perf_release_counter == 9'h1; // @[Edges.scala 231:25]
  assign io_cpu_perf_release_last = _io_cpu_perf_release_last_T | _last_T_3; // @[Edges.scala 231:37]
  assign auto_out_a_valid = s2_valid_uncached_pending | _tl_out_a_valid_T_12; // @[LazyModule.scala 311:12]
  assign auto_out_a_bits_opcode = s2_uncached ? _tl_out_a_bits_T_8_opcode : 3'h6; // @[LazyModule.scala 311:12]
  assign auto_out_a_bits_param = s2_uncached ? _tl_out_a_bits_T_8_param : tl_out_a_bits_a_param; // @[LazyModule.scala 311:12]
  assign auto_out_a_bits_size = s2_uncached ? _tl_out_a_bits_T_8_size : 4'h6; // @[LazyModule.scala 311:12]
  assign auto_out_a_bits_source = s2_uncached ? _tl_out_a_bits_T_8_source : 1'h0; // @[LazyModule.scala 311:12]
  assign auto_out_a_bits_address = s2_uncached ? _tl_out_a_bits_T_8_address : tl_out_a_bits_a_address; // @[LazyModule.scala 311:12]
  assign auto_out_a_bits_mask = s2_uncached ? _tl_out_a_bits_T_8_mask : 8'hff; // @[LazyModule.scala 311:12]
  assign auto_out_a_bits_data = s2_uncached ? _tl_out_a_bits_T_8_data : 64'h0; // @[LazyModule.scala 311:12]
  assign auto_out_b_ready = metaArb_io_in_6_ready & ~_bundleOut_0_b_ready_T_2; // @[LazyModule.scala 311:12]
  assign auto_out_c_valid = _T_306 | _GEN_302; // @[LazyModule.scala 311:12]
  assign auto_out_c_bits_opcode = _T_312 ? _GEN_323 : _GEN_315; // @[LazyModule.scala 311:12]
  assign auto_out_c_bits_param = _T_312 ? s2_shrink_param : _GEN_316; // @[LazyModule.scala 311:12]
  assign auto_out_c_bits_size = _T_312 ? 4'h6 : probe_bits_size; // @[LazyModule.scala 311:12]
  assign auto_out_c_bits_source = probe_bits_source; // @[LazyModule.scala 311:12]
  assign auto_out_c_bits_address = probe_bits_address; // @[LazyModule.scala 311:12]
  assign auto_out_c_bits_data = {s2_data_corrected_hi,s2_data_corrected_lo}; // @[LazyModule.scala 311:12]
  assign auto_out_d_ready = _T_294 ? 1'h0 : _GEN_233; // @[LazyModule.scala 311:12]
  assign auto_out_e_valid = _T_292 ? 1'h0 : _bundleOut_0_e_valid_T_2; // @[LazyModule.scala 311:12]
  assign auto_out_e_bits_sink = auto_out_d_bits_sink; // @[LazyModule.scala 311:12]
  assign io_cpu_req_ready = _T_294 ? _GEN_234 : _GEN_32; // @[DCache.scala 211:20 DCache.scala 236:64 DCache.scala 245:53 DCache.scala 253:98 DCache.scala 727:26]
  assign io_cpu_s2_nack = _io_cpu_s2_nack_T_3 & ~s2_valid_hit_pre_data_ecc_and_waw; // @[DCache.scala 416:18]
  assign io_cpu_resp_valid = s2_valid_hit_pre_data_ecc_and_waw | doUncachedResp; // @[DCache.scala 917:21]
  assign io_cpu_resp_bits_tag = s2_req_tag; // @[DCache.scala 888:20]
  assign io_cpu_resp_bits_size = s2_req_size; // @[DCache.scala 888:20]
  assign io_cpu_resp_bits_data = _io_cpu_resp_bits_data_T_23 | _GEN_364; // @[DCache.scala 888:20 DCache.scala 942:25]
  assign io_cpu_resp_bits_replay = doUncachedResp; // @[DCache.scala 890:27 DCache.scala 921:29]
  assign io_cpu_resp_bits_has_data = _s2_read_T_4 | _s2_write_T_21; // @[DCache.scala 889:29]
  assign io_cpu_resp_bits_data_word_bypass = {io_cpu_resp_bits_data_hi,io_cpu_resp_bits_data_shifted}; // @[DCache.scala 943:37]
  assign io_cpu_replay_next = _T_271 & grantIsUncachedData; // @[DCache.scala 918:22]
  assign io_cpu_s2_xcpt_ma_ld = io_cpu_s2_xcpt_REG & s2_tlb_xcpt_ma_ld; // @[DCache.scala 901:18]
  assign io_cpu_s2_xcpt_ma_st = io_cpu_s2_xcpt_REG & s2_tlb_xcpt_ma_st; // @[DCache.scala 901:18]
  assign io_cpu_s2_xcpt_pf_ld = io_cpu_s2_xcpt_REG & s2_tlb_xcpt_pf_ld; // @[DCache.scala 901:18]
  assign io_cpu_s2_xcpt_pf_st = io_cpu_s2_xcpt_REG & s2_tlb_xcpt_pf_st; // @[DCache.scala 901:18]
  assign io_cpu_s2_xcpt_ae_ld = io_cpu_s2_xcpt_REG & s2_tlb_xcpt_ae_ld; // @[DCache.scala 901:18]
  assign io_cpu_s2_xcpt_ae_st = io_cpu_s2_xcpt_REG & s2_tlb_xcpt_ae_st; // @[DCache.scala 901:18]
  assign io_cpu_ordered = ~_io_cpu_ordered_T_7; // @[DCache.scala 898:18]
  assign io_cpu_perf_release = io_cpu_perf_release_last & _T_297; // @[DCache.scala 1045:23]
  assign io_cpu_perf_grant = auto_out_d_valid & d_last; // @[DCache.scala 1046:21]
  assign io_ptw_req_valid = tlb_io_ptw_req_valid; // @[DCache.scala 249:10]
  assign io_ptw_req_bits_bits_addr = tlb_io_ptw_req_bits_bits_addr; // @[DCache.scala 249:10]
  assign tlb_clock = gated_clock;
  assign tlb_reset = reset;
  assign tlb_io_req_valid = s1_valid_masked & s1_cmd_uses_tlb; // @[DCache.scala 251:20]
  assign tlb_io_req_bits_vaddr = s1_tlb_req_vaddr; // @[DCache.scala 252:19]
  assign tlb_io_req_bits_passthrough = s1_tlb_req_passthrough; // @[DCache.scala 252:19]
  assign tlb_io_req_bits_size = s1_tlb_req_size; // @[DCache.scala 252:19]
  assign tlb_io_req_bits_cmd = s1_tlb_req_cmd; // @[DCache.scala 252:19]
  assign tlb_io_sfence_valid = s1_valid_masked & s1_sfence; // @[DCache.scala 256:23]
  assign tlb_io_sfence_bits_rs1 = s1_req_size[0]; // @[DCache.scala 257:26]
  assign tlb_io_sfence_bits_rs2 = s1_req_size[1]; // @[DCache.scala 258:26]
  assign tlb_io_sfence_bits_addr = s1_req_addr[38:0]; // @[DCache.scala 260:27]
  assign tlb_io_ptw_req_ready = io_ptw_req_ready; // @[DCache.scala 249:10]
  assign tlb_io_ptw_resp_valid = io_ptw_resp_valid; // @[DCache.scala 249:10]
  assign tlb_io_ptw_resp_bits_ae = io_ptw_resp_bits_ae; // @[DCache.scala 249:10]
  assign tlb_io_ptw_resp_bits_pte_ppn = io_ptw_resp_bits_pte_ppn; // @[DCache.scala 249:10]
  assign tlb_io_ptw_resp_bits_pte_d = io_ptw_resp_bits_pte_d; // @[DCache.scala 249:10]
  assign tlb_io_ptw_resp_bits_pte_a = io_ptw_resp_bits_pte_a; // @[DCache.scala 249:10]
  assign tlb_io_ptw_resp_bits_pte_g = io_ptw_resp_bits_pte_g; // @[DCache.scala 249:10]
  assign tlb_io_ptw_resp_bits_pte_u = io_ptw_resp_bits_pte_u; // @[DCache.scala 249:10]
  assign tlb_io_ptw_resp_bits_pte_x = io_ptw_resp_bits_pte_x; // @[DCache.scala 249:10]
  assign tlb_io_ptw_resp_bits_pte_w = io_ptw_resp_bits_pte_w; // @[DCache.scala 249:10]
  assign tlb_io_ptw_resp_bits_pte_r = io_ptw_resp_bits_pte_r; // @[DCache.scala 249:10]
  assign tlb_io_ptw_resp_bits_pte_v = io_ptw_resp_bits_pte_v; // @[DCache.scala 249:10]
  assign tlb_io_ptw_resp_bits_level = io_ptw_resp_bits_level; // @[DCache.scala 249:10]
  assign tlb_io_ptw_resp_bits_homogeneous = io_ptw_resp_bits_homogeneous; // @[DCache.scala 249:10]
  assign tlb_io_ptw_ptbr_mode = io_ptw_ptbr_mode; // @[DCache.scala 249:10]
  assign tlb_io_ptw_status_debug = io_ptw_status_debug; // @[DCache.scala 249:10]
  assign tlb_io_ptw_status_dprv = io_ptw_status_dprv; // @[DCache.scala 249:10]
  assign tlb_io_ptw_status_mxr = io_ptw_status_mxr; // @[DCache.scala 249:10]
  assign tlb_io_ptw_status_sum = io_ptw_status_sum; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_0_cfg_l = io_ptw_pmp_0_cfg_l; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_0_cfg_a = io_ptw_pmp_0_cfg_a; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_0_cfg_x = io_ptw_pmp_0_cfg_x; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_0_cfg_w = io_ptw_pmp_0_cfg_w; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_0_cfg_r = io_ptw_pmp_0_cfg_r; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_0_addr = io_ptw_pmp_0_addr; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_0_mask = io_ptw_pmp_0_mask; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_1_cfg_l = io_ptw_pmp_1_cfg_l; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_1_cfg_a = io_ptw_pmp_1_cfg_a; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_1_cfg_x = io_ptw_pmp_1_cfg_x; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_1_cfg_w = io_ptw_pmp_1_cfg_w; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_1_cfg_r = io_ptw_pmp_1_cfg_r; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_1_addr = io_ptw_pmp_1_addr; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_1_mask = io_ptw_pmp_1_mask; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_2_cfg_l = io_ptw_pmp_2_cfg_l; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_2_cfg_a = io_ptw_pmp_2_cfg_a; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_2_cfg_x = io_ptw_pmp_2_cfg_x; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_2_cfg_w = io_ptw_pmp_2_cfg_w; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_2_cfg_r = io_ptw_pmp_2_cfg_r; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_2_addr = io_ptw_pmp_2_addr; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_2_mask = io_ptw_pmp_2_mask; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_3_cfg_l = io_ptw_pmp_3_cfg_l; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_3_cfg_a = io_ptw_pmp_3_cfg_a; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_3_cfg_x = io_ptw_pmp_3_cfg_x; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_3_cfg_w = io_ptw_pmp_3_cfg_w; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_3_cfg_r = io_ptw_pmp_3_cfg_r; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_3_addr = io_ptw_pmp_3_addr; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_3_mask = io_ptw_pmp_3_mask; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_4_cfg_l = io_ptw_pmp_4_cfg_l; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_4_cfg_a = io_ptw_pmp_4_cfg_a; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_4_cfg_x = io_ptw_pmp_4_cfg_x; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_4_cfg_w = io_ptw_pmp_4_cfg_w; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_4_cfg_r = io_ptw_pmp_4_cfg_r; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_4_addr = io_ptw_pmp_4_addr; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_4_mask = io_ptw_pmp_4_mask; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_5_cfg_l = io_ptw_pmp_5_cfg_l; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_5_cfg_a = io_ptw_pmp_5_cfg_a; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_5_cfg_x = io_ptw_pmp_5_cfg_x; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_5_cfg_w = io_ptw_pmp_5_cfg_w; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_5_cfg_r = io_ptw_pmp_5_cfg_r; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_5_addr = io_ptw_pmp_5_addr; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_5_mask = io_ptw_pmp_5_mask; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_6_cfg_l = io_ptw_pmp_6_cfg_l; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_6_cfg_a = io_ptw_pmp_6_cfg_a; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_6_cfg_x = io_ptw_pmp_6_cfg_x; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_6_cfg_w = io_ptw_pmp_6_cfg_w; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_6_cfg_r = io_ptw_pmp_6_cfg_r; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_6_addr = io_ptw_pmp_6_addr; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_6_mask = io_ptw_pmp_6_mask; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_7_cfg_l = io_ptw_pmp_7_cfg_l; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_7_cfg_a = io_ptw_pmp_7_cfg_a; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_7_cfg_x = io_ptw_pmp_7_cfg_x; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_7_cfg_w = io_ptw_pmp_7_cfg_w; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_7_cfg_r = io_ptw_pmp_7_cfg_r; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_7_addr = io_ptw_pmp_7_addr; // @[DCache.scala 249:10]
  assign tlb_io_ptw_pmp_7_mask = io_ptw_pmp_7_mask; // @[DCache.scala 249:10]
  assign pma_checker_clock = gated_clock;
  assign pma_checker_reset = reset;
  assign pma_checker_io_req_valid = 1'h0;
  assign pma_checker_io_req_bits_vaddr = 40'h0;
  assign pma_checker_io_req_bits_passthrough = 1'h1; // @[DCache.scala 266:39]
  assign pma_checker_io_req_bits_size = s1_req_size; // @[DCache.scala 267:27]
  assign pma_checker_io_req_bits_cmd = s1_req_cmd; // @[DCache.scala 267:27]
  assign pma_checker_io_sfence_valid = 1'h0;
  assign pma_checker_io_sfence_bits_rs1 = 1'h0;
  assign pma_checker_io_sfence_bits_rs2 = 1'h0;
  assign pma_checker_io_sfence_bits_addr = 39'h0;
  assign pma_checker_io_ptw_req_ready = 1'h0;
  assign pma_checker_io_ptw_resp_valid = 1'h0;
  assign pma_checker_io_ptw_resp_bits_ae = 1'h0;
  assign pma_checker_io_ptw_resp_bits_pte_ppn = 54'h0;
  assign pma_checker_io_ptw_resp_bits_pte_d = 1'h0;
  assign pma_checker_io_ptw_resp_bits_pte_a = 1'h0;
  assign pma_checker_io_ptw_resp_bits_pte_g = 1'h0;
  assign pma_checker_io_ptw_resp_bits_pte_u = 1'h0;
  assign pma_checker_io_ptw_resp_bits_pte_x = 1'h0;
  assign pma_checker_io_ptw_resp_bits_pte_w = 1'h0;
  assign pma_checker_io_ptw_resp_bits_pte_r = 1'h0;
  assign pma_checker_io_ptw_resp_bits_pte_v = 1'h0;
  assign pma_checker_io_ptw_resp_bits_level = 2'h0;
  assign pma_checker_io_ptw_resp_bits_homogeneous = 1'h0;
  assign pma_checker_io_ptw_ptbr_mode = 4'h0;
  assign pma_checker_io_ptw_status_debug = 1'h0;
  assign pma_checker_io_ptw_status_dprv = 2'h0;
  assign pma_checker_io_ptw_status_mxr = 1'h0;
  assign pma_checker_io_ptw_status_sum = 1'h0;
  assign pma_checker_io_ptw_pmp_0_cfg_l = 1'h0;
  assign pma_checker_io_ptw_pmp_0_cfg_a = 2'h0;
  assign pma_checker_io_ptw_pmp_0_cfg_x = 1'h0;
  assign pma_checker_io_ptw_pmp_0_cfg_w = 1'h0;
  assign pma_checker_io_ptw_pmp_0_cfg_r = 1'h0;
  assign pma_checker_io_ptw_pmp_0_addr = 30'h0;
  assign pma_checker_io_ptw_pmp_0_mask = 32'h0;
  assign pma_checker_io_ptw_pmp_1_cfg_l = 1'h0;
  assign pma_checker_io_ptw_pmp_1_cfg_a = 2'h0;
  assign pma_checker_io_ptw_pmp_1_cfg_x = 1'h0;
  assign pma_checker_io_ptw_pmp_1_cfg_w = 1'h0;
  assign pma_checker_io_ptw_pmp_1_cfg_r = 1'h0;
  assign pma_checker_io_ptw_pmp_1_addr = 30'h0;
  assign pma_checker_io_ptw_pmp_1_mask = 32'h0;
  assign pma_checker_io_ptw_pmp_2_cfg_l = 1'h0;
  assign pma_checker_io_ptw_pmp_2_cfg_a = 2'h0;
  assign pma_checker_io_ptw_pmp_2_cfg_x = 1'h0;
  assign pma_checker_io_ptw_pmp_2_cfg_w = 1'h0;
  assign pma_checker_io_ptw_pmp_2_cfg_r = 1'h0;
  assign pma_checker_io_ptw_pmp_2_addr = 30'h0;
  assign pma_checker_io_ptw_pmp_2_mask = 32'h0;
  assign pma_checker_io_ptw_pmp_3_cfg_l = 1'h0;
  assign pma_checker_io_ptw_pmp_3_cfg_a = 2'h0;
  assign pma_checker_io_ptw_pmp_3_cfg_x = 1'h0;
  assign pma_checker_io_ptw_pmp_3_cfg_w = 1'h0;
  assign pma_checker_io_ptw_pmp_3_cfg_r = 1'h0;
  assign pma_checker_io_ptw_pmp_3_addr = 30'h0;
  assign pma_checker_io_ptw_pmp_3_mask = 32'h0;
  assign pma_checker_io_ptw_pmp_4_cfg_l = 1'h0;
  assign pma_checker_io_ptw_pmp_4_cfg_a = 2'h0;
  assign pma_checker_io_ptw_pmp_4_cfg_x = 1'h0;
  assign pma_checker_io_ptw_pmp_4_cfg_w = 1'h0;
  assign pma_checker_io_ptw_pmp_4_cfg_r = 1'h0;
  assign pma_checker_io_ptw_pmp_4_addr = 30'h0;
  assign pma_checker_io_ptw_pmp_4_mask = 32'h0;
  assign pma_checker_io_ptw_pmp_5_cfg_l = 1'h0;
  assign pma_checker_io_ptw_pmp_5_cfg_a = 2'h0;
  assign pma_checker_io_ptw_pmp_5_cfg_x = 1'h0;
  assign pma_checker_io_ptw_pmp_5_cfg_w = 1'h0;
  assign pma_checker_io_ptw_pmp_5_cfg_r = 1'h0;
  assign pma_checker_io_ptw_pmp_5_addr = 30'h0;
  assign pma_checker_io_ptw_pmp_5_mask = 32'h0;
  assign pma_checker_io_ptw_pmp_6_cfg_l = 1'h0;
  assign pma_checker_io_ptw_pmp_6_cfg_a = 2'h0;
  assign pma_checker_io_ptw_pmp_6_cfg_x = 1'h0;
  assign pma_checker_io_ptw_pmp_6_cfg_w = 1'h0;
  assign pma_checker_io_ptw_pmp_6_cfg_r = 1'h0;
  assign pma_checker_io_ptw_pmp_6_addr = 30'h0;
  assign pma_checker_io_ptw_pmp_6_mask = 32'h0;
  assign pma_checker_io_ptw_pmp_7_cfg_l = 1'h0;
  assign pma_checker_io_ptw_pmp_7_cfg_a = 2'h0;
  assign pma_checker_io_ptw_pmp_7_cfg_x = 1'h0;
  assign pma_checker_io_ptw_pmp_7_cfg_w = 1'h0;
  assign pma_checker_io_ptw_pmp_7_cfg_r = 1'h0;
  assign pma_checker_io_ptw_pmp_7_addr = 30'h0;
  assign pma_checker_io_ptw_pmp_7_mask = 32'h0;
  assign lfsr_prng_clock = gated_clock;
  assign lfsr_prng_reset = reset;
  assign lfsr_prng_io_increment = _T_271 & _GEN_209; // @[PRNG.scala 85:23]
  assign metaArb_io_in_0_valid = resetting; // @[DCache.scala 1014:26]
  assign metaArb_io_in_0_bits_addr = metaArb_io_in_5_bits_addr; // @[DCache.scala 1015:25]
  assign metaArb_io_in_0_bits_idx = metaArb_io_in_5_bits_idx; // @[DCache.scala 1015:25]
  assign metaArb_io_in_1_valid = s2_meta_error & _metaArb_io_in_1_valid_T_1; // @[DCache.scala 421:26]
  assign metaArb_io_in_1_bits_addr = {dataArb_io_in_3_bits_addr_hi,metaArb_io_in_1_bits_addr_lo}; // @[DCache.scala 425:30]
  assign metaArb_io_in_1_bits_idx = s2_probe ? probe_bits_address[11:6] : s2_vaddr[11:6]; // @[DCache.scala 424:29]
  assign metaArb_io_in_1_bits_data = {new_meta_coh_state,s2_meta_corrected_3_tag}; // @[DCache.scala 426:30]
  assign metaArb_io_in_2_valid = s2_valid_hit_pre_data_ecc_and_waw & s2_update_meta; // @[DCache.scala 433:26]
  assign metaArb_io_in_2_bits_addr = {dataArb_io_in_3_bits_addr_hi,metaArb_io_in_2_bits_addr_lo}; // @[DCache.scala 437:30]
  assign metaArb_io_in_2_bits_idx = s2_vaddr[11:6]; // @[DCache.scala 436:29]
  assign metaArb_io_in_2_bits_way_en = s2_hit_valid ? s2_hit_way : s2_victim_way; // @[DCache.scala 435:32]
  assign metaArb_io_in_2_bits_data = {s2_grow_param,metaArb_io_in_2_bits_data_meta_tag}; // @[DCache.scala 438:30]
  assign metaArb_io_in_3_valid = _metaArb_io_in_3_valid_T & ~auto_out_d_bits_denied; // @[DCache.scala 712:26]
  assign metaArb_io_in_3_bits_addr = {dataArb_io_in_3_bits_addr_hi,metaArb_io_in_2_bits_addr_lo}; // @[DCache.scala 716:30]
  assign metaArb_io_in_3_bits_idx = s2_vaddr[11:6]; // @[DCache.scala 715:29]
  assign metaArb_io_in_3_bits_way_en = refill_way; // @[DCache.scala 714:32]
  assign metaArb_io_in_3_bits_data = {metaArb_io_in_3_bits_data_meta_state,metaArb_io_in_2_bits_data_meta_tag}; // @[DCache.scala 717:30]
  assign metaArb_io_in_4_valid = _T_309 | _metaArb_io_in_4_valid_T_1; // @[DCache.scala 879:26]
  assign metaArb_io_in_4_bits_addr = {dataArb_io_in_3_bits_addr_hi,metaArb_io_in_4_bits_addr_lo}; // @[DCache.scala 883:30]
  assign metaArb_io_in_4_bits_idx = probe_bits_address[11:6]; // @[DCache.scala 882:29]
  assign metaArb_io_in_4_bits_way_en = _T_312 ? s2_victim_or_hit_way : s2_probe_way; // @[DCache.scala 881:32]
  assign metaArb_io_in_4_bits_data = {newCoh_state,metaArb_io_in_4_bits_data_meta_tag}; // @[DCache.scala 884:30]
  assign metaArb_io_in_5_valid = 1'h0; // @[DCache.scala 983:26]
  assign metaArb_io_in_5_bits_addr = {dataArb_io_in_3_bits_addr_hi,metaArb_io_in_5_bits_addr_lo}; // @[DCache.scala 986:30]
  assign metaArb_io_in_5_bits_idx = flushCounter[5:0]; // @[DCache.scala 985:29]
  assign metaArb_io_in_6_valid = _T_304 | _metaArb_io_in_6_valid_T_2; // @[DCache.scala 740:26 DCache.scala 813:30]
  assign metaArb_io_in_6_bits_addr = _T_304 ? _metaArb_io_in_6_bits_addr_T_1 : _metaArb_io_in_6_bits_addr_T; // @[DCache.scala 744:30 DCache.scala 815:34]
  assign metaArb_io_in_6_bits_idx = _T_304 ? probe_bits_address[11:6] : auto_out_b_bits_address[11:6]; // @[DCache.scala 743:29 DCache.scala 814:33]
  assign metaArb_io_in_6_bits_way_en = metaArb_io_in_4_bits_way_en; // @[DCache.scala 745:32]
  assign metaArb_io_in_6_bits_data = metaArb_io_in_4_bits_data; // @[DCache.scala 746:30]
  assign metaArb_io_in_7_valid = io_cpu_req_valid; // @[DCache.scala 239:26]
  assign metaArb_io_in_7_bits_addr = io_cpu_req_bits_addr; // @[DCache.scala 242:30]
  assign metaArb_io_in_7_bits_idx = dataArb_io_in_3_bits_addr[11:6]; // @[DCache.scala 241:29]
  assign metaArb_io_in_7_bits_way_en = metaArb_io_in_4_bits_way_en; // @[DCache.scala 243:32]
  assign metaArb_io_in_7_bits_data = metaArb_io_in_4_bits_data; // @[DCache.scala 244:30]
  assign data_clock = gated_clock;
  assign data_io_req_valid = dataArb_io_out_valid; // @[DCache.scala 135:15]
  assign data_io_req_bits_addr = dataArb_io_out_bits_addr; // @[DCache.scala 135:15]
  assign data_io_req_bits_write = dataArb_io_out_bits_write; // @[DCache.scala 135:15]
  assign data_io_req_bits_wdata = dataArb_io_out_bits_wdata; // @[DCache.scala 135:15]
  assign data_io_req_bits_eccMask = dataArb_io_out_bits_eccMask; // @[DCache.scala 135:15]
  assign data_io_req_bits_way_en = dataArb_io_out_bits_way_en; // @[DCache.scala 135:15]
  assign dataArb_io_in_0_valid = pstore_drain_structural | _pstore_drain_T_10; // @[DCache.scala 518:26]
  assign dataArb_io_in_0_bits_addr = _dataArb_io_in_0_bits_addr_T[11:0]; // @[DCache.scala 520:30]
  assign dataArb_io_in_0_bits_write = pstore_drain_structural | _pstore_drain_T_10; // @[DCache.scala 519:31]
  assign dataArb_io_in_0_bits_wdata = {dataArb_io_in_0_bits_wdata_hi,dataArb_io_in_0_bits_wdata_lo}; // @[DCache.scala 522:31]
  assign dataArb_io_in_0_bits_eccMask = {dataArb_io_in_0_bits_eccMask_hi,dataArb_io_in_0_bits_eccMask_lo}; // @[DCache.scala 528:33]
  assign dataArb_io_in_0_bits_way_en = pstore2_valid ? pstore2_way : pstore1_way; // @[DCache.scala 521:32]
  assign dataArb_io_in_1_valid = _T_294 ? _GEN_235 : _dataArb_io_in_1_valid_T_1; // @[DCache.scala 692:26 DCache.scala 728:32]
  assign dataArb_io_in_1_bits_addr = _dataArb_io_in_1_bits_addr_T_2[11:0]; // @[DCache.scala 699:32]
  assign dataArb_io_in_1_bits_write = _T_294 ? _GEN_236 : 1'h1; // @[DCache.scala 698:33 DCache.scala 729:37]
  assign dataArb_io_in_1_bits_wdata = {tl_d_data_encoded_hi,tl_d_data_encoded_lo}; // @[DCache.scala 134:43 DCache.scala 701:33]
  assign dataArb_io_in_1_bits_way_en = refill_way; // @[DCache.scala 700:34]
  assign dataArb_io_in_2_valid = inWriteback & _dataArb_io_in_2_valid_T; // @[DCache.scala 871:26]
  assign dataArb_io_in_2_bits_addr = _dataArb_io_in_2_bits_addr_T_1 | _GEN_363; // @[DCache.scala 872:25 DCache.scala 874:30]
  assign dataArb_io_in_2_bits_wdata = dataArb_io_in_1_bits_wdata; // @[DCache.scala 134:43 DCache.scala 872:25]
  assign dataArb_io_in_3_valid = io_cpu_req_valid & res; // @[DCache.scala 220:26]
  assign dataArb_io_in_3_bits_addr = _dataArb_io_in_3_bits_addr_T[11:0]; // @[DCache.scala 221:25 DCache.scala 223:30]
  assign dataArb_io_in_3_bits_wdata = dataArb_io_in_1_bits_wdata; // @[DCache.scala 134:43 DCache.scala 221:25]
  assign dataArb_io_in_3_bits_wordMask = 1'h1; // @[DCache.scala 221:25 DCache.scala 224:34]
  assign amoalu_io_mask = pstore1_mask; // @[DCache.scala 951:22]
  assign amoalu_io_cmd = pstore1_cmd; // @[DCache.scala 952:21]
  assign amoalu_io_lhs = {s2_data_corrected_hi,s2_data_corrected_lo}; // @[DCache.scala 953:21]
  assign amoalu_io_rhs = pstore1_data; // @[DCache.scala 954:21]
  assign _GEN_367 = _T_271 & grantIsCached; // @[DCache.scala 648:13]
  assign _GEN_370 = _T_271 & ~grantIsCached; // @[DCache.scala 658:17]
  assign _GEN_371 = _GEN_370 & grantIsUncached; // @[DCache.scala 658:17]
  assign _GEN_372 = _GEN_371 & _T_276; // @[DCache.scala 658:17]
  assign _GEN_380 = _GEN_370 & ~grantIsUncached; // @[DCache.scala 679:13]
  assign _GEN_381 = _GEN_380 & grantIsVoluntary; // @[DCache.scala 679:13]
  assign DCache_cov_read_addr = DCache_state;
  assign DCache_cov_read_data = DCache_cov[DCache_cov_read_addr]; // @[Coverage map for DCache]
  assign DCache_cov_write_data = 1'h1;
  assign DCache_cov_write_addr = DCache_state;
  assign DCache_cov_write_mask = 1'h1;
  assign DCache_cov_write_en = 1'h1;
  assign mux_cond_0 = s1_req_addr[0];
  assign mux_cond_1 = get_a_mask_bit_2;
  assign mux_cond_2 = s1_req_addr[2];
  assign mux_cond_3 = get_a_mask_bit;
  assign mux_cond_4 = get_a_mask_bit_1;
  assign mux_cond_5 = s1_req_addr[1];
  assign s2_req_size_shl = {s2_req_size, 3'h0};
  assign s2_req_size_pad = {15'h0,s2_req_size_shl};
  assign pstore1_held_shl = {pstore1_held, 9'h0};
  assign pstore1_held_pad = {10'h0,pstore1_held_shl};
  assign s2_req_signed_shl = {s2_req_signed, 5'h0};
  assign s2_req_signed_pad = {14'h0,s2_req_signed_shl};
  assign pstore2_valid_shl = {pstore2_valid, 10'h0};
  assign pstore2_valid_pad = {9'h0,pstore2_valid_shl};
  assign s1_flush_valid_shl = {s1_flush_valid, 17'h0};
  assign s1_flush_valid_pad = {2'h0,s1_flush_valid_shl};
  assign uncachedInFlight_0_shl = {uncachedInFlight_0, 8'h0};
  assign uncachedInFlight_0_pad = {11'h0,uncachedInFlight_0_shl};
  assign blockUncachedGrant_shl = {blockUncachedGrant, 18'h0};
  assign blockUncachedGrant_pad = {1'h0,blockUncachedGrant_shl};
  assign probe_bits_param_shl = {probe_bits_param, 12'h0};
  assign probe_bits_param_pad = {6'h0,probe_bits_param_shl};
  assign s2_flush_valid_pre_tag_ecc_shl = {s2_flush_valid_pre_tag_ecc, 16'h0};
  assign s2_flush_valid_pre_tag_ecc_pad = {3'h0,s2_flush_valid_pre_tag_ecc_shl};
  assign s1_read_mask_shl = {s1_read_mask, 10'h0};
  assign s1_read_mask_pad = {9'h0,s1_read_mask_shl};
  assign s2_victim_way_r_shl = {s2_victim_way_r, 12'h0};
  assign s2_victim_way_r_pad = {6'h0,s2_victim_way_r_shl};
  assign s1_probe_shl = {s1_probe, 13'h0};
  assign s1_probe_pad = {6'h0,s1_probe_shl};
  assign release_ack_wait_shl = {release_ack_wait, 2'h0};
  assign release_ack_wait_pad = {17'h0,release_ack_wait_shl};
  assign s2_hit_state_state_shl = {s2_hit_state_state, 11'h0};
  assign s2_hit_state_state_pad = {7'h0,s2_hit_state_state_shl};
  assign cached_grant_wait_shl = {cached_grant_wait, 15'h0};
  assign cached_grant_wait_pad = {4'h0,cached_grant_wait_shl};
  assign s1_valid_shl = {s1_valid, 19'h0};
  assign s1_valid_pad = s1_valid_shl;
  assign s2_pma_cacheable_shl = {s2_pma_cacheable, 18'h0};
  assign s2_pma_cacheable_pad = {1'h0,s2_pma_cacheable_shl};
  assign s1_did_read_shl = {s1_did_read, 17'h0};
  assign s1_did_read_pad = {2'h0,s1_did_read_shl};
  assign s2_probe_shl = {s2_probe, 19'h0};
  assign s2_probe_pad = s2_probe_shl;
  assign s2_hit_way_shl = {s2_hit_way, 3'h0};
  assign s2_hit_way_pad = {13'h0,s2_hit_way_shl};
  assign s2_not_nacked_in_s1_shl = {s2_not_nacked_in_s1, 9'h0};
  assign s2_not_nacked_in_s1_pad = {10'h0,s2_not_nacked_in_s1_shl};
  assign s2_probe_state_state_shl = {s2_probe_state_state, 17'h0};
  assign s2_probe_state_state_pad = {1'h0,s2_probe_state_state_shl};
  assign s1_req_size_shl = {s1_req_size, 3'h0};
  assign s1_req_size_pad = {15'h0,s1_req_size_shl};
  assign pstore1_rmw_r_shl = {pstore1_rmw_r, 14'h0};
  assign pstore1_rmw_r_pad = {5'h0,pstore1_rmw_r_shl};
  assign s2_release_data_valid_shl = {s2_release_data_valid, 7'h0};
  assign s2_release_data_valid_pad = {12'h0,s2_release_data_valid_shl};
  assign s2_valid_shl = {s2_valid, 8'h0};
  assign s2_valid_pad = {11'h0,s2_valid_shl};
  assign pstore_drain_on_miss_REG_shl = {pstore_drain_on_miss_REG, 19'h0};
  assign pstore_drain_on_miss_REG_pad = pstore_drain_on_miss_REG_shl;
  assign resetting_shl = {resetting, 15'h0};
  assign resetting_pad = {4'h0,resetting_shl};
  assign grantInProgress_shl = {grantInProgress, 19'h0};
  assign grantInProgress_pad = grantInProgress_shl;
  assign s2_probe_way_shl = {s2_probe_way, 9'h0};
  assign s2_probe_way_pad = {7'h0,s2_probe_way_shl};
  assign mux_cond_0_shl = {mux_cond_0, 11'h0};
  assign mux_cond_0_pad = {8'h0,mux_cond_0_shl};
  assign mux_cond_1_shl = {mux_cond_1, 1'h0};
  assign mux_cond_1_pad = {18'h0,mux_cond_1_shl};
  assign mux_cond_2_shl = {mux_cond_2, 15'h0};
  assign mux_cond_2_pad = {4'h0,mux_cond_2_shl};
  assign mux_cond_3_shl = {mux_cond_3, 6'h0};
  assign mux_cond_3_pad = {13'h0,mux_cond_3_shl};
  assign mux_cond_4_shl = {mux_cond_4, 7'h0};
  assign mux_cond_4_pad = {12'h0,mux_cond_4_shl};
  assign mux_cond_5_shl = {mux_cond_5, 7'h0};
  assign mux_cond_5_pad = {12'h0,mux_cond_5_shl};
  assign DCache_xor15 = s2_req_size_pad ^ pstore1_held_pad;
  assign DCache_xor16 = s2_req_signed_pad ^ pstore2_valid_pad;
  assign DCache_xor7 = DCache_xor15 ^ DCache_xor16;
  assign DCache_xor17 = s1_flush_valid_pad ^ uncachedInFlight_0_pad;
  assign DCache_xor38 = probe_bits_param_pad ^ s2_flush_valid_pre_tag_ecc_pad;
  assign DCache_xor18 = blockUncachedGrant_pad ^ DCache_xor38;
  assign DCache_xor8 = DCache_xor17 ^ DCache_xor18;
  assign DCache_xor3 = DCache_xor7 ^ DCache_xor8;
  assign DCache_xor19 = s1_read_mask_pad ^ s2_victim_way_r_pad;
  assign DCache_xor20 = s1_probe_pad ^ release_ack_wait_pad;
  assign DCache_xor9 = DCache_xor19 ^ DCache_xor20;
  assign DCache_xor21 = s2_hit_state_state_pad ^ cached_grant_wait_pad;
  assign DCache_xor46 = s2_pma_cacheable_pad ^ s1_did_read_pad;
  assign DCache_xor22 = s1_valid_pad ^ DCache_xor46;
  assign DCache_xor10 = DCache_xor21 ^ DCache_xor22;
  assign DCache_xor4 = DCache_xor9 ^ DCache_xor10;
  assign DCache_xor1 = DCache_xor3 ^ DCache_xor4;
  assign DCache_xor23 = s2_probe_pad ^ s2_hit_way_pad;
  assign DCache_xor24 = s2_not_nacked_in_s1_pad ^ s2_probe_state_state_pad;
  assign DCache_xor11 = DCache_xor23 ^ DCache_xor24;
  assign DCache_xor25 = s1_req_size_pad ^ pstore1_rmw_r_pad;
  assign DCache_xor54 = s2_valid_pad ^ pstore_drain_on_miss_REG_pad;
  assign DCache_xor26 = s2_release_data_valid_pad ^ DCache_xor54;
  assign DCache_xor12 = DCache_xor25 ^ DCache_xor26;
  assign DCache_xor5 = DCache_xor11 ^ DCache_xor12;
  assign DCache_xor27 = resetting_pad ^ grantInProgress_pad;
  assign DCache_xor28 = s2_probe_way_pad ^ mux_cond_0_pad;
  assign DCache_xor13 = DCache_xor27 ^ DCache_xor28;
  assign DCache_xor29 = mux_cond_1_pad ^ mux_cond_2_pad;
  assign DCache_xor62 = mux_cond_4_pad ^ mux_cond_5_pad;
  assign DCache_xor30 = mux_cond_3_pad ^ DCache_xor62;
  assign DCache_xor14 = DCache_xor29 ^ DCache_xor30;
  assign DCache_xor6 = DCache_xor13 ^ DCache_xor14;
  assign DCache_xor2 = DCache_xor5 ^ DCache_xor6;
  assign DCache_xor0 = DCache_xor1 ^ DCache_xor2;
  assign data_sum = DCache_covSum + data_io_covSum;
  assign tlb_sum = data_sum + tlb_io_covSum;
  assign pma_checker_sum = tlb_sum + pma_checker_io_covSum;
  assign metaArb_sum = pma_checker_sum + metaArb_io_covSum;
  assign lfsr_prng_sum = metaArb_sum + lfsr_prng_io_covSum;
  assign amoalu_sum = lfsr_prng_sum + amoalu_io_covSum;
  assign dataArb_sum = amoalu_sum + dataArb_io_covSum;
  assign io_covSum = dataArb_sum;
  assign stopEn0 = ~_dataArb_io_in_3_valid_T_54;
  assign stopEn1 = ~_T_68;
  assign stopEn2 = ~_dataArb_io_in_3_valid_T_54;
  assign stopEn3 = ~_T_258;
  assign stopEn4 = _GEN_367 & ~_T_273;
  assign stopEn5 = _GEN_372 & ~_T_278;
  assign stopEn6 = _GEN_381 & ~_T_281;
  assign stopEn7 = ~_T_289;
  assign stopEn8 = s2_want_victimize & ~_T_301;
  assign stopEn9 = doUncachedResp & ~_T_321;
  assign lfsr_prng_metaAssert_wire = lfsr_prng_metaAssert;
  assign tlb_metaAssert_wire = tlb_metaAssert;
  assign amoalu_metaAssert_wire = amoalu_metaAssert;
  assign data_metaAssert_wire = data_metaAssert;
  assign dataArb_metaAssert_wire = dataArb_metaAssert;
  assign pma_checker_metaAssert_wire = pma_checker_metaAssert;
  assign metaArb_metaAssert_wire = metaArb_metaAssert;
  assign DCache_or7 = stopEn0 | stopEn1;
  assign DCache_or8 = stopEn2 | stopEn3;
  assign DCache_or3 = DCache_or7 | DCache_or8;
  assign DCache_or9 = stopEn4 | stopEn5;
  assign DCache_or10 = stopEn6 | stopEn7;
  assign DCache_or4 = DCache_or9 | DCache_or10;
  assign DCache_or1 = DCache_or3 | DCache_or4;
  assign DCache_or11 = stopEn8 | stopEn9;
  assign DCache_or12 = dataArb_metaAssert_wire | tlb_metaAssert_wire;
  assign DCache_or5 = DCache_or11 | DCache_or12;
  assign DCache_or13 = amoalu_metaAssert_wire | lfsr_prng_metaAssert_wire;
  assign DCache_or30 = pma_checker_metaAssert_wire | metaArb_metaAssert_wire;
  assign DCache_or14 = data_metaAssert_wire | DCache_or30;
  assign DCache_or6 = DCache_or13 | DCache_or14;
  assign DCache_or2 = DCache_or5 | DCache_or6;
  assign DCache_or0 = DCache_or1 | DCache_or2;
  assign metaAssert = DCache_or0;
  assign data_metaReset = metaReset | data_halt;
  assign tlb_metaReset = metaReset | tlb_halt;
  assign pma_checker_metaReset = metaReset | pma_checker_halt;
  assign lfsr_prng_metaReset = metaReset | lfsr_prng_halt;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tag_array_0[initvar] = _RAND_0[21:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  tag_array_0_s1_meta_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  tag_array_0_s1_meta_addr_pipe_0 = _RAND_2[5:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tag_array_1[initvar] = _RAND_3[21:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  tag_array_1_s1_meta_en_pipe_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  tag_array_1_s1_meta_addr_pipe_0 = _RAND_5[5:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tag_array_2[initvar] = _RAND_6[21:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  tag_array_2_s1_meta_en_pipe_0 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  tag_array_2_s1_meta_addr_pipe_0 = _RAND_8[5:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tag_array_3[initvar] = _RAND_9[21:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  tag_array_3_s1_meta_en_pipe_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  tag_array_3_s1_meta_addr_pipe_0 = _RAND_11[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  s1_valid = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  blockProbeAfterGrantCount = _RAND_13[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  lrscCount = _RAND_14[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  s1_probe = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  s2_probe = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  release_state = _RAND_17[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  release_ack_wait = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  release_ack_addr = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  grantInProgress = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  s2_valid = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  probe_bits_param = _RAND_22[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  probe_bits_size = _RAND_23[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  probe_bits_source = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  probe_bits_address = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  s2_probe_state_state = _RAND_26[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  counter_1 = _RAND_27[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  s2_release_data_valid = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  s1_req_cmd = _RAND_29[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  s2_req_cmd = _RAND_30[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  pstore1_held = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {2{`RANDOM}};
  pstore1_addr = _RAND_32[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {2{`RANDOM}};
  s1_req_addr = _RAND_33[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  pstore1_mask = _RAND_34[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  s1_req_size = _RAND_35[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  pstore2_valid = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {2{`RANDOM}};
  pstore2_addr = _RAND_37[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  mask = _RAND_38[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  s2_not_nacked_in_s1 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  s2_hit_state_state = _RAND_40[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  s1_req_tag = _RAND_41[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  s1_req_signed = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {2{`RANDOM}};
  s1_tlb_req_vaddr = _RAND_43[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  s1_tlb_req_passthrough = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  s1_tlb_req_size = _RAND_45[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  s1_tlb_req_cmd = _RAND_46[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  s1_flush_valid = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  cached_grant_wait = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  resetting = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  flushCounter = _RAND_50[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  refill_way = _RAND_51[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  uncachedInFlight_0 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {2{`RANDOM}};
  uncachedReqs_0_addr = _RAND_53[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  uncachedReqs_0_tag = _RAND_54[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  uncachedReqs_0_size = _RAND_55[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  uncachedReqs_0_signed = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  s1_did_read = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  s1_read_mask = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  s2_hit_way = _RAND_59[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  s2_victim_way_r = _RAND_60[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  s2_probe_way = _RAND_61[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {2{`RANDOM}};
  s2_req_addr = _RAND_62[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  s2_req_tag = _RAND_63[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  s2_req_size = _RAND_64[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  s2_req_signed = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  s2_tlb_xcpt_pf_ld = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  s2_tlb_xcpt_pf_st = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  s2_tlb_xcpt_ae_ld = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  s2_tlb_xcpt_ae_st = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  s2_tlb_xcpt_ma_ld = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  s2_tlb_xcpt_ma_st = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  s2_pma_cacheable = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {2{`RANDOM}};
  s2_vaddr_r = _RAND_73[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  s2_flush_valid_pre_tag_ecc = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  s2_meta_corrected_r = _RAND_75[21:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  s2_meta_corrected_r_1 = _RAND_76[21:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  s2_meta_corrected_r_2 = _RAND_77[21:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  s2_meta_corrected_r_3 = _RAND_78[21:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  blockUncachedGrant = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  counter = _RAND_80[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {2{`RANDOM}};
  s2_data = _RAND_81[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {2{`RANDOM}};
  lrscAddr = _RAND_82[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  pstore1_cmd = _RAND_83[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {2{`RANDOM}};
  pstore1_data = _RAND_84[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  pstore1_way = _RAND_85[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  pstore1_rmw_r = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  pstore_drain_on_miss_REG = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  pstore2_way = _RAND_88[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  pstore2_storegen_data_lo_lo_lo = _RAND_89[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  pstore2_storegen_data_lo_lo_hi = _RAND_90[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  pstore2_storegen_data_lo_hi_lo = _RAND_91[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  pstore2_storegen_data_lo_hi_hi = _RAND_92[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  pstore2_storegen_data_hi_lo_lo = _RAND_93[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  pstore2_storegen_data_hi_lo_hi = _RAND_94[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  pstore2_storegen_data_hi_hi_lo = _RAND_95[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  pstore2_storegen_data_hi_hi_hi = _RAND_96[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  s1_release_data_valid = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  io_cpu_s2_xcpt_REG = _RAND_98[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  doUncachedResp = _RAND_99[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  REG = _RAND_100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  io_cpu_perf_release_counter = _RAND_101[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  DCache_state = _RAND_102[19:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1048576; initvar = initvar+1)
    DCache_cov[initvar] = _RAND_103[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  DCache_covSum = _RAND_104[29:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge gated_clock) begin
    if(tag_array_0_MPORT_en & tag_array_0_MPORT_mask) begin
      tag_array_0[tag_array_0_MPORT_addr] <= tag_array_0_MPORT_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      tag_array_0_s1_meta_en_pipe_0 <= 1'h0;
    end else begin
      tag_array_0_s1_meta_en_pipe_0 <= metaArb_io_out_valid & ~metaArb_io_out_bits_write;
    end
    if (metaReset) begin
      tag_array_0_s1_meta_addr_pipe_0 <= 6'h0;
    end else if (metaArb_io_out_valid & ~metaArb_io_out_bits_write) begin
      tag_array_0_s1_meta_addr_pipe_0 <= metaArb_io_out_bits_idx;
    end
    if(tag_array_1_MPORT_en & tag_array_1_MPORT_mask) begin
      tag_array_1[tag_array_1_MPORT_addr] <= tag_array_1_MPORT_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      tag_array_1_s1_meta_en_pipe_0 <= 1'h0;
    end else begin
      tag_array_1_s1_meta_en_pipe_0 <= metaArb_io_out_valid & ~metaArb_io_out_bits_write;
    end
    if (metaReset) begin
      tag_array_1_s1_meta_addr_pipe_0 <= 6'h0;
    end else if (metaArb_io_out_valid & ~metaArb_io_out_bits_write) begin
      tag_array_1_s1_meta_addr_pipe_0 <= metaArb_io_out_bits_idx;
    end
    if(tag_array_2_MPORT_en & tag_array_2_MPORT_mask) begin
      tag_array_2[tag_array_2_MPORT_addr] <= tag_array_2_MPORT_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      tag_array_2_s1_meta_en_pipe_0 <= 1'h0;
    end else begin
      tag_array_2_s1_meta_en_pipe_0 <= metaArb_io_out_valid & ~metaArb_io_out_bits_write;
    end
    if (metaReset) begin
      tag_array_2_s1_meta_addr_pipe_0 <= 6'h0;
    end else if (metaArb_io_out_valid & ~metaArb_io_out_bits_write) begin
      tag_array_2_s1_meta_addr_pipe_0 <= metaArb_io_out_bits_idx;
    end
    if(tag_array_3_MPORT_en & tag_array_3_MPORT_mask) begin
      tag_array_3[tag_array_3_MPORT_addr] <= tag_array_3_MPORT_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      tag_array_3_s1_meta_en_pipe_0 <= 1'h0;
    end else begin
      tag_array_3_s1_meta_en_pipe_0 <= metaArb_io_out_valid & ~metaArb_io_out_bits_write;
    end
    if (metaReset) begin
      tag_array_3_s1_meta_addr_pipe_0 <= 6'h0;
    end else if (metaArb_io_out_valid & ~metaArb_io_out_bits_write) begin
      tag_array_3_s1_meta_addr_pipe_0 <= metaArb_io_out_bits_idx;
    end
    if (metaReset) begin
      s1_valid <= 1'h0;
    end else if (reset) begin
      s1_valid <= 1'h0;
    end else begin
      s1_valid <= s1_valid_x9;
    end
    if (metaReset) begin
      blockProbeAfterGrantCount <= 3'h0;
    end else if (reset) begin
      blockProbeAfterGrantCount <= 3'h0;
    end else if (_T_271) begin
      if (grantIsCached) begin
        if (d_last) begin
          blockProbeAfterGrantCount <= 3'h7;
        end else if (_block_probe_for_core_progress_T) begin
          blockProbeAfterGrantCount <= _blockProbeAfterGrantCount_T_1;
        end
      end else if (_block_probe_for_core_progress_T) begin
        blockProbeAfterGrantCount <= _blockProbeAfterGrantCount_T_1;
      end
    end else if (_block_probe_for_core_progress_T) begin
      blockProbeAfterGrantCount <= _blockProbeAfterGrantCount_T_1;
    end
    if (metaReset) begin
      lrscCount <= 7'h0;
    end else if (reset) begin
      lrscCount <= 7'h0;
    end else if (s1_probe) begin
      lrscCount <= 7'h0;
    end else if (_T_250) begin
      lrscCount <= 7'h3;
    end else if (_lrscBackingOff_T) begin
      lrscCount <= _lrscCount_T_2;
    end else if (_T_246) begin
      if (s2_hit) begin
        lrscCount <= 7'h4f;
      end else begin
        lrscCount <= 7'h0;
      end
    end
    if (metaReset) begin
      s1_probe <= 1'h0;
    end else if (reset) begin
      s1_probe <= 1'h0;
    end else if (_T_304) begin
      s1_probe <= _GEN_295;
    end else begin
      s1_probe <= s1_probe_x12;
    end
    if (metaReset) begin
      s2_probe <= 1'h0;
    end else if (reset) begin
      s2_probe <= 1'h0;
    end else begin
      s2_probe <= s1_probe;
    end
    if (metaReset) begin
      release_state <= 4'h0;
    end else if (reset) begin
      release_state <= 4'h0;
    end else if (_T_316) begin
      release_state <= 4'h0;
    end else if (_T_312) begin
      if (releaseDone) begin
        release_state <= 4'h6;
      end else if (_T_307) begin
        if (releaseDone) begin
          release_state <= 4'h7;
        end else if (_T_306) begin
          if (releaseDone) begin
            release_state <= 4'h7;
          end else if (_T_305) begin
            if (releaseDone) begin
              release_state <= 4'h0;
            end else if (_T_304) begin
              if (metaArb_io_in_6_ready) begin
                release_state <= 4'h0;
              end else if (s2_probe) begin
                if (s2_meta_error) begin
                  release_state <= 4'h4;
                end else if (s2_prb_ack_data) begin
                  release_state <= 4'h2;
                end else if (_T_303) begin
                  if (releaseDone) begin
                    release_state <= 4'h7;
                  end else begin
                    release_state <= 4'h3;
                  end
                end else if (releaseDone) begin
                  release_state <= 4'h0;
                end else begin
                  release_state <= 4'h5;
                end
              end else if (s2_want_victimize) begin
                if (_release_state_T_1) begin
                  release_state <= 4'h1;
                end else begin
                  release_state <= 4'h6;
                end
              end
            end else if (s2_probe) begin
              if (s2_meta_error) begin
                release_state <= 4'h4;
              end else if (s2_prb_ack_data) begin
                release_state <= 4'h2;
              end else if (_T_303) begin
                if (releaseDone) begin
                  release_state <= 4'h7;
                end else begin
                  release_state <= 4'h3;
                end
              end else if (releaseDone) begin
                release_state <= 4'h0;
              end else begin
                release_state <= 4'h5;
              end
            end else if (s2_want_victimize) begin
              if (_release_state_T_1) begin
                release_state <= 4'h1;
              end else begin
                release_state <= 4'h6;
              end
            end
          end else if (_T_304) begin
            if (metaArb_io_in_6_ready) begin
              release_state <= 4'h0;
            end else if (s2_probe) begin
              if (s2_meta_error) begin
                release_state <= 4'h4;
              end else if (s2_prb_ack_data) begin
                release_state <= 4'h2;
              end else if (_T_303) begin
                if (releaseDone) begin
                  release_state <= 4'h7;
                end else begin
                  release_state <= 4'h3;
                end
              end else if (releaseDone) begin
                release_state <= 4'h0;
              end else begin
                release_state <= 4'h5;
              end
            end else if (s2_want_victimize) begin
              if (_release_state_T_1) begin
                release_state <= 4'h1;
              end else begin
                release_state <= 4'h6;
              end
            end
          end else if (s2_probe) begin
            if (s2_meta_error) begin
              release_state <= 4'h4;
            end else if (s2_prb_ack_data) begin
              release_state <= 4'h2;
            end else if (_T_303) begin
              if (releaseDone) begin
                release_state <= 4'h7;
              end else begin
                release_state <= 4'h3;
              end
            end else if (releaseDone) begin
              release_state <= 4'h0;
            end else begin
              release_state <= 4'h5;
            end
          end else if (s2_want_victimize) begin
            if (_release_state_T_1) begin
              release_state <= 4'h1;
            end else begin
              release_state <= 4'h6;
            end
          end
        end else if (_T_305) begin
          if (releaseDone) begin
            release_state <= 4'h0;
          end else if (_T_304) begin
            if (metaArb_io_in_6_ready) begin
              release_state <= 4'h0;
            end else begin
              release_state <= _GEN_284;
            end
          end else begin
            release_state <= _GEN_284;
          end
        end else if (_T_304) begin
          if (metaArb_io_in_6_ready) begin
            release_state <= 4'h0;
          end else begin
            release_state <= _GEN_284;
          end
        end else begin
          release_state <= _GEN_284;
        end
      end else if (_T_306) begin
        if (releaseDone) begin
          release_state <= 4'h7;
        end else if (_T_305) begin
          if (releaseDone) begin
            release_state <= 4'h0;
          end else begin
            release_state <= _GEN_299;
          end
        end else begin
          release_state <= _GEN_299;
        end
      end else if (_T_305) begin
        if (releaseDone) begin
          release_state <= 4'h0;
        end else begin
          release_state <= _GEN_299;
        end
      end else begin
        release_state <= _GEN_299;
      end
    end else if (_T_307) begin
      if (releaseDone) begin
        release_state <= 4'h7;
      end else if (_T_306) begin
        if (releaseDone) begin
          release_state <= 4'h7;
        end else begin
          release_state <= _GEN_303;
        end
      end else begin
        release_state <= _GEN_303;
      end
    end else if (_T_306) begin
      if (releaseDone) begin
        release_state <= 4'h7;
      end else begin
        release_state <= _GEN_303;
      end
    end else begin
      release_state <= _GEN_303;
    end
    if (metaReset) begin
      release_ack_wait <= 1'h0;
    end else if (reset) begin
      release_ack_wait <= 1'h0;
    end else if (_T_312) begin
      release_ack_wait <= _GEN_331;
    end else if (_T_271) begin
      if (!(grantIsCached)) begin
        if (!(grantIsUncached)) begin
          if (grantIsVoluntary) begin
            release_ack_wait <= 1'h0;
          end
        end
      end
    end
    if (metaReset) begin
      release_ack_addr <= 32'h0;
    end else if (_T_312) begin
      if (_T_315) begin
        release_ack_addr <= probe_bits_address;
      end
    end
    if (metaReset) begin
      grantInProgress <= 1'h0;
    end else if (reset) begin
      grantInProgress <= 1'h0;
    end else if (_T_271) begin
      if (grantIsCached) begin
        if (d_last) begin
          grantInProgress <= 1'h0;
        end else begin
          grantInProgress <= 1'h1;
        end
      end
    end
    if (metaReset) begin
      s2_valid <= 1'h0;
    end else if (reset) begin
      s2_valid <= 1'h0;
    end else begin
      s2_valid <= s2_valid_x37;
    end
    if (metaReset) begin
      probe_bits_param <= 2'h0;
    end else if (s2_want_victimize) begin
      probe_bits_param <= 2'h0;
    end else if (s1_probe_x12) begin
      probe_bits_param <= auto_out_b_bits_param;
    end
    if (metaReset) begin
      probe_bits_size <= 4'h0;
    end else if (s2_want_victimize) begin
      probe_bits_size <= 4'h0;
    end else if (s1_probe_x12) begin
      probe_bits_size <= auto_out_b_bits_size;
    end
    if (metaReset) begin
      probe_bits_source <= 1'h0;
    end else if (s2_want_victimize) begin
      probe_bits_source <= 1'h0;
    end else if (s1_probe_x12) begin
      probe_bits_source <= auto_out_b_bits_source;
    end
    if (metaReset) begin
      probe_bits_address <= 32'h0;
    end else if (s2_want_victimize) begin
      probe_bits_address <= res_2_address;
    end else if (s1_probe_x12) begin
      probe_bits_address <= auto_out_b_bits_address;
    end
    if (metaReset) begin
      s2_probe_state_state <= 2'h0;
    end else if (s1_probe) begin
      s2_probe_state_state <= s1_meta_hit_state_state;
    end
    if (metaReset) begin
      counter_1 <= 9'h0;
    end else if (reset) begin
      counter_1 <= 9'h0;
    end else if (_T_297) begin
      if (c_first) begin
        if (beats1_opdata_1) begin
          counter_1 <= beats1_decode_1;
        end else begin
          counter_1 <= 9'h0;
        end
      end else begin
        counter_1 <= counter1_1;
      end
    end
    if (metaReset) begin
      s2_release_data_valid <= 1'h0;
    end else begin
      s2_release_data_valid <= s1_release_data_valid & ~releaseRejected;
    end
    if (metaReset) begin
      s1_req_cmd <= 5'h0;
    end else if (s0_clk_en) begin
      s1_req_cmd <= io_cpu_req_bits_cmd;
    end
    if (metaReset) begin
      s2_req_cmd <= 5'h0;
    end else if (_T_271) begin
      if (grantIsCached) begin
        if (_T_70) begin
          s2_req_cmd <= s1_req_cmd;
        end
      end else if (grantIsUncached) begin
        if (grantIsUncachedData) begin
          s2_req_cmd <= 5'h0;
        end else if (_T_70) begin
          s2_req_cmd <= s1_req_cmd;
        end
      end else if (_T_70) begin
        s2_req_cmd <= s1_req_cmd;
      end
    end else if (_T_70) begin
      s2_req_cmd <= s1_req_cmd;
    end
    if (metaReset) begin
      pstore1_held <= 1'h0;
    end else if (reset) begin
      pstore1_held <= 1'h0;
    end else begin
      pstore1_held <= _pstore1_held_T_10;
    end
    if (metaReset) begin
      pstore1_addr <= 40'h0;
    end else if (_pstore1_cmd_T) begin
      pstore1_addr <= s1_vaddr;
    end
    if (metaReset) begin
      s1_req_addr <= 40'h0;
    end else if (s0_clk_en) begin
      s1_req_addr <= s0_req_addr;
    end
    if (metaReset) begin
      pstore1_mask <= 8'h0;
    end else if (_pstore1_cmd_T) begin
      if (_s1_write_T_1) begin
        pstore1_mask <= 8'h0;
      end else begin
        pstore1_mask <= s1_mask_xwr;
      end
    end
    if (metaReset) begin
      s1_req_size <= 2'h0;
    end else if (s0_clk_en) begin
      s1_req_size <= io_cpu_req_bits_size;
    end
    if (metaReset) begin
      pstore2_valid <= 1'h0;
    end else if (reset) begin
      pstore2_valid <= 1'h0;
    end else begin
      pstore2_valid <= _pstore2_valid_T_2;
    end
    if (metaReset) begin
      pstore2_addr <= 40'h0;
    end else if (advance_pstore1) begin
      pstore2_addr <= pstore1_addr;
    end
    if (metaReset) begin
      mask <= 8'h0;
    end else if (advance_pstore1) begin
      mask <= pstore1_mask[7:0];
    end
    if (metaReset) begin
      s2_not_nacked_in_s1 <= 1'h0;
    end else begin
      s2_not_nacked_in_s1 <= ~s1_nack;
    end
    if (metaReset) begin
      s2_hit_state_state <= 2'h0;
    end else if (_T_70) begin
      s2_hit_state_state <= s1_meta_hit_state_state;
    end
    if (metaReset) begin
      s1_req_tag <= 7'h0;
    end else if (s0_clk_en) begin
      s1_req_tag <= io_cpu_req_bits_tag;
    end
    if (metaReset) begin
      s1_req_signed <= 1'h0;
    end else if (s0_clk_en) begin
      s1_req_signed <= io_cpu_req_bits_signed;
    end
    if (metaReset) begin
      s1_tlb_req_vaddr <= 40'h0;
    end else if (s0_clk_en) begin
      s1_tlb_req_vaddr <= s0_req_addr;
    end
    if (metaReset) begin
      s1_tlb_req_passthrough <= 1'h0;
    end else if (s0_clk_en) begin
      s1_tlb_req_passthrough <= s0_req_phys;
    end
    if (metaReset) begin
      s1_tlb_req_size <= 2'h0;
    end else if (s0_clk_en) begin
      s1_tlb_req_size <= io_cpu_req_bits_size;
    end
    if (metaReset) begin
      s1_tlb_req_cmd <= 5'h0;
    end else if (s0_clk_en) begin
      s1_tlb_req_cmd <= io_cpu_req_bits_cmd;
    end
    if (metaReset) begin
      s1_flush_valid <= 1'h0;
    end else begin
      s1_flush_valid <= _s1_flush_valid_T_6 & ~release_ack_wait;
    end
    if (metaReset) begin
      cached_grant_wait <= 1'h0;
    end else if (reset) begin
      cached_grant_wait <= 1'h0;
    end else if (_T_271) begin
      if (grantIsCached) begin
        if (d_last) begin
          cached_grant_wait <= 1'h0;
        end else if (_T_263) begin
          if (!(s2_uncached)) begin
            cached_grant_wait <= 1'h1;
          end
        end
      end else if (_T_263) begin
        if (!(s2_uncached)) begin
          cached_grant_wait <= 1'h1;
        end
      end
    end else if (_T_263) begin
      if (!(s2_uncached)) begin
        cached_grant_wait <= 1'h1;
      end
    end
    if (metaReset) begin
      resetting <= 1'h0;
    end else if (reset) begin
      resetting <= 1'h0;
    end else if (resetting) begin
      if (flushDone) begin
        resetting <= 1'h0;
      end else begin
        resetting <= _GEN_349;
      end
    end else begin
      resetting <= _GEN_349;
    end
    if (metaReset) begin
      flushCounter <= 8'h0;
    end else if (reset) begin
      flushCounter <= 8'hc0;
    end else begin
      flushCounter <= _GEN_351[7:0];
    end
    if (metaReset) begin
      refill_way <= 4'h0;
    end else if (_T_263) begin
      if (!(s2_uncached)) begin
        if (s2_hit_valid) begin
          refill_way <= s2_hit_way;
        end else begin
          refill_way <= s2_victim_way;
        end
      end
    end
    if (metaReset) begin
      uncachedInFlight_0 <= 1'h0;
    end else if (reset) begin
      uncachedInFlight_0 <= 1'h0;
    end else if (_T_271) begin
      if (grantIsCached) begin
        if (_T_263) begin
          if (s2_uncached) begin
            uncachedInFlight_0 <= _GEN_142;
          end
        end
      end else if (grantIsUncached) begin
        if (_T_276) begin
          uncachedInFlight_0 <= 1'h0;
        end else if (_T_263) begin
          if (s2_uncached) begin
            uncachedInFlight_0 <= _GEN_142;
          end
        end
      end else if (_T_263) begin
        if (s2_uncached) begin
          uncachedInFlight_0 <= _GEN_142;
        end
      end
    end else if (_T_263) begin
      if (s2_uncached) begin
        uncachedInFlight_0 <= _GEN_142;
      end
    end
    if (metaReset) begin
      uncachedReqs_0_addr <= 40'h0;
    end else if (_T_263) begin
      if (s2_uncached) begin
        if (a_sel) begin
          uncachedReqs_0_addr <= s2_req_addr;
        end
      end
    end
    if (metaReset) begin
      uncachedReqs_0_tag <= 7'h0;
    end else if (_T_263) begin
      if (s2_uncached) begin
        if (a_sel) begin
          uncachedReqs_0_tag <= s2_req_tag;
        end
      end
    end
    if (metaReset) begin
      uncachedReqs_0_size <= 2'h0;
    end else if (_T_263) begin
      if (s2_uncached) begin
        if (a_sel) begin
          uncachedReqs_0_size <= s2_req_size;
        end
      end
    end
    if (metaReset) begin
      uncachedReqs_0_signed <= 1'h0;
    end else if (_T_263) begin
      if (s2_uncached) begin
        if (a_sel) begin
          uncachedReqs_0_signed <= s2_req_signed;
        end
      end
    end
    if (metaReset) begin
      s1_did_read <= 1'h0;
    end else if (s0_clk_en) begin
      s1_did_read <= _s1_did_read_T_52;
    end
    if (metaReset) begin
      s1_read_mask <= 1'h0;
    end else if (s0_clk_en) begin
      s1_read_mask <= dataArb_io_in_3_bits_wordMask;
    end
    if (metaReset) begin
      s2_hit_way <= 4'h0;
    end else if (s1_valid_not_nacked) begin
      s2_hit_way <= s1_meta_hit_way;
    end
    if (metaReset) begin
      s2_victim_way_r <= 2'h0;
    end else if (_T_70) begin
      s2_victim_way_r <= s1_victim_way;
    end
    if (metaReset) begin
      s2_probe_way <= 4'h0;
    end else if (s1_probe) begin
      s2_probe_way <= s1_meta_hit_way;
    end
    if (metaReset) begin
      s2_req_addr <= 40'h0;
    end else if (_T_271) begin
      if (grantIsCached) begin
        if (_T_70) begin
          s2_req_addr <= {{8'd0}, s1_paddr};
        end
      end else if (grantIsUncached) begin
        if (grantIsUncachedData) begin
          s2_req_addr <= {{8'd0}, _s2_req_addr_T_1};
        end else if (_T_70) begin
          s2_req_addr <= {{8'd0}, s1_paddr};
        end
      end else if (_T_70) begin
        s2_req_addr <= {{8'd0}, s1_paddr};
      end
    end else if (_T_70) begin
      s2_req_addr <= {{8'd0}, s1_paddr};
    end
    if (metaReset) begin
      s2_req_tag <= 7'h0;
    end else if (_T_271) begin
      if (grantIsCached) begin
        if (_T_70) begin
          s2_req_tag <= s1_req_tag;
        end
      end else if (grantIsUncached) begin
        if (grantIsUncachedData) begin
          s2_req_tag <= uncachedReqs_0_tag;
        end else if (_T_70) begin
          s2_req_tag <= s1_req_tag;
        end
      end else if (_T_70) begin
        s2_req_tag <= s1_req_tag;
      end
    end else if (_T_70) begin
      s2_req_tag <= s1_req_tag;
    end
    if (metaReset) begin
      s2_req_size <= 2'h0;
    end else if (_T_271) begin
      if (grantIsCached) begin
        if (_T_70) begin
          s2_req_size <= s1_req_size;
        end
      end else if (grantIsUncached) begin
        if (grantIsUncachedData) begin
          s2_req_size <= uncachedReqs_0_size;
        end else if (_T_70) begin
          s2_req_size <= s1_req_size;
        end
      end else if (_T_70) begin
        s2_req_size <= s1_req_size;
      end
    end else if (_T_70) begin
      s2_req_size <= s1_req_size;
    end
    if (metaReset) begin
      s2_req_signed <= 1'h0;
    end else if (_T_271) begin
      if (grantIsCached) begin
        if (_T_70) begin
          s2_req_signed <= s1_req_signed;
        end
      end else if (grantIsUncached) begin
        if (grantIsUncachedData) begin
          s2_req_signed <= uncachedReqs_0_signed;
        end else if (_T_70) begin
          s2_req_signed <= s1_req_signed;
        end
      end else if (_T_70) begin
        s2_req_signed <= s1_req_signed;
      end
    end else if (_T_70) begin
      s2_req_signed <= s1_req_signed;
    end
    if (metaReset) begin
      s2_tlb_xcpt_pf_ld <= 1'h0;
    end else if (_T_70) begin
      s2_tlb_xcpt_pf_ld <= tlb_io_resp_pf_ld;
    end
    if (metaReset) begin
      s2_tlb_xcpt_pf_st <= 1'h0;
    end else if (_T_70) begin
      s2_tlb_xcpt_pf_st <= tlb_io_resp_pf_st;
    end
    if (metaReset) begin
      s2_tlb_xcpt_ae_ld <= 1'h0;
    end else if (_T_70) begin
      s2_tlb_xcpt_ae_ld <= tlb_io_resp_ae_ld;
    end
    if (metaReset) begin
      s2_tlb_xcpt_ae_st <= 1'h0;
    end else if (_T_70) begin
      s2_tlb_xcpt_ae_st <= tlb_io_resp_ae_st;
    end
    if (metaReset) begin
      s2_tlb_xcpt_ma_ld <= 1'h0;
    end else if (_T_70) begin
      s2_tlb_xcpt_ma_ld <= tlb_io_resp_ma_ld;
    end
    if (metaReset) begin
      s2_tlb_xcpt_ma_st <= 1'h0;
    end else if (_T_70) begin
      s2_tlb_xcpt_ma_st <= tlb_io_resp_ma_st;
    end
    if (metaReset) begin
      s2_pma_cacheable <= 1'h0;
    end else if (_T_70) begin
      s2_pma_cacheable <= _s2_pma_T_cacheable;
    end
    if (metaReset) begin
      s2_vaddr_r <= 40'h0;
    end else if (_T_70) begin
      s2_vaddr_r <= s1_vaddr;
    end
    if (metaReset) begin
      s2_flush_valid_pre_tag_ecc <= 1'h0;
    end else begin
      s2_flush_valid_pre_tag_ecc <= s1_flush_valid;
    end
    if (metaReset) begin
      s2_meta_corrected_r <= 22'h0;
    end else if (s1_meta_clk_en) begin
      s2_meta_corrected_r <= tag_array_0_s1_meta_data;
    end
    if (metaReset) begin
      s2_meta_corrected_r_1 <= 22'h0;
    end else if (s1_meta_clk_en) begin
      s2_meta_corrected_r_1 <= tag_array_1_s1_meta_data;
    end
    if (metaReset) begin
      s2_meta_corrected_r_2 <= 22'h0;
    end else if (s1_meta_clk_en) begin
      s2_meta_corrected_r_2 <= tag_array_2_s1_meta_data;
    end
    if (metaReset) begin
      s2_meta_corrected_r_3 <= 22'h0;
    end else if (s1_meta_clk_en) begin
      s2_meta_corrected_r_3 <= tag_array_3_s1_meta_data;
    end
    if (metaReset) begin
      blockUncachedGrant <= 1'h0;
    end else if (_T_294) begin
      if (auto_out_d_valid) begin
        blockUncachedGrant <= ~dataArb_io_in_1_ready;
      end else begin
        blockUncachedGrant <= dataArb_io_out_valid;
      end
    end else begin
      blockUncachedGrant <= dataArb_io_out_valid;
    end
    if (metaReset) begin
      counter <= 9'h0;
    end else if (reset) begin
      counter <= 9'h0;
    end else if (_T_271) begin
      if (d_first) begin
        if (beats1_opdata) begin
          counter <= beats1_decode;
        end else begin
          counter <= 9'h0;
        end
      end else begin
        counter <= counter1;
      end
    end
    if (metaReset) begin
      s2_data <= 64'h0;
    end else if (en) begin
      s2_data <= _s2_data_T_15;
    end
    if (metaReset) begin
      lrscAddr <= 34'h0;
    end else if (_T_246) begin
      lrscAddr <= s2_req_addr[39:6];
    end
    if (metaReset) begin
      pstore1_cmd <= 5'h0;
    end else if (_pstore1_cmd_T) begin
      pstore1_cmd <= s1_req_cmd;
    end
    if (metaReset) begin
      pstore1_data <= 64'h0;
    end else if (_pstore1_cmd_T) begin
      pstore1_data <= io_cpu_s1_data_data;
    end
    if (metaReset) begin
      pstore1_way <= 4'h0;
    end else if (_pstore1_cmd_T) begin
      pstore1_way <= s1_meta_hit_way;
    end
    if (metaReset) begin
      pstore1_rmw_r <= 1'h0;
    end else if (_pstore1_cmd_T) begin
      pstore1_rmw_r <= _pstore1_rmw_T_50;
    end
    if (metaReset) begin
      pstore_drain_on_miss_REG <= 1'h0;
    end else begin
      pstore_drain_on_miss_REG <= io_cpu_s2_nack;
    end
    if (metaReset) begin
      pstore2_way <= 4'h0;
    end else if (advance_pstore1) begin
      pstore2_way <= pstore1_way;
    end
    if (metaReset) begin
      pstore2_storegen_data_lo_lo_lo <= 8'h0;
    end else if (advance_pstore1) begin
      pstore2_storegen_data_lo_lo_lo <= pstore1_storegen_data[7:0];
    end
    if (metaReset) begin
      pstore2_storegen_data_lo_lo_hi <= 8'h0;
    end else if (advance_pstore1) begin
      pstore2_storegen_data_lo_lo_hi <= pstore1_storegen_data[15:8];
    end
    if (metaReset) begin
      pstore2_storegen_data_lo_hi_lo <= 8'h0;
    end else if (advance_pstore1) begin
      pstore2_storegen_data_lo_hi_lo <= pstore1_storegen_data[23:16];
    end
    if (metaReset) begin
      pstore2_storegen_data_lo_hi_hi <= 8'h0;
    end else if (advance_pstore1) begin
      pstore2_storegen_data_lo_hi_hi <= pstore1_storegen_data[31:24];
    end
    if (metaReset) begin
      pstore2_storegen_data_hi_lo_lo <= 8'h0;
    end else if (advance_pstore1) begin
      pstore2_storegen_data_hi_lo_lo <= pstore1_storegen_data[39:32];
    end
    if (metaReset) begin
      pstore2_storegen_data_hi_lo_hi <= 8'h0;
    end else if (advance_pstore1) begin
      pstore2_storegen_data_hi_lo_hi <= pstore1_storegen_data[47:40];
    end
    if (metaReset) begin
      pstore2_storegen_data_hi_hi_lo <= 8'h0;
    end else if (advance_pstore1) begin
      pstore2_storegen_data_hi_hi_lo <= pstore1_storegen_data[55:48];
    end
    if (metaReset) begin
      pstore2_storegen_data_hi_hi_hi <= 8'h0;
    end else if (advance_pstore1) begin
      pstore2_storegen_data_hi_hi_hi <= pstore1_storegen_data[63:56];
    end
    if (metaReset) begin
      s1_release_data_valid <= 1'h0;
    end else begin
      s1_release_data_valid <= dataArb_io_in_2_ready & dataArb_io_in_2_valid;
    end
    if (metaReset) begin
      io_cpu_s2_xcpt_REG <= 1'h0;
    end else begin
      io_cpu_s2_xcpt_REG <= _s1_xcpt_valid_T_1 & ~s1_nack;
    end
    if (metaReset) begin
      doUncachedResp <= 1'h0;
    end else begin
      doUncachedResp <= io_cpu_replay_next;
    end
    if (metaReset) begin
      REG <= 1'h0;
    end else begin
      REG <= reset;
    end
    if (metaReset) begin
      io_cpu_perf_release_counter <= 9'h0;
    end else if (reset) begin
      io_cpu_perf_release_counter <= 9'h0;
    end else if (_T_297) begin
      if (io_cpu_perf_release_first) begin
        if (beats1_opdata_1) begin
          io_cpu_perf_release_counter <= beats1_decode_1;
        end else begin
          io_cpu_perf_release_counter <= 9'h0;
        end
      end else begin
        io_cpu_perf_release_counter <= io_cpu_perf_release_counter1;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_dataArb_io_in_3_valid_T_54) begin
          $fwrite(32'h80000002,"Assertion failed\n    at DCache.scala:1154 assert(!needsRead(req) || res)\n"); // @[DCache.scala 1154:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_dataArb_io_in_3_valid_T_54) begin
          $fatal; // @[DCache.scala 1154:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_68) begin
          $fwrite(32'h80000002,"Assertion failed\n    at DCache.scala:300 assert(!(s1_valid_masked && s1_req.cmd === M_PWR) || (s1_mask_xwr | ~io.cpu.s1_data.mask).andR)\n"); // @[DCache.scala 300:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_68) begin
          $fatal; // @[DCache.scala 300:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_dataArb_io_in_3_valid_T_54) begin
          $fwrite(32'h80000002,"Assertion failed\n    at DCache.scala:1154 assert(!needsRead(req) || res)\n"); // @[DCache.scala 1154:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_dataArb_io_in_3_valid_T_54) begin
          $fatal; // @[DCache.scala 1154:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_258) begin
          $fwrite(32'h80000002,"Assertion failed\n    at DCache.scala:481 assert(pstore1_rmw || pstore1_valid_not_rmw(io.cpu.s2_kill) === pstore1_valid)\n"); // @[DCache.scala 481:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_258) begin
          $fatal; // @[DCache.scala 481:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_367 & ~_T_273) begin
          $fwrite(32'h80000002,"Assertion failed: A GrantData was unexpected by the dcache.\n    at DCache.scala:648 assert(cached_grant_wait, \"A GrantData was unexpected by the dcache.\")\n"); // @[DCache.scala 648:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_367 & ~_T_273) begin
          $fatal; // @[DCache.scala 648:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_372 & ~_T_278) begin
          $fwrite(32'h80000002,"Assertion failed: An AccessAck was unexpected by the dcache.\n    at DCache.scala:658 assert(f, \"An AccessAck was unexpected by the dcache.\") // TODO must handle Ack coming back on same cycle!\n"); // @[DCache.scala 658:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_372 & ~_T_278) begin
          $fatal; // @[DCache.scala 658:17]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_381 & ~_T_281) begin
          $fwrite(32'h80000002,"Assertion failed: A ReleaseAck was unexpected by the dcache.\n    at DCache.scala:679 assert(release_ack_wait, \"A ReleaseAck was unexpected by the dcache.\") // TODO should handle Ack coming back on same cycle!\n"); // @[DCache.scala 679:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_381 & ~_T_281) begin
          $fatal; // @[DCache.scala 679:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_289) begin
          $fwrite(32'h80000002,"Assertion failed\n    at DCache.scala:687 assert(tl_out.e.fire() === (tl_out.d.fire() && d_first && grantIsCached))\n"); // @[DCache.scala 687:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_289) begin
          $fatal; // @[DCache.scala 687:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (s2_want_victimize & ~_T_301) begin
          $fwrite(32'h80000002,"Assertion failed\n    at DCache.scala:788 assert(s2_valid_flush_line || s2_flush_valid || io.cpu.s2_nack)\n"); // @[DCache.scala 788:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (s2_want_victimize & ~_T_301) begin
          $fatal; // @[DCache.scala 788:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (doUncachedResp & ~_T_321) begin
          $fwrite(32'h80000002,"Assertion failed\n    at DCache.scala:920 assert(!s2_valid_hit)\n"); // @[DCache.scala 920:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (doUncachedResp & ~_T_321) begin
          $fatal; // @[DCache.scala 920:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    DCache_state <= DCache_xor0;
    if (!(DCache_cov_read_data)) begin
      DCache_covSum <= DCache_covSum + 1'h1;
    end
  end
  always @(posedge gated_clock) begin
    if(DCache_cov_write_en & DCache_cov_write_mask) begin
      DCache_cov[DCache_cov_write_addr] <= DCache_cov_write_data; // @[Coverage map for DCache]
    end
  end
endmodule
module Frontend(
  input         gated_clock,
  input         reset,
  input         auto_icache_master_out_a_ready,
  output        auto_icache_master_out_a_valid,
  output [31:0] auto_icache_master_out_a_bits_address,
  input         auto_icache_master_out_d_valid,
  input  [2:0]  auto_icache_master_out_d_bits_opcode,
  input  [3:0]  auto_icache_master_out_d_bits_size,
  input  [63:0] auto_icache_master_out_d_bits_data,
  input         auto_icache_master_out_d_bits_corrupt,
  input  [31:0] auto_reset_vector_sink_in,
  input         io_cpu_might_request,
  input         io_cpu_req_valid,
  input  [39:0] io_cpu_req_bits_pc,
  input         io_cpu_req_bits_speculative,
  input         io_cpu_sfence_valid,
  input         io_cpu_sfence_bits_rs1,
  input         io_cpu_sfence_bits_rs2,
  input  [38:0] io_cpu_sfence_bits_addr,
  input         io_cpu_resp_ready,
  output        io_cpu_resp_valid,
  output        io_cpu_resp_bits_btb_taken,
  output        io_cpu_resp_bits_btb_bridx,
  output [4:0]  io_cpu_resp_bits_btb_entry,
  output [7:0]  io_cpu_resp_bits_btb_bht_history,
  output [39:0] io_cpu_resp_bits_pc,
  output [31:0] io_cpu_resp_bits_data,
  output        io_cpu_resp_bits_xcpt_pf_inst,
  output        io_cpu_resp_bits_xcpt_ae_inst,
  output        io_cpu_resp_bits_replay,
  input         io_cpu_btb_update_valid,
  input  [4:0]  io_cpu_btb_update_bits_prediction_entry,
  input  [38:0] io_cpu_btb_update_bits_pc,
  input         io_cpu_btb_update_bits_isValid,
  input  [38:0] io_cpu_btb_update_bits_br_pc,
  input  [1:0]  io_cpu_btb_update_bits_cfiType,
  input         io_cpu_bht_update_valid,
  input  [7:0]  io_cpu_bht_update_bits_prediction_history,
  input  [38:0] io_cpu_bht_update_bits_pc,
  input         io_cpu_bht_update_bits_branch,
  input         io_cpu_bht_update_bits_taken,
  input         io_cpu_bht_update_bits_mispredict,
  input         io_cpu_flush_icache,
  output [39:0] io_cpu_npc,
  input         io_ptw_req_ready,
  output        io_ptw_req_valid,
  output        io_ptw_req_bits_valid,
  output [26:0] io_ptw_req_bits_bits_addr,
  input         io_ptw_resp_valid,
  input         io_ptw_resp_bits_ae,
  input  [53:0] io_ptw_resp_bits_pte_ppn,
  input         io_ptw_resp_bits_pte_d,
  input         io_ptw_resp_bits_pte_a,
  input         io_ptw_resp_bits_pte_g,
  input         io_ptw_resp_bits_pte_u,
  input         io_ptw_resp_bits_pte_x,
  input         io_ptw_resp_bits_pte_w,
  input         io_ptw_resp_bits_pte_r,
  input         io_ptw_resp_bits_pte_v,
  input  [1:0]  io_ptw_resp_bits_level,
  input         io_ptw_resp_bits_homogeneous,
  input  [3:0]  io_ptw_ptbr_mode,
  input         io_ptw_status_debug,
  input  [1:0]  io_ptw_status_prv,
  input         io_ptw_pmp_0_cfg_l,
  input  [1:0]  io_ptw_pmp_0_cfg_a,
  input         io_ptw_pmp_0_cfg_x,
  input         io_ptw_pmp_0_cfg_w,
  input         io_ptw_pmp_0_cfg_r,
  input  [29:0] io_ptw_pmp_0_addr,
  input  [31:0] io_ptw_pmp_0_mask,
  input         io_ptw_pmp_1_cfg_l,
  input  [1:0]  io_ptw_pmp_1_cfg_a,
  input         io_ptw_pmp_1_cfg_x,
  input         io_ptw_pmp_1_cfg_w,
  input         io_ptw_pmp_1_cfg_r,
  input  [29:0] io_ptw_pmp_1_addr,
  input  [31:0] io_ptw_pmp_1_mask,
  input         io_ptw_pmp_2_cfg_l,
  input  [1:0]  io_ptw_pmp_2_cfg_a,
  input         io_ptw_pmp_2_cfg_x,
  input         io_ptw_pmp_2_cfg_w,
  input         io_ptw_pmp_2_cfg_r,
  input  [29:0] io_ptw_pmp_2_addr,
  input  [31:0] io_ptw_pmp_2_mask,
  input         io_ptw_pmp_3_cfg_l,
  input  [1:0]  io_ptw_pmp_3_cfg_a,
  input         io_ptw_pmp_3_cfg_x,
  input         io_ptw_pmp_3_cfg_w,
  input         io_ptw_pmp_3_cfg_r,
  input  [29:0] io_ptw_pmp_3_addr,
  input  [31:0] io_ptw_pmp_3_mask,
  input         io_ptw_pmp_4_cfg_l,
  input  [1:0]  io_ptw_pmp_4_cfg_a,
  input         io_ptw_pmp_4_cfg_x,
  input         io_ptw_pmp_4_cfg_w,
  input         io_ptw_pmp_4_cfg_r,
  input  [29:0] io_ptw_pmp_4_addr,
  input  [31:0] io_ptw_pmp_4_mask,
  input         io_ptw_pmp_5_cfg_l,
  input  [1:0]  io_ptw_pmp_5_cfg_a,
  input         io_ptw_pmp_5_cfg_x,
  input         io_ptw_pmp_5_cfg_w,
  input         io_ptw_pmp_5_cfg_r,
  input  [29:0] io_ptw_pmp_5_addr,
  input  [31:0] io_ptw_pmp_5_mask,
  input         io_ptw_pmp_6_cfg_l,
  input  [1:0]  io_ptw_pmp_6_cfg_a,
  input         io_ptw_pmp_6_cfg_x,
  input         io_ptw_pmp_6_cfg_w,
  input         io_ptw_pmp_6_cfg_r,
  input  [29:0] io_ptw_pmp_6_addr,
  input  [31:0] io_ptw_pmp_6_mask,
  input         io_ptw_pmp_7_cfg_l,
  input  [1:0]  io_ptw_pmp_7_cfg_a,
  input         io_ptw_pmp_7_cfg_x,
  input         io_ptw_pmp_7_cfg_w,
  input         io_ptw_pmp_7_cfg_r,
  input  [29:0] io_ptw_pmp_7_addr,
  input  [31:0] io_ptw_pmp_7_mask,
  input  [63:0] io_ptw_customCSRs_csrs_0_value,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset,
  input         icache_halt,
  input         fq_halt,
  input         tlb_halt,
  input         btb_halt
);
  wire  icache_clock; // @[Frontend.scala 62:26]
  wire  icache_reset; // @[Frontend.scala 62:26]
  wire  icache_auto_master_out_a_ready; // @[Frontend.scala 62:26]
  wire  icache_auto_master_out_a_valid; // @[Frontend.scala 62:26]
  wire [31:0] icache_auto_master_out_a_bits_address; // @[Frontend.scala 62:26]
  wire  icache_auto_master_out_d_valid; // @[Frontend.scala 62:26]
  wire [2:0] icache_auto_master_out_d_bits_opcode; // @[Frontend.scala 62:26]
  wire [3:0] icache_auto_master_out_d_bits_size; // @[Frontend.scala 62:26]
  wire [63:0] icache_auto_master_out_d_bits_data; // @[Frontend.scala 62:26]
  wire  icache_auto_master_out_d_bits_corrupt; // @[Frontend.scala 62:26]
  wire  icache_io_req_ready; // @[Frontend.scala 62:26]
  wire  icache_io_req_valid; // @[Frontend.scala 62:26]
  wire [38:0] icache_io_req_bits_addr; // @[Frontend.scala 62:26]
  wire [31:0] icache_io_s1_paddr; // @[Frontend.scala 62:26]
  wire  icache_io_s1_kill; // @[Frontend.scala 62:26]
  wire  icache_io_s2_kill; // @[Frontend.scala 62:26]
  wire  icache_io_resp_valid; // @[Frontend.scala 62:26]
  wire [31:0] icache_io_resp_bits_data; // @[Frontend.scala 62:26]
  wire  icache_io_resp_bits_replay; // @[Frontend.scala 62:26]
  wire  icache_io_resp_bits_ae; // @[Frontend.scala 62:26]
  wire  icache_io_invalidate; // @[Frontend.scala 62:26]
  wire [29:0] icache_io_covSum; // @[Frontend.scala 62:26]
  wire  icache_metaAssert; // @[Frontend.scala 62:26]
  wire  icache_metaReset; // @[Frontend.scala 62:26]
  wire  icache_repl_way_v0_prng_halt; // @[Frontend.scala 62:26]
  wire  fq_clock; // @[Frontend.scala 84:57]
  wire  fq_reset; // @[Frontend.scala 84:57]
  wire  fq_io_enq_ready; // @[Frontend.scala 84:57]
  wire  fq_io_enq_valid; // @[Frontend.scala 84:57]
  wire  fq_io_enq_bits_btb_taken; // @[Frontend.scala 84:57]
  wire  fq_io_enq_bits_btb_bridx; // @[Frontend.scala 84:57]
  wire [4:0] fq_io_enq_bits_btb_entry; // @[Frontend.scala 84:57]
  wire [7:0] fq_io_enq_bits_btb_bht_history; // @[Frontend.scala 84:57]
  wire [39:0] fq_io_enq_bits_pc; // @[Frontend.scala 84:57]
  wire [31:0] fq_io_enq_bits_data; // @[Frontend.scala 84:57]
  wire [1:0] fq_io_enq_bits_mask; // @[Frontend.scala 84:57]
  wire  fq_io_enq_bits_xcpt_pf_inst; // @[Frontend.scala 84:57]
  wire  fq_io_enq_bits_xcpt_ae_inst; // @[Frontend.scala 84:57]
  wire  fq_io_enq_bits_replay; // @[Frontend.scala 84:57]
  wire  fq_io_deq_ready; // @[Frontend.scala 84:57]
  wire  fq_io_deq_valid; // @[Frontend.scala 84:57]
  wire  fq_io_deq_bits_btb_taken; // @[Frontend.scala 84:57]
  wire  fq_io_deq_bits_btb_bridx; // @[Frontend.scala 84:57]
  wire [4:0] fq_io_deq_bits_btb_entry; // @[Frontend.scala 84:57]
  wire [7:0] fq_io_deq_bits_btb_bht_history; // @[Frontend.scala 84:57]
  wire [39:0] fq_io_deq_bits_pc; // @[Frontend.scala 84:57]
  wire [31:0] fq_io_deq_bits_data; // @[Frontend.scala 84:57]
  wire  fq_io_deq_bits_xcpt_pf_inst; // @[Frontend.scala 84:57]
  wire  fq_io_deq_bits_xcpt_ae_inst; // @[Frontend.scala 84:57]
  wire  fq_io_deq_bits_replay; // @[Frontend.scala 84:57]
  wire [4:0] fq_io_mask; // @[Frontend.scala 84:57]
  wire [29:0] fq_io_covSum; // @[Frontend.scala 84:57]
  wire  fq_metaAssert; // @[Frontend.scala 84:57]
  wire  fq_metaReset; // @[Frontend.scala 84:57]
  wire  tlb_clock; // @[Frontend.scala 98:19]
  wire  tlb_reset; // @[Frontend.scala 98:19]
  wire  tlb_io_req_ready; // @[Frontend.scala 98:19]
  wire  tlb_io_req_valid; // @[Frontend.scala 98:19]
  wire [39:0] tlb_io_req_bits_vaddr; // @[Frontend.scala 98:19]
  wire  tlb_io_resp_miss; // @[Frontend.scala 98:19]
  wire [31:0] tlb_io_resp_paddr; // @[Frontend.scala 98:19]
  wire  tlb_io_resp_pf_inst; // @[Frontend.scala 98:19]
  wire  tlb_io_resp_ae_inst; // @[Frontend.scala 98:19]
  wire  tlb_io_resp_cacheable; // @[Frontend.scala 98:19]
  wire  tlb_io_sfence_valid; // @[Frontend.scala 98:19]
  wire  tlb_io_sfence_bits_rs1; // @[Frontend.scala 98:19]
  wire  tlb_io_sfence_bits_rs2; // @[Frontend.scala 98:19]
  wire [38:0] tlb_io_sfence_bits_addr; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_req_ready; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_req_valid; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_req_bits_valid; // @[Frontend.scala 98:19]
  wire [26:0] tlb_io_ptw_req_bits_bits_addr; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_resp_valid; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_resp_bits_ae; // @[Frontend.scala 98:19]
  wire [53:0] tlb_io_ptw_resp_bits_pte_ppn; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_resp_bits_pte_d; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_resp_bits_pte_a; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_resp_bits_pte_g; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_resp_bits_pte_u; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_resp_bits_pte_x; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_resp_bits_pte_w; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_resp_bits_pte_r; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_resp_bits_pte_v; // @[Frontend.scala 98:19]
  wire [1:0] tlb_io_ptw_resp_bits_level; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_resp_bits_homogeneous; // @[Frontend.scala 98:19]
  wire [3:0] tlb_io_ptw_ptbr_mode; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_status_debug; // @[Frontend.scala 98:19]
  wire [1:0] tlb_io_ptw_status_prv; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_pmp_0_cfg_l; // @[Frontend.scala 98:19]
  wire [1:0] tlb_io_ptw_pmp_0_cfg_a; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_pmp_0_cfg_x; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_pmp_0_cfg_w; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_pmp_0_cfg_r; // @[Frontend.scala 98:19]
  wire [29:0] tlb_io_ptw_pmp_0_addr; // @[Frontend.scala 98:19]
  wire [31:0] tlb_io_ptw_pmp_0_mask; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_pmp_1_cfg_l; // @[Frontend.scala 98:19]
  wire [1:0] tlb_io_ptw_pmp_1_cfg_a; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_pmp_1_cfg_x; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_pmp_1_cfg_w; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_pmp_1_cfg_r; // @[Frontend.scala 98:19]
  wire [29:0] tlb_io_ptw_pmp_1_addr; // @[Frontend.scala 98:19]
  wire [31:0] tlb_io_ptw_pmp_1_mask; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_pmp_2_cfg_l; // @[Frontend.scala 98:19]
  wire [1:0] tlb_io_ptw_pmp_2_cfg_a; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_pmp_2_cfg_x; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_pmp_2_cfg_w; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_pmp_2_cfg_r; // @[Frontend.scala 98:19]
  wire [29:0] tlb_io_ptw_pmp_2_addr; // @[Frontend.scala 98:19]
  wire [31:0] tlb_io_ptw_pmp_2_mask; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_pmp_3_cfg_l; // @[Frontend.scala 98:19]
  wire [1:0] tlb_io_ptw_pmp_3_cfg_a; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_pmp_3_cfg_x; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_pmp_3_cfg_w; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_pmp_3_cfg_r; // @[Frontend.scala 98:19]
  wire [29:0] tlb_io_ptw_pmp_3_addr; // @[Frontend.scala 98:19]
  wire [31:0] tlb_io_ptw_pmp_3_mask; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_pmp_4_cfg_l; // @[Frontend.scala 98:19]
  wire [1:0] tlb_io_ptw_pmp_4_cfg_a; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_pmp_4_cfg_x; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_pmp_4_cfg_w; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_pmp_4_cfg_r; // @[Frontend.scala 98:19]
  wire [29:0] tlb_io_ptw_pmp_4_addr; // @[Frontend.scala 98:19]
  wire [31:0] tlb_io_ptw_pmp_4_mask; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_pmp_5_cfg_l; // @[Frontend.scala 98:19]
  wire [1:0] tlb_io_ptw_pmp_5_cfg_a; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_pmp_5_cfg_x; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_pmp_5_cfg_w; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_pmp_5_cfg_r; // @[Frontend.scala 98:19]
  wire [29:0] tlb_io_ptw_pmp_5_addr; // @[Frontend.scala 98:19]
  wire [31:0] tlb_io_ptw_pmp_5_mask; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_pmp_6_cfg_l; // @[Frontend.scala 98:19]
  wire [1:0] tlb_io_ptw_pmp_6_cfg_a; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_pmp_6_cfg_x; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_pmp_6_cfg_w; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_pmp_6_cfg_r; // @[Frontend.scala 98:19]
  wire [29:0] tlb_io_ptw_pmp_6_addr; // @[Frontend.scala 98:19]
  wire [31:0] tlb_io_ptw_pmp_6_mask; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_pmp_7_cfg_l; // @[Frontend.scala 98:19]
  wire [1:0] tlb_io_ptw_pmp_7_cfg_a; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_pmp_7_cfg_x; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_pmp_7_cfg_w; // @[Frontend.scala 98:19]
  wire  tlb_io_ptw_pmp_7_cfg_r; // @[Frontend.scala 98:19]
  wire [29:0] tlb_io_ptw_pmp_7_addr; // @[Frontend.scala 98:19]
  wire [31:0] tlb_io_ptw_pmp_7_mask; // @[Frontend.scala 98:19]
  wire  tlb_io_kill; // @[Frontend.scala 98:19]
  wire [29:0] tlb_io_covSum; // @[Frontend.scala 98:19]
  wire  tlb_metaAssert; // @[Frontend.scala 98:19]
  wire  tlb_metaReset; // @[Frontend.scala 98:19]
  wire  btb_clock; // @[Frontend.scala 179:21]
  wire  btb_reset; // @[Frontend.scala 179:21]
  wire [38:0] btb_io_req_bits_addr; // @[Frontend.scala 179:21]
  wire  btb_io_resp_valid; // @[Frontend.scala 179:21]
  wire  btb_io_resp_bits_taken; // @[Frontend.scala 179:21]
  wire  btb_io_resp_bits_bridx; // @[Frontend.scala 179:21]
  wire [38:0] btb_io_resp_bits_target; // @[Frontend.scala 179:21]
  wire [4:0] btb_io_resp_bits_entry; // @[Frontend.scala 179:21]
  wire [7:0] btb_io_resp_bits_bht_history; // @[Frontend.scala 179:21]
  wire  btb_io_resp_bits_bht_value; // @[Frontend.scala 179:21]
  wire  btb_io_btb_update_valid; // @[Frontend.scala 179:21]
  wire [4:0] btb_io_btb_update_bits_prediction_entry; // @[Frontend.scala 179:21]
  wire [38:0] btb_io_btb_update_bits_pc; // @[Frontend.scala 179:21]
  wire  btb_io_btb_update_bits_isValid; // @[Frontend.scala 179:21]
  wire [38:0] btb_io_btb_update_bits_br_pc; // @[Frontend.scala 179:21]
  wire [1:0] btb_io_btb_update_bits_cfiType; // @[Frontend.scala 179:21]
  wire  btb_io_bht_update_valid; // @[Frontend.scala 179:21]
  wire [7:0] btb_io_bht_update_bits_prediction_history; // @[Frontend.scala 179:21]
  wire [38:0] btb_io_bht_update_bits_pc; // @[Frontend.scala 179:21]
  wire  btb_io_bht_update_bits_branch; // @[Frontend.scala 179:21]
  wire  btb_io_bht_update_bits_taken; // @[Frontend.scala 179:21]
  wire  btb_io_bht_update_bits_mispredict; // @[Frontend.scala 179:21]
  wire  btb_io_bht_advance_valid; // @[Frontend.scala 179:21]
  wire  btb_io_bht_advance_bits_bht_value; // @[Frontend.scala 179:21]
  wire  btb_io_ras_update_valid; // @[Frontend.scala 179:21]
  wire [1:0] btb_io_ras_update_bits_cfiType; // @[Frontend.scala 179:21]
  wire [38:0] btb_io_ras_update_bits_returnAddr; // @[Frontend.scala 179:21]
  wire  btb_io_ras_head_valid; // @[Frontend.scala 179:21]
  wire [38:0] btb_io_ras_head_bits; // @[Frontend.scala 179:21]
  wire  btb_io_flush; // @[Frontend.scala 179:21]
  wire [29:0] btb_io_covSum; // @[Frontend.scala 179:21]
  wire  btb_metaAssert; // @[Frontend.scala 179:21]
  wire  btb_metaReset; // @[Frontend.scala 179:21]
  wire  _T_2; // @[Frontend.scala 89:29]
  wire  _T_3; // @[Frontend.scala 89:52]
  wire  _T_4; // @[Frontend.scala 89:75]
  wire  _T_5; // @[Frontend.scala 89:102]
  wire  _T_7; // @[Frontend.scala 89:130]
  wire  _T_9; // @[Frontend.scala 89:9]
  reg  s1_valid; // @[Frontend.scala 100:21]
  reg [31:0] _RAND_0;
  reg  s2_valid; // @[Frontend.scala 101:25]
  reg [31:0] _RAND_1;
  wire  _s0_fq_has_space_T_6; // @[Frontend.scala 104:55]
  wire  _s0_fq_has_space_T_7; // @[Frontend.scala 104:41]
  wire  _s0_fq_has_space_T_8; // @[Frontend.scala 103:40]
  wire  _s0_fq_has_space_T_13; // @[Frontend.scala 105:55]
  wire  _s0_fq_has_space_T_14; // @[Frontend.scala 105:41]
  wire  s0_fq_has_space; // @[Frontend.scala 104:70]
  wire  s0_valid; // @[Frontend.scala 106:35]
  reg [39:0] s1_pc; // @[Frontend.scala 108:18]
  reg [63:0] _RAND_2;
  reg  s1_speculative; // @[Frontend.scala 109:27]
  reg [31:0] _RAND_3;
  wire [31:0] _s2_pc_T_1; // @[Frontend.scala 341:33]
  reg [39:0] s2_pc; // @[Frontend.scala 110:22]
  reg [63:0] _RAND_4;
  reg  s2_btb_resp_valid; // @[Frontend.scala 111:44]
  reg [31:0] _RAND_5;
  reg  s2_btb_resp_bits_taken; // @[Frontend.scala 112:29]
  reg [31:0] _RAND_6;
  reg  s2_btb_resp_bits_bridx; // @[Frontend.scala 112:29]
  reg [31:0] _RAND_7;
  reg [4:0] s2_btb_resp_bits_entry; // @[Frontend.scala 112:29]
  reg [31:0] _RAND_8;
  reg [7:0] s2_btb_resp_bits_bht_history; // @[Frontend.scala 112:29]
  reg [31:0] _RAND_9;
  reg  s2_btb_resp_bits_bht_value; // @[Frontend.scala 112:29]
  reg [31:0] _RAND_10;
  wire  s2_btb_taken; // @[Frontend.scala 113:40]
  reg  s2_tlb_resp_miss; // @[Frontend.scala 114:24]
  reg [31:0] _RAND_11;
  reg  s2_tlb_resp_pf_inst; // @[Frontend.scala 114:24]
  reg [31:0] _RAND_12;
  reg  s2_tlb_resp_ae_inst; // @[Frontend.scala 114:24]
  reg [31:0] _RAND_13;
  reg  s2_tlb_resp_cacheable; // @[Frontend.scala 114:24]
  reg [31:0] _RAND_14;
  wire  s2_xcpt; // @[Frontend.scala 115:37]
  reg  s2_speculative; // @[Frontend.scala 116:27]
  reg [31:0] _RAND_15;
  reg  s2_partial_insn_valid; // @[Frontend.scala 117:38]
  reg [31:0] _RAND_16;
  reg [15:0] s2_partial_insn; // @[Frontend.scala 118:28]
  reg [31:0] _RAND_17;
  reg  wrong_path; // @[Frontend.scala 119:27]
  reg [31:0] _RAND_18;
  wire [39:0] _s1_base_pc_T_1; // @[Frontend.scala 121:29]
  wire [39:0] s1_base_pc; // @[Frontend.scala 121:20]
  wire [39:0] ntpc; // @[Frontend.scala 122:25]
  wire  _s2_replay_T; // @[Decoupled.scala 40:37]
  wire  _s2_replay_T_2; // @[Frontend.scala 127:26]
  reg  s2_replay_REG; // @[Frontend.scala 127:58]
  reg [31:0] _RAND_19;
  wire  s2_replay; // @[Frontend.scala 127:48]
  wire  _s2_replay_T_4; // @[Frontend.scala 127:69]
  wire  _taken_prevRVI_T_1; // @[Frontend.scala 208:45]
  wire  taken_prevRVI; // @[Frontend.scala 209:31]
  wire [15:0] taken_bits; // @[Frontend.scala 211:37]
  wire [31:0] taken_rviBits; // @[Cat.scala 30:58]
  wire  taken_rviJump; // @[Frontend.scala 215:34]
  wire  taken_rviJALR; // @[Frontend.scala 216:34]
  wire  _taken_taken_T; // @[Frontend.scala 230:29]
  wire  taken_rviBranch; // @[Frontend.scala 214:36]
  wire  _taken_taken_T_1; // @[Frontend.scala 230:53]
  wire  _taken_taken_T_2; // @[Frontend.scala 230:40]
  wire  _taken_taken_T_3; // @[Frontend.scala 230:17]
  wire  taken_valid; // @[Frontend.scala 210:44]
  wire [15:0] _taken_rvcJump_T; // @[Frontend.scala 221:26]
  wire  taken_rvcJump; // @[Frontend.scala 221:26]
  wire [15:0] _taken_rvcJALR_T; // @[Frontend.scala 225:26]
  wire  _taken_rvcJALR_T_1; // @[Frontend.scala 225:26]
  wire  _taken_rvcJALR_T_3; // @[Frontend.scala 225:62]
  wire  taken_rvcJALR; // @[Frontend.scala 225:49]
  wire  _taken_taken_T_4; // @[Frontend.scala 231:27]
  wire  _taken_rvcJR_T_1; // @[Frontend.scala 223:24]
  wire  taken_rvcJR; // @[Frontend.scala 223:46]
  wire  _taken_taken_T_5; // @[Frontend.scala 231:38]
  wire  _taken_rvcBranch_T_1; // @[Frontend.scala 219:28]
  wire  _taken_rvcBranch_T_3; // @[Frontend.scala 219:60]
  wire  taken_rvcBranch; // @[Frontend.scala 219:52]
  wire  _taken_taken_T_6; // @[Frontend.scala 231:60]
  wire  _taken_taken_T_7; // @[Frontend.scala 231:47]
  wire  _taken_taken_T_8; // @[Frontend.scala 231:15]
  wire  taken_taken; // @[Frontend.scala 230:71]
  wire  taken_idx; // @[Frontend.scala 245:13]
  wire  _taken_prevRVI_T_4; // @[Frontend.scala 208:45]
  wire  taken_prevRVI_1; // @[Frontend.scala 209:31]
  wire [15:0] taken_bits_1; // @[Frontend.scala 211:37]
  wire [31:0] taken_rviBits_1; // @[Cat.scala 30:58]
  wire  taken_rviJALR_1; // @[Frontend.scala 216:34]
  wire  _taken_rviReturn_T_8; // @[Frontend.scala 217:31]
  wire [4:0] _taken_rviReturn_T_10; // @[Frontend.scala 217:66]
  wire  _taken_rviReturn_T_11; // @[Frontend.scala 217:66]
  wire  taken_rviReturn_1; // @[Frontend.scala 217:46]
  wire  _taken_predictReturn_T_3; // @[Frontend.scala 232:61]
  wire  taken_valid_1; // @[Frontend.scala 210:44]
  wire [15:0] _taken_rvcJR_T_4; // @[Frontend.scala 223:24]
  wire  _taken_rvcJR_T_5; // @[Frontend.scala 223:24]
  wire  _taken_rvcJR_T_7; // @[Frontend.scala 223:59]
  wire  taken_rvcJR_1; // @[Frontend.scala 223:46]
  wire [4:0] _taken_rvcReturn_T_4; // @[Frontend.scala 224:49]
  wire  _taken_rvcReturn_T_5; // @[Frontend.scala 224:49]
  wire  taken_rvcReturn_1; // @[Frontend.scala 224:29]
  wire  _taken_predictReturn_T_4; // @[Frontend.scala 232:83]
  wire  _taken_predictReturn_T_5; // @[Frontend.scala 232:74]
  wire  taken_predictReturn_1; // @[Frontend.scala 232:49]
  wire  _taken_T_45; // @[Frontend.scala 258:26]
  wire  _taken_rviReturn_T_2; // @[Frontend.scala 217:31]
  wire [4:0] _taken_rviReturn_T_4; // @[Frontend.scala 217:66]
  wire  _taken_rviReturn_T_5; // @[Frontend.scala 217:66]
  wire  taken_rviReturn; // @[Frontend.scala 217:46]
  wire  _taken_predictReturn_T; // @[Frontend.scala 232:61]
  wire [4:0] _taken_rvcReturn_T_1; // @[Frontend.scala 224:49]
  wire  _taken_rvcReturn_T_2; // @[Frontend.scala 224:49]
  wire  taken_rvcReturn; // @[Frontend.scala 224:29]
  wire  _taken_predictReturn_T_1; // @[Frontend.scala 232:83]
  wire  _taken_predictReturn_T_2; // @[Frontend.scala 232:74]
  wire  taken_predictReturn; // @[Frontend.scala 232:49]
  wire  _taken_T_16; // @[Frontend.scala 258:26]
  wire  _GEN_45; // @[Frontend.scala 254:30]
  wire  _GEN_78; // @[Frontend.scala 258:44]
  wire  _GEN_81; // @[Frontend.scala 254:30]
  wire  useRAS; // @[Frontend.scala 245:25]
  wire  taken_rviBranch_1; // @[Frontend.scala 214:36]
  wire  _taken_predictBranch_T_3; // @[Frontend.scala 234:53]
  wire [15:0] _taken_rvcBranch_T_4; // @[Frontend.scala 219:28]
  wire  _taken_rvcBranch_T_5; // @[Frontend.scala 219:28]
  wire  _taken_rvcBranch_T_7; // @[Frontend.scala 219:60]
  wire  taken_rvcBranch_1; // @[Frontend.scala 219:52]
  wire  _taken_predictBranch_T_4; // @[Frontend.scala 234:75]
  wire  _taken_predictBranch_T_5; // @[Frontend.scala 234:66]
  wire  taken_predictBranch_1; // @[Frontend.scala 234:41]
  wire  taken_rviJump_1; // @[Frontend.scala 215:34]
  wire  _taken_predictJump_T_2; // @[Frontend.scala 233:33]
  wire  taken_rvcJump_1; // @[Frontend.scala 221:26]
  wire  _taken_predictJump_T_3; // @[Frontend.scala 233:53]
  wire  taken_predictJump_1; // @[Frontend.scala 233:44]
  wire  _taken_T_46; // @[Frontend.scala 261:44]
  wire  _taken_T_47; // @[Frontend.scala 261:26]
  wire [39:0] _s2_base_pc_T_1; // @[Frontend.scala 201:31]
  wire [39:0] s2_base_pc; // @[Frontend.scala 201:22]
  wire [39:0] taken_pc_1; // @[Frontend.scala 262:33]
  wire [39:0] _taken_npc_T_6; // @[Frontend.scala 265:36]
  wire [39:0] _taken_npc_T_8; // @[Frontend.scala 265:57]
  wire  taken_rviImm_sign_2; // @[RocketCore.scala 1037:53]
  wire  taken_rviImm_hi_hi_hi_2; // @[Cat.scala 30:58]
  wire [10:0] taken_rviImm_hi_hi_lo_2; // @[Cat.scala 30:58]
  wire [7:0] taken_rviImm_hi_lo_hi_2; // @[Cat.scala 30:58]
  wire  taken_rviImm_hi_lo_lo_2; // @[Cat.scala 30:58]
  wire [5:0] taken_rviImm_lo_hi_hi_2; // @[RocketCore.scala 1043:66]
  wire [3:0] taken_rviImm_lo_hi_lo_2; // @[RocketCore.scala 1046:52]
  wire [31:0] _taken_rviImm_T_7; // @[RocketCore.scala 1051:53]
  wire [7:0] taken_rviImm_hi_lo_hi_3; // @[Cat.scala 30:58]
  wire  taken_rviImm_hi_lo_lo_3; // @[Cat.scala 30:58]
  wire [31:0] _taken_rviImm_T_9; // @[RocketCore.scala 1051:53]
  wire [31:0] taken_rviImm_1; // @[Frontend.scala 227:23]
  wire [4:0] taken_rvcImm_hi_hi_hi_2; // @[Bitwise.scala 72:12]
  wire [1:0] taken_rvcImm_hi_hi_lo_2; // @[RVC.scala 45:35]
  wire  taken_rvcImm_hi_lo_2; // @[RVC.scala 45:43]
  wire [1:0] taken_rvcImm_lo_hi_hi_2; // @[RVC.scala 45:49]
  wire [1:0] taken_rvcImm_lo_hi_lo_2; // @[RVC.scala 45:59]
  wire [12:0] _taken_rvcImm_T_13; // @[Frontend.scala 222:66]
  wire [9:0] taken_rvcImm_hi_hi_hi_hi_1; // @[Bitwise.scala 72:12]
  wire  taken_rvcImm_hi_hi_hi_lo_1; // @[RVC.scala 44:36]
  wire [1:0] taken_rvcImm_hi_hi_lo_3; // @[RVC.scala 44:42]
  wire  taken_rvcImm_hi_lo_hi_1; // @[RVC.scala 44:51]
  wire  taken_rvcImm_hi_lo_lo_1; // @[RVC.scala 44:57]
  wire  taken_rvcImm_lo_hi_lo_3; // @[RVC.scala 44:69]
  wire [2:0] taken_rvcImm_lo_lo_hi_1; // @[RVC.scala 44:76]
  wire [20:0] _taken_rvcImm_T_17; // @[Frontend.scala 222:106]
  wire [20:0] taken_rvcImm_1; // @[Frontend.scala 222:23]
  wire [31:0] _taken_npc_T_9; // @[Frontend.scala 265:69]
  wire [39:0] _GEN_127; // @[Frontend.scala 265:64]
  wire [39:0] _taken_predicted_npc_T_1; // @[Frontend.scala 266:34]
  wire  _taken_predictBranch_T; // @[Frontend.scala 234:53]
  wire  _taken_predictBranch_T_1; // @[Frontend.scala 234:75]
  wire  _taken_predictBranch_T_2; // @[Frontend.scala 234:66]
  wire  taken_predictBranch; // @[Frontend.scala 234:41]
  wire  _taken_predictJump_T; // @[Frontend.scala 233:33]
  wire  _taken_predictJump_T_1; // @[Frontend.scala 233:53]
  wire  taken_predictJump; // @[Frontend.scala 233:44]
  wire  _taken_T_17; // @[Frontend.scala 261:44]
  wire  _taken_T_18; // @[Frontend.scala 261:26]
  wire [39:0] _taken_npc_T; // @[Frontend.scala 264:32]
  wire  taken_rviImm_sign; // @[RocketCore.scala 1037:53]
  wire  taken_rviImm_hi_hi_hi; // @[Cat.scala 30:58]
  wire [10:0] taken_rviImm_hi_hi_lo; // @[Cat.scala 30:58]
  wire [7:0] taken_rviImm_hi_lo_hi; // @[Cat.scala 30:58]
  wire  taken_rviImm_hi_lo_lo; // @[Cat.scala 30:58]
  wire [5:0] taken_rviImm_lo_hi_hi; // @[RocketCore.scala 1043:66]
  wire [3:0] taken_rviImm_lo_hi_lo; // @[RocketCore.scala 1046:52]
  wire [31:0] _taken_rviImm_T_2; // @[RocketCore.scala 1051:53]
  wire [7:0] taken_rviImm_hi_lo_hi_1; // @[Cat.scala 30:58]
  wire  taken_rviImm_hi_lo_lo_1; // @[Cat.scala 30:58]
  wire [31:0] _taken_rviImm_T_4; // @[RocketCore.scala 1051:53]
  wire [31:0] taken_rviImm; // @[Frontend.scala 227:23]
  wire [32:0] _taken_npc_T_1; // @[Frontend.scala 264:61]
  wire [4:0] taken_rvcImm_hi_hi_hi; // @[Bitwise.scala 72:12]
  wire [1:0] taken_rvcImm_hi_hi_lo; // @[RVC.scala 45:35]
  wire  taken_rvcImm_hi_lo; // @[RVC.scala 45:43]
  wire [1:0] taken_rvcImm_lo_hi_hi; // @[RVC.scala 45:49]
  wire [1:0] taken_rvcImm_lo_hi_lo; // @[RVC.scala 45:59]
  wire [12:0] _taken_rvcImm_T_4; // @[Frontend.scala 222:66]
  wire [9:0] taken_rvcImm_hi_hi_hi_hi; // @[Bitwise.scala 72:12]
  wire  taken_rvcImm_hi_hi_hi_lo; // @[RVC.scala 44:36]
  wire [1:0] taken_rvcImm_hi_hi_lo_1; // @[RVC.scala 44:42]
  wire  taken_rvcImm_hi_lo_hi; // @[RVC.scala 44:51]
  wire  taken_rvcImm_hi_lo_lo; // @[RVC.scala 44:57]
  wire  taken_rvcImm_lo_hi_lo_1; // @[RVC.scala 44:69]
  wire [2:0] taken_rvcImm_lo_lo_hi; // @[RVC.scala 44:76]
  wire [20:0] _taken_rvcImm_T_8; // @[Frontend.scala 222:106]
  wire [20:0] taken_rvcImm; // @[Frontend.scala 222:23]
  wire [32:0] _taken_npc_T_2; // @[Frontend.scala 264:44]
  wire [39:0] _GEN_128; // @[Frontend.scala 264:39]
  wire [39:0] _taken_predicted_npc_T; // @[Frontend.scala 266:34]
  wire  predicted_taken; // @[Frontend.scala 192:29]
  wire  predicted_npc_hi; // @[package.scala 123:38]
  wire [39:0] _predicted_npc_T; // @[Cat.scala 30:58]
  wire [39:0] _GEN_28; // @[Frontend.scala 192:56]
  wire [39:0] _GEN_43; // @[Frontend.scala 261:61]
  wire [39:0] _GEN_46; // @[Frontend.scala 254:30]
  wire [39:0] _GEN_79; // @[Frontend.scala 261:61]
  wire [39:0] _GEN_82; // @[Frontend.scala 254:30]
  wire [39:0] _GEN_99; // @[Frontend.scala 245:25]
  wire [39:0] predicted_npc; // @[Frontend.scala 305:19]
  wire [39:0] npc; // @[Frontend.scala 128:16]
  wire  _s0_speculative_T_1; // @[Frontend.scala 134:53]
  wire  _s0_speculative_T_2; // @[Frontend.scala 134:41]
  wire  s0_speculative; // @[Frontend.scala 134:72]
  wire  _taken_taken_T_9; // @[Frontend.scala 230:29]
  wire  _taken_taken_T_10; // @[Frontend.scala 230:53]
  wire  _taken_taken_T_11; // @[Frontend.scala 230:40]
  wire  _taken_taken_T_12; // @[Frontend.scala 230:17]
  wire  _taken_rvcJALR_T_5; // @[Frontend.scala 225:26]
  wire  taken_rvcJALR_1; // @[Frontend.scala 225:49]
  wire  _taken_taken_T_13; // @[Frontend.scala 231:27]
  wire  _taken_taken_T_14; // @[Frontend.scala 231:38]
  wire  _taken_taken_T_15; // @[Frontend.scala 231:60]
  wire  _taken_taken_T_16; // @[Frontend.scala 231:47]
  wire  _taken_taken_T_17; // @[Frontend.scala 231:15]
  wire  taken_taken_1; // @[Frontend.scala 230:71]
  wire  taken; // @[Frontend.scala 286:19]
  wire  _GEN_116; // @[Frontend.scala 316:33]
  wire  _GEN_120; // @[Frontend.scala 312:20]
  wire  s2_redirect; // @[Frontend.scala 311:26]
  wire  _GEN_0; // @[Frontend.scala 140:21]
  wire  _icache_io_s1_kill_T; // @[Frontend.scala 160:36]
  wire  s2_can_speculatively_refill; // @[Frontend.scala 161:59]
  wire  _icache_io_s2_kill_T_1; // @[Frontend.scala 162:39]
  reg  fq_io_enq_valid_REG; // @[Frontend.scala 165:29]
  reg [31:0] _RAND_20;
  wire  _fq_io_enq_valid_T; // @[Frontend.scala 165:40]
  wire  _fq_io_enq_valid_T_2; // @[Frontend.scala 165:98]
  wire  _fq_io_enq_valid_T_3; // @[Frontend.scala 165:77]
  wire [39:0] _io_cpu_npc_T; // @[Frontend.scala 167:28]
  wire [39:0] _io_cpu_npc_T_2; // @[Frontend.scala 341:33]
  wire [2:0] _fq_io_enq_bits_mask_T_1; // @[Frontend.scala 170:52]
  wire  _fq_io_enq_bits_replay_T_1; // @[Frontend.scala 171:76]
  wire  _fq_io_enq_bits_replay_T_3; // @[Frontend.scala 171:101]
  wire  _fq_io_enq_bits_replay_T_4; // @[Frontend.scala 171:55]
  wire  _T_13; // @[Frontend.scala 175:27]
  wire  _T_15; // @[Frontend.scala 175:110]
  wire  _T_18; // @[Frontend.scala 175:9]
  wire  _T_20; // @[Frontend.scala 176:30]
  wire  fetch_bubble_likely; // @[Frontend.scala 293:33]
  wire  _btb_io_btb_update_valid_T_2; // @[Frontend.scala 294:51]
  wire  _btb_io_btb_update_valid_T_3; // @[Frontend.scala 294:66]
  wire  _taken_T_53; // @[Frontend.scala 273:52]
  wire  _taken_T_54; // @[Frontend.scala 273:91]
  wire  _taken_T_55; // @[Frontend.scala 273:106]
  wire  _taken_T_56; // @[Frontend.scala 273:34]
  wire  _taken_T_24; // @[Frontend.scala 273:52]
  wire  _taken_T_25; // @[Frontend.scala 273:91]
  wire  _taken_T_26; // @[Frontend.scala 273:106]
  wire  _taken_T_27; // @[Frontend.scala 273:34]
  wire  _GEN_92; // @[Frontend.scala 273:125]
  wire  updateBTB; // @[Frontend.scala 245:25]
  wire  _btb_io_btb_update_valid_T_4; // @[Frontend.scala 294:89]
  wire [1:0] _btb_io_btb_update_bits_br_pc_T; // @[Frontend.scala 298:63]
  wire [39:0] _GEN_129; // @[Frontend.scala 298:50]
  wire [39:0] _btb_io_btb_update_bits_br_pc_T_1; // @[Frontend.scala 298:50]
  wire [39:0] _GEN_36; // @[Frontend.scala 292:37]
  wire [39:0] _GEN_37; // @[Frontend.scala 292:37]
  wire [1:0] after_idx; // @[Frontend.scala 245:25]
  wire [2:0] _btb_io_ras_update_bits_returnAddr_T; // @[Frontend.scala 302:66]
  wire [39:0] _GEN_130; // @[Frontend.scala 302:53]
  wire [39:0] _btb_io_ras_update_bits_returnAddr_T_2; // @[Frontend.scala 302:53]
  wire  _taken_rviCall_T; // @[Frontend.scala 218:30]
  wire  taken_rviCall; // @[Frontend.scala 218:42]
  wire  _taken_T; // @[Frontend.scala 236:22]
  wire  _taken_T_2; // @[Frontend.scala 236:43]
  wire  _taken_T_3; // @[Frontend.scala 236:77]
  wire  _taken_T_5; // @[Frontend.scala 236:86]
  wire  _GEN_39; // @[Frontend.scala 236:95]
  wire  _GEN_40; // @[Frontend.scala 236:95]
  wire  _taken_btb_io_ras_update_valid_T_3; // @[Frontend.scala 248:92]
  wire  _taken_btb_io_ras_update_valid_T_4; // @[Frontend.scala 248:80]
  wire  _taken_btb_io_ras_update_valid_T_5; // @[Frontend.scala 248:127]
  wire  _taken_btb_io_ras_update_valid_T_6; // @[Frontend.scala 248:115]
  wire  _taken_btb_io_ras_update_valid_T_7; // @[Frontend.scala 248:106]
  wire  _taken_btb_io_ras_update_valid_T_8; // @[Frontend.scala 248:68]
  wire  _taken_btb_io_ras_update_bits_cfiType_T; // @[Frontend.scala 249:50]
  wire  _taken_btb_io_ras_update_bits_cfiType_T_1; // @[Frontend.scala 250:50]
  wire  _taken_btb_io_ras_update_bits_cfiType_T_2; // @[Frontend.scala 251:50]
  wire  _taken_btb_io_ras_update_bits_cfiType_T_5; // @[Frontend.scala 251:46]
  wire [1:0] _taken_btb_io_ras_update_bits_cfiType_T_6; // @[Frontend.scala 250:46]
  wire [1:0] _taken_btb_io_ras_update_bits_cfiType_T_7; // @[Frontend.scala 249:46]
  wire  _taken_T_9; // @[Frontend.scala 255:34]
  wire  _taken_T_11; // @[Frontend.scala 255:43]
  wire  _taken_T_13; // @[Frontend.scala 255:61]
  wire  _taken_T_15; // @[Frontend.scala 255:77]
  wire  _GEN_41; // @[Frontend.scala 255:96]
  wire  _GEN_44; // @[Frontend.scala 254:30]
  wire  _GEN_47; // @[Frontend.scala 269:59]
  wire  taken_rvc_1; // @[Frontend.scala 208:45]
  wire  _taken_rviCall_T_2; // @[Frontend.scala 218:30]
  wire  taken_rviCall_1; // @[Frontend.scala 218:42]
  wire  _taken_T_31; // @[Frontend.scala 236:43]
  wire  _taken_T_32; // @[Frontend.scala 236:77]
  wire  _taken_T_34; // @[Frontend.scala 236:86]
  wire  _GEN_76; // @[Frontend.scala 236:95]
  wire  _taken_btb_io_ras_update_valid_T_12; // @[Frontend.scala 248:92]
  wire  _taken_btb_io_ras_update_valid_T_13; // @[Frontend.scala 248:80]
  wire  _taken_btb_io_ras_update_valid_T_14; // @[Frontend.scala 248:127]
  wire  _taken_btb_io_ras_update_valid_T_15; // @[Frontend.scala 248:115]
  wire  _taken_btb_io_ras_update_valid_T_16; // @[Frontend.scala 248:106]
  wire  _taken_btb_io_ras_update_valid_T_17; // @[Frontend.scala 248:68]
  wire  _taken_btb_io_ras_update_bits_cfiType_T_8; // @[Frontend.scala 249:50]
  wire  _taken_btb_io_ras_update_bits_cfiType_T_9; // @[Frontend.scala 250:50]
  wire  _taken_btb_io_ras_update_bits_cfiType_T_10; // @[Frontend.scala 251:50]
  wire  _taken_btb_io_ras_update_bits_cfiType_T_13; // @[Frontend.scala 251:46]
  wire [1:0] _taken_btb_io_ras_update_bits_cfiType_T_14; // @[Frontend.scala 250:46]
  wire [1:0] _taken_btb_io_ras_update_bits_cfiType_T_15; // @[Frontend.scala 249:46]
  wire  _taken_T_38; // @[Frontend.scala 255:34]
  wire  _taken_T_40; // @[Frontend.scala 255:43]
  wire  _taken_T_42; // @[Frontend.scala 255:61]
  wire  _taken_T_44; // @[Frontend.scala 255:77]
  wire  _GEN_77; // @[Frontend.scala 255:96]
  wire  _GEN_83; // @[Frontend.scala 269:59]
  wire  _taken_T_59; // @[Frontend.scala 281:23]
  wire  _taken_T_61; // @[Frontend.scala 281:37]
  wire [15:0] _taken_lo_T; // @[Frontend.scala 283:37]
  wire  _T_25; // @[Frontend.scala 308:45]
  wire  _T_26; // @[Frontend.scala 308:28]
  wire  _GEN_117; // @[Frontend.scala 312:20]
  wire  _GEN_118; // @[Frontend.scala 312:20]
  wire [4:0] _GEN_119; // @[Frontend.scala 312:20]
  wire  _T_31; // @[Frontend.scala 320:35]
  wire  _T_33; // @[Frontend.scala 320:11]
  reg [5:0] Frontend_state; // @[Register tracking Frontend state]
  reg [31:0] _RAND_21;
  reg  Frontend_cov [0:63]; // @[Coverage map for Frontend]
  reg [31:0] _RAND_22;
  wire  Frontend_cov_read_data; // @[Coverage map for Frontend]
  wire [5:0] Frontend_cov_read_addr; // @[Coverage map for Frontend]
  wire  Frontend_cov_write_data; // @[Coverage map for Frontend]
  wire [5:0] Frontend_cov_write_addr; // @[Coverage map for Frontend]
  wire  Frontend_cov_write_mask; // @[Coverage map for Frontend]
  wire  Frontend_cov_write_en; // @[Coverage map for Frontend]
  reg [29:0] Frontend_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_23;
  wire  s2_partial_insn_valid_shl;
  wire [5:0] s2_partial_insn_valid_pad;
  wire [1:0] s2_btb_resp_valid_shl;
  wire [5:0] s2_btb_resp_valid_pad;
  wire [2:0] s2_replay_REG_shl;
  wire [5:0] s2_replay_REG_pad;
  wire [3:0] s2_btb_resp_bits_bht_value_shl;
  wire [5:0] s2_btb_resp_bits_bht_value_pad;
  wire [4:0] s2_valid_shl;
  wire [5:0] s2_valid_pad;
  wire [5:0] s2_btb_resp_bits_taken_shl;
  wire [5:0] s2_btb_resp_bits_taken_pad;
  wire [5:0] Frontend_xor4;
  wire [5:0] Frontend_xor1;
  wire [5:0] Frontend_xor6;
  wire [5:0] Frontend_xor2;
  wire [5:0] Frontend_xor0;
  wire [29:0] icache_sum;
  wire [29:0] fq_sum;
  wire [29:0] tlb_sum;
  wire [29:0] btb_sum;
  wire  stopEn0;
  wire  stopEn1;
  wire  stopEn2;
  wire  icache_metaAssert_wire;
  wire  fq_metaAssert_wire;
  wire  tlb_metaAssert_wire;
  wire  btb_metaAssert_wire;
  wire  Frontend_or4;
  wire  Frontend_or1;
  wire  Frontend_or5;
  wire  Frontend_or6;
  wire  Frontend_or2;
  wire  Frontend_or0;
  ICache icache ( // @[Frontend.scala 62:26]
    .clock(icache_clock),
    .reset(icache_reset),
    .auto_master_out_a_ready(icache_auto_master_out_a_ready),
    .auto_master_out_a_valid(icache_auto_master_out_a_valid),
    .auto_master_out_a_bits_address(icache_auto_master_out_a_bits_address),
    .auto_master_out_d_valid(icache_auto_master_out_d_valid),
    .auto_master_out_d_bits_opcode(icache_auto_master_out_d_bits_opcode),
    .auto_master_out_d_bits_size(icache_auto_master_out_d_bits_size),
    .auto_master_out_d_bits_data(icache_auto_master_out_d_bits_data),
    .auto_master_out_d_bits_corrupt(icache_auto_master_out_d_bits_corrupt),
    .io_req_ready(icache_io_req_ready),
    .io_req_valid(icache_io_req_valid),
    .io_req_bits_addr(icache_io_req_bits_addr),
    .io_s1_paddr(icache_io_s1_paddr),
    .io_s1_kill(icache_io_s1_kill),
    .io_s2_kill(icache_io_s2_kill),
    .io_resp_valid(icache_io_resp_valid),
    .io_resp_bits_data(icache_io_resp_bits_data),
    .io_resp_bits_replay(icache_io_resp_bits_replay),
    .io_resp_bits_ae(icache_io_resp_bits_ae),
    .io_invalidate(icache_io_invalidate),
    .io_covSum(icache_io_covSum),
    .metaAssert(icache_metaAssert),
    .metaReset(icache_metaReset),
    .repl_way_v0_prng_halt(icache_repl_way_v0_prng_halt)
  );
  ShiftQueue fq ( // @[Frontend.scala 84:57]
    .clock(fq_clock),
    .reset(fq_reset),
    .io_enq_ready(fq_io_enq_ready),
    .io_enq_valid(fq_io_enq_valid),
    .io_enq_bits_btb_taken(fq_io_enq_bits_btb_taken),
    .io_enq_bits_btb_bridx(fq_io_enq_bits_btb_bridx),
    .io_enq_bits_btb_entry(fq_io_enq_bits_btb_entry),
    .io_enq_bits_btb_bht_history(fq_io_enq_bits_btb_bht_history),
    .io_enq_bits_pc(fq_io_enq_bits_pc),
    .io_enq_bits_data(fq_io_enq_bits_data),
    .io_enq_bits_mask(fq_io_enq_bits_mask),
    .io_enq_bits_xcpt_pf_inst(fq_io_enq_bits_xcpt_pf_inst),
    .io_enq_bits_xcpt_ae_inst(fq_io_enq_bits_xcpt_ae_inst),
    .io_enq_bits_replay(fq_io_enq_bits_replay),
    .io_deq_ready(fq_io_deq_ready),
    .io_deq_valid(fq_io_deq_valid),
    .io_deq_bits_btb_taken(fq_io_deq_bits_btb_taken),
    .io_deq_bits_btb_bridx(fq_io_deq_bits_btb_bridx),
    .io_deq_bits_btb_entry(fq_io_deq_bits_btb_entry),
    .io_deq_bits_btb_bht_history(fq_io_deq_bits_btb_bht_history),
    .io_deq_bits_pc(fq_io_deq_bits_pc),
    .io_deq_bits_data(fq_io_deq_bits_data),
    .io_deq_bits_xcpt_pf_inst(fq_io_deq_bits_xcpt_pf_inst),
    .io_deq_bits_xcpt_ae_inst(fq_io_deq_bits_xcpt_ae_inst),
    .io_deq_bits_replay(fq_io_deq_bits_replay),
    .io_mask(fq_io_mask),
    .io_covSum(fq_io_covSum),
    .metaAssert(fq_metaAssert),
    .metaReset(fq_metaReset)
  );
  TLB_1 tlb ( // @[Frontend.scala 98:19]
    .clock(tlb_clock),
    .reset(tlb_reset),
    .io_req_ready(tlb_io_req_ready),
    .io_req_valid(tlb_io_req_valid),
    .io_req_bits_vaddr(tlb_io_req_bits_vaddr),
    .io_resp_miss(tlb_io_resp_miss),
    .io_resp_paddr(tlb_io_resp_paddr),
    .io_resp_pf_inst(tlb_io_resp_pf_inst),
    .io_resp_ae_inst(tlb_io_resp_ae_inst),
    .io_resp_cacheable(tlb_io_resp_cacheable),
    .io_sfence_valid(tlb_io_sfence_valid),
    .io_sfence_bits_rs1(tlb_io_sfence_bits_rs1),
    .io_sfence_bits_rs2(tlb_io_sfence_bits_rs2),
    .io_sfence_bits_addr(tlb_io_sfence_bits_addr),
    .io_ptw_req_ready(tlb_io_ptw_req_ready),
    .io_ptw_req_valid(tlb_io_ptw_req_valid),
    .io_ptw_req_bits_valid(tlb_io_ptw_req_bits_valid),
    .io_ptw_req_bits_bits_addr(tlb_io_ptw_req_bits_bits_addr),
    .io_ptw_resp_valid(tlb_io_ptw_resp_valid),
    .io_ptw_resp_bits_ae(tlb_io_ptw_resp_bits_ae),
    .io_ptw_resp_bits_pte_ppn(tlb_io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_d(tlb_io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_a(tlb_io_ptw_resp_bits_pte_a),
    .io_ptw_resp_bits_pte_g(tlb_io_ptw_resp_bits_pte_g),
    .io_ptw_resp_bits_pte_u(tlb_io_ptw_resp_bits_pte_u),
    .io_ptw_resp_bits_pte_x(tlb_io_ptw_resp_bits_pte_x),
    .io_ptw_resp_bits_pte_w(tlb_io_ptw_resp_bits_pte_w),
    .io_ptw_resp_bits_pte_r(tlb_io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_v(tlb_io_ptw_resp_bits_pte_v),
    .io_ptw_resp_bits_level(tlb_io_ptw_resp_bits_level),
    .io_ptw_resp_bits_homogeneous(tlb_io_ptw_resp_bits_homogeneous),
    .io_ptw_ptbr_mode(tlb_io_ptw_ptbr_mode),
    .io_ptw_status_debug(tlb_io_ptw_status_debug),
    .io_ptw_status_prv(tlb_io_ptw_status_prv),
    .io_ptw_pmp_0_cfg_l(tlb_io_ptw_pmp_0_cfg_l),
    .io_ptw_pmp_0_cfg_a(tlb_io_ptw_pmp_0_cfg_a),
    .io_ptw_pmp_0_cfg_x(tlb_io_ptw_pmp_0_cfg_x),
    .io_ptw_pmp_0_cfg_w(tlb_io_ptw_pmp_0_cfg_w),
    .io_ptw_pmp_0_cfg_r(tlb_io_ptw_pmp_0_cfg_r),
    .io_ptw_pmp_0_addr(tlb_io_ptw_pmp_0_addr),
    .io_ptw_pmp_0_mask(tlb_io_ptw_pmp_0_mask),
    .io_ptw_pmp_1_cfg_l(tlb_io_ptw_pmp_1_cfg_l),
    .io_ptw_pmp_1_cfg_a(tlb_io_ptw_pmp_1_cfg_a),
    .io_ptw_pmp_1_cfg_x(tlb_io_ptw_pmp_1_cfg_x),
    .io_ptw_pmp_1_cfg_w(tlb_io_ptw_pmp_1_cfg_w),
    .io_ptw_pmp_1_cfg_r(tlb_io_ptw_pmp_1_cfg_r),
    .io_ptw_pmp_1_addr(tlb_io_ptw_pmp_1_addr),
    .io_ptw_pmp_1_mask(tlb_io_ptw_pmp_1_mask),
    .io_ptw_pmp_2_cfg_l(tlb_io_ptw_pmp_2_cfg_l),
    .io_ptw_pmp_2_cfg_a(tlb_io_ptw_pmp_2_cfg_a),
    .io_ptw_pmp_2_cfg_x(tlb_io_ptw_pmp_2_cfg_x),
    .io_ptw_pmp_2_cfg_w(tlb_io_ptw_pmp_2_cfg_w),
    .io_ptw_pmp_2_cfg_r(tlb_io_ptw_pmp_2_cfg_r),
    .io_ptw_pmp_2_addr(tlb_io_ptw_pmp_2_addr),
    .io_ptw_pmp_2_mask(tlb_io_ptw_pmp_2_mask),
    .io_ptw_pmp_3_cfg_l(tlb_io_ptw_pmp_3_cfg_l),
    .io_ptw_pmp_3_cfg_a(tlb_io_ptw_pmp_3_cfg_a),
    .io_ptw_pmp_3_cfg_x(tlb_io_ptw_pmp_3_cfg_x),
    .io_ptw_pmp_3_cfg_w(tlb_io_ptw_pmp_3_cfg_w),
    .io_ptw_pmp_3_cfg_r(tlb_io_ptw_pmp_3_cfg_r),
    .io_ptw_pmp_3_addr(tlb_io_ptw_pmp_3_addr),
    .io_ptw_pmp_3_mask(tlb_io_ptw_pmp_3_mask),
    .io_ptw_pmp_4_cfg_l(tlb_io_ptw_pmp_4_cfg_l),
    .io_ptw_pmp_4_cfg_a(tlb_io_ptw_pmp_4_cfg_a),
    .io_ptw_pmp_4_cfg_x(tlb_io_ptw_pmp_4_cfg_x),
    .io_ptw_pmp_4_cfg_w(tlb_io_ptw_pmp_4_cfg_w),
    .io_ptw_pmp_4_cfg_r(tlb_io_ptw_pmp_4_cfg_r),
    .io_ptw_pmp_4_addr(tlb_io_ptw_pmp_4_addr),
    .io_ptw_pmp_4_mask(tlb_io_ptw_pmp_4_mask),
    .io_ptw_pmp_5_cfg_l(tlb_io_ptw_pmp_5_cfg_l),
    .io_ptw_pmp_5_cfg_a(tlb_io_ptw_pmp_5_cfg_a),
    .io_ptw_pmp_5_cfg_x(tlb_io_ptw_pmp_5_cfg_x),
    .io_ptw_pmp_5_cfg_w(tlb_io_ptw_pmp_5_cfg_w),
    .io_ptw_pmp_5_cfg_r(tlb_io_ptw_pmp_5_cfg_r),
    .io_ptw_pmp_5_addr(tlb_io_ptw_pmp_5_addr),
    .io_ptw_pmp_5_mask(tlb_io_ptw_pmp_5_mask),
    .io_ptw_pmp_6_cfg_l(tlb_io_ptw_pmp_6_cfg_l),
    .io_ptw_pmp_6_cfg_a(tlb_io_ptw_pmp_6_cfg_a),
    .io_ptw_pmp_6_cfg_x(tlb_io_ptw_pmp_6_cfg_x),
    .io_ptw_pmp_6_cfg_w(tlb_io_ptw_pmp_6_cfg_w),
    .io_ptw_pmp_6_cfg_r(tlb_io_ptw_pmp_6_cfg_r),
    .io_ptw_pmp_6_addr(tlb_io_ptw_pmp_6_addr),
    .io_ptw_pmp_6_mask(tlb_io_ptw_pmp_6_mask),
    .io_ptw_pmp_7_cfg_l(tlb_io_ptw_pmp_7_cfg_l),
    .io_ptw_pmp_7_cfg_a(tlb_io_ptw_pmp_7_cfg_a),
    .io_ptw_pmp_7_cfg_x(tlb_io_ptw_pmp_7_cfg_x),
    .io_ptw_pmp_7_cfg_w(tlb_io_ptw_pmp_7_cfg_w),
    .io_ptw_pmp_7_cfg_r(tlb_io_ptw_pmp_7_cfg_r),
    .io_ptw_pmp_7_addr(tlb_io_ptw_pmp_7_addr),
    .io_ptw_pmp_7_mask(tlb_io_ptw_pmp_7_mask),
    .io_kill(tlb_io_kill),
    .io_covSum(tlb_io_covSum),
    .metaAssert(tlb_metaAssert),
    .metaReset(tlb_metaReset)
  );
  BTB btb ( // @[Frontend.scala 179:21]
    .clock(btb_clock),
    .reset(btb_reset),
    .io_req_bits_addr(btb_io_req_bits_addr),
    .io_resp_valid(btb_io_resp_valid),
    .io_resp_bits_taken(btb_io_resp_bits_taken),
    .io_resp_bits_bridx(btb_io_resp_bits_bridx),
    .io_resp_bits_target(btb_io_resp_bits_target),
    .io_resp_bits_entry(btb_io_resp_bits_entry),
    .io_resp_bits_bht_history(btb_io_resp_bits_bht_history),
    .io_resp_bits_bht_value(btb_io_resp_bits_bht_value),
    .io_btb_update_valid(btb_io_btb_update_valid),
    .io_btb_update_bits_prediction_entry(btb_io_btb_update_bits_prediction_entry),
    .io_btb_update_bits_pc(btb_io_btb_update_bits_pc),
    .io_btb_update_bits_isValid(btb_io_btb_update_bits_isValid),
    .io_btb_update_bits_br_pc(btb_io_btb_update_bits_br_pc),
    .io_btb_update_bits_cfiType(btb_io_btb_update_bits_cfiType),
    .io_bht_update_valid(btb_io_bht_update_valid),
    .io_bht_update_bits_prediction_history(btb_io_bht_update_bits_prediction_history),
    .io_bht_update_bits_pc(btb_io_bht_update_bits_pc),
    .io_bht_update_bits_branch(btb_io_bht_update_bits_branch),
    .io_bht_update_bits_taken(btb_io_bht_update_bits_taken),
    .io_bht_update_bits_mispredict(btb_io_bht_update_bits_mispredict),
    .io_bht_advance_valid(btb_io_bht_advance_valid),
    .io_bht_advance_bits_bht_value(btb_io_bht_advance_bits_bht_value),
    .io_ras_update_valid(btb_io_ras_update_valid),
    .io_ras_update_bits_cfiType(btb_io_ras_update_bits_cfiType),
    .io_ras_update_bits_returnAddr(btb_io_ras_update_bits_returnAddr),
    .io_ras_head_valid(btb_io_ras_head_valid),
    .io_ras_head_bits(btb_io_ras_head_bits),
    .io_flush(btb_io_flush),
    .io_covSum(btb_io_covSum),
    .metaAssert(btb_metaAssert),
    .metaReset(btb_metaReset)
  );
  assign _T_2 = io_cpu_req_valid | io_cpu_sfence_valid; // @[Frontend.scala 89:29]
  assign _T_3 = _T_2 | io_cpu_flush_icache; // @[Frontend.scala 89:52]
  assign _T_4 = _T_3 | io_cpu_bht_update_valid; // @[Frontend.scala 89:75]
  assign _T_5 = _T_4 | io_cpu_btb_update_valid; // @[Frontend.scala 89:102]
  assign _T_7 = ~_T_5 | io_cpu_might_request; // @[Frontend.scala 89:130]
  assign _T_9 = _T_7 | reset; // @[Frontend.scala 89:9]
  assign _s0_fq_has_space_T_6 = ~s1_valid | ~s2_valid; // @[Frontend.scala 104:55]
  assign _s0_fq_has_space_T_7 = ~fq_io_mask[3] & _s0_fq_has_space_T_6; // @[Frontend.scala 104:41]
  assign _s0_fq_has_space_T_8 = ~fq_io_mask[2] | _s0_fq_has_space_T_7; // @[Frontend.scala 103:40]
  assign _s0_fq_has_space_T_13 = ~s1_valid & ~s2_valid; // @[Frontend.scala 105:55]
  assign _s0_fq_has_space_T_14 = ~fq_io_mask[4] & _s0_fq_has_space_T_13; // @[Frontend.scala 105:41]
  assign s0_fq_has_space = _s0_fq_has_space_T_8 | _s0_fq_has_space_T_14; // @[Frontend.scala 104:70]
  assign s0_valid = io_cpu_req_valid | s0_fq_has_space; // @[Frontend.scala 106:35]
  assign _s2_pc_T_1 = ~auto_reset_vector_sink_in | 32'h1; // @[Frontend.scala 341:33]
  assign s2_btb_taken = s2_btb_resp_valid & s2_btb_resp_bits_taken; // @[Frontend.scala 113:40]
  assign s2_xcpt = s2_tlb_resp_ae_inst | s2_tlb_resp_pf_inst; // @[Frontend.scala 115:37]
  assign _s1_base_pc_T_1 = ~s1_pc | 40'h3; // @[Frontend.scala 121:29]
  assign s1_base_pc = ~_s1_base_pc_T_1; // @[Frontend.scala 121:20]
  assign ntpc = s1_base_pc + 40'h4; // @[Frontend.scala 122:25]
  assign _s2_replay_T = fq_io_enq_ready & fq_io_enq_valid; // @[Decoupled.scala 40:37]
  assign _s2_replay_T_2 = s2_valid & ~_s2_replay_T; // @[Frontend.scala 127:26]
  assign s2_replay = _s2_replay_T_2 | s2_replay_REG; // @[Frontend.scala 127:48]
  assign _s2_replay_T_4 = s2_replay & ~s0_valid; // @[Frontend.scala 127:69]
  assign _taken_prevRVI_T_1 = s2_partial_insn[1:0] != 2'h3; // @[Frontend.scala 208:45]
  assign taken_prevRVI = s2_partial_insn_valid & ~_taken_prevRVI_T_1; // @[Frontend.scala 209:31]
  assign taken_bits = fq_io_enq_bits_data[15:0]; // @[Frontend.scala 211:37]
  assign taken_rviBits = {taken_bits,s2_partial_insn}; // @[Cat.scala 30:58]
  assign taken_rviJump = taken_rviBits[6:0] == 7'h6f; // @[Frontend.scala 215:34]
  assign taken_rviJALR = taken_rviBits[6:0] == 7'h67; // @[Frontend.scala 216:34]
  assign _taken_taken_T = taken_rviJump | taken_rviJALR; // @[Frontend.scala 230:29]
  assign taken_rviBranch = taken_rviBits[6:0] == 7'h63; // @[Frontend.scala 214:36]
  assign _taken_taken_T_1 = taken_rviBranch & s2_btb_resp_bits_bht_value; // @[Frontend.scala 230:53]
  assign _taken_taken_T_2 = _taken_taken_T | _taken_taken_T_1; // @[Frontend.scala 230:40]
  assign _taken_taken_T_3 = taken_prevRVI & _taken_taken_T_2; // @[Frontend.scala 230:17]
  assign taken_valid = fq_io_enq_bits_mask[0] & ~taken_prevRVI; // @[Frontend.scala 210:44]
  assign _taken_rvcJump_T = taken_bits & 16'he003; // @[Frontend.scala 221:26]
  assign taken_rvcJump = 16'ha001 == _taken_rvcJump_T; // @[Frontend.scala 221:26]
  assign _taken_rvcJALR_T = taken_bits & 16'hf003; // @[Frontend.scala 225:26]
  assign _taken_rvcJALR_T_1 = 16'h9002 == _taken_rvcJALR_T; // @[Frontend.scala 225:26]
  assign _taken_rvcJALR_T_3 = taken_bits[6:2] == 5'h0; // @[Frontend.scala 225:62]
  assign taken_rvcJALR = _taken_rvcJALR_T_1 & _taken_rvcJALR_T_3; // @[Frontend.scala 225:49]
  assign _taken_taken_T_4 = taken_rvcJump | taken_rvcJALR; // @[Frontend.scala 231:27]
  assign _taken_rvcJR_T_1 = 16'h8002 == _taken_rvcJALR_T; // @[Frontend.scala 223:24]
  assign taken_rvcJR = _taken_rvcJR_T_1 & _taken_rvcJALR_T_3; // @[Frontend.scala 223:46]
  assign _taken_taken_T_5 = _taken_taken_T_4 | taken_rvcJR; // @[Frontend.scala 231:38]
  assign _taken_rvcBranch_T_1 = 16'hc001 == _taken_rvcJump_T; // @[Frontend.scala 219:28]
  assign _taken_rvcBranch_T_3 = 16'he001 == _taken_rvcJump_T; // @[Frontend.scala 219:60]
  assign taken_rvcBranch = _taken_rvcBranch_T_1 | _taken_rvcBranch_T_3; // @[Frontend.scala 219:52]
  assign _taken_taken_T_6 = taken_rvcBranch & s2_btb_resp_bits_bht_value; // @[Frontend.scala 231:60]
  assign _taken_taken_T_7 = _taken_taken_T_5 | _taken_taken_T_6; // @[Frontend.scala 231:47]
  assign _taken_taken_T_8 = taken_valid & _taken_taken_T_7; // @[Frontend.scala 231:15]
  assign taken_taken = _taken_taken_T_3 | _taken_taken_T_8; // @[Frontend.scala 230:71]
  assign taken_idx = ~taken_taken; // @[Frontend.scala 245:13]
  assign _taken_prevRVI_T_4 = taken_bits[1:0] != 2'h3; // @[Frontend.scala 208:45]
  assign taken_prevRVI_1 = taken_valid & ~_taken_prevRVI_T_4; // @[Frontend.scala 209:31]
  assign taken_bits_1 = fq_io_enq_bits_data[31:16]; // @[Frontend.scala 211:37]
  assign taken_rviBits_1 = {taken_bits_1,taken_bits}; // @[Cat.scala 30:58]
  assign taken_rviJALR_1 = taken_rviBits_1[6:0] == 7'h67; // @[Frontend.scala 216:34]
  assign _taken_rviReturn_T_8 = taken_rviJALR_1 & ~taken_rviBits_1[7]; // @[Frontend.scala 217:31]
  assign _taken_rviReturn_T_10 = taken_rviBits_1[19:15] & 5'h1b; // @[Frontend.scala 217:66]
  assign _taken_rviReturn_T_11 = 5'h1 == _taken_rviReturn_T_10; // @[Frontend.scala 217:66]
  assign taken_rviReturn_1 = _taken_rviReturn_T_8 & _taken_rviReturn_T_11; // @[Frontend.scala 217:46]
  assign _taken_predictReturn_T_3 = taken_prevRVI_1 & taken_rviReturn_1; // @[Frontend.scala 232:61]
  assign taken_valid_1 = fq_io_enq_bits_mask[1] & ~taken_prevRVI_1; // @[Frontend.scala 210:44]
  assign _taken_rvcJR_T_4 = taken_bits_1 & 16'hf003; // @[Frontend.scala 223:24]
  assign _taken_rvcJR_T_5 = 16'h8002 == _taken_rvcJR_T_4; // @[Frontend.scala 223:24]
  assign _taken_rvcJR_T_7 = taken_bits_1[6:2] == 5'h0; // @[Frontend.scala 223:59]
  assign taken_rvcJR_1 = _taken_rvcJR_T_5 & _taken_rvcJR_T_7; // @[Frontend.scala 223:46]
  assign _taken_rvcReturn_T_4 = taken_bits_1[11:7] & 5'h1b; // @[Frontend.scala 224:49]
  assign _taken_rvcReturn_T_5 = 5'h1 == _taken_rvcReturn_T_4; // @[Frontend.scala 224:49]
  assign taken_rvcReturn_1 = taken_rvcJR_1 & _taken_rvcReturn_T_5; // @[Frontend.scala 224:29]
  assign _taken_predictReturn_T_4 = taken_valid_1 & taken_rvcReturn_1; // @[Frontend.scala 232:83]
  assign _taken_predictReturn_T_5 = _taken_predictReturn_T_3 | _taken_predictReturn_T_4; // @[Frontend.scala 232:74]
  assign taken_predictReturn_1 = btb_io_ras_head_valid & _taken_predictReturn_T_5; // @[Frontend.scala 232:49]
  assign _taken_T_45 = s2_valid & taken_predictReturn_1; // @[Frontend.scala 258:26]
  assign _taken_rviReturn_T_2 = taken_rviJALR & ~taken_rviBits[7]; // @[Frontend.scala 217:31]
  assign _taken_rviReturn_T_4 = taken_rviBits[19:15] & 5'h1b; // @[Frontend.scala 217:66]
  assign _taken_rviReturn_T_5 = 5'h1 == _taken_rviReturn_T_4; // @[Frontend.scala 217:66]
  assign taken_rviReturn = _taken_rviReturn_T_2 & _taken_rviReturn_T_5; // @[Frontend.scala 217:46]
  assign _taken_predictReturn_T = taken_prevRVI & taken_rviReturn; // @[Frontend.scala 232:61]
  assign _taken_rvcReturn_T_1 = taken_bits[11:7] & 5'h1b; // @[Frontend.scala 224:49]
  assign _taken_rvcReturn_T_2 = 5'h1 == _taken_rvcReturn_T_1; // @[Frontend.scala 224:49]
  assign taken_rvcReturn = taken_rvcJR & _taken_rvcReturn_T_2; // @[Frontend.scala 224:29]
  assign _taken_predictReturn_T_1 = taken_valid & taken_rvcReturn; // @[Frontend.scala 232:83]
  assign _taken_predictReturn_T_2 = _taken_predictReturn_T | _taken_predictReturn_T_1; // @[Frontend.scala 232:74]
  assign taken_predictReturn = btb_io_ras_head_valid & _taken_predictReturn_T_2; // @[Frontend.scala 232:49]
  assign _taken_T_16 = s2_valid & taken_predictReturn; // @[Frontend.scala 258:26]
  assign _GEN_45 = ~s2_btb_taken & _taken_T_16; // @[Frontend.scala 254:30]
  assign _GEN_78 = _taken_T_45 | _GEN_45; // @[Frontend.scala 258:44]
  assign _GEN_81 = s2_btb_taken ? _GEN_45 : _GEN_78; // @[Frontend.scala 254:30]
  assign useRAS = taken_idx ? _GEN_81 : _GEN_45; // @[Frontend.scala 245:25]
  assign taken_rviBranch_1 = taken_rviBits_1[6:0] == 7'h63; // @[Frontend.scala 214:36]
  assign _taken_predictBranch_T_3 = taken_prevRVI_1 & taken_rviBranch_1; // @[Frontend.scala 234:53]
  assign _taken_rvcBranch_T_4 = taken_bits_1 & 16'he003; // @[Frontend.scala 219:28]
  assign _taken_rvcBranch_T_5 = 16'hc001 == _taken_rvcBranch_T_4; // @[Frontend.scala 219:28]
  assign _taken_rvcBranch_T_7 = 16'he001 == _taken_rvcBranch_T_4; // @[Frontend.scala 219:60]
  assign taken_rvcBranch_1 = _taken_rvcBranch_T_5 | _taken_rvcBranch_T_7; // @[Frontend.scala 219:52]
  assign _taken_predictBranch_T_4 = taken_valid_1 & taken_rvcBranch_1; // @[Frontend.scala 234:75]
  assign _taken_predictBranch_T_5 = _taken_predictBranch_T_3 | _taken_predictBranch_T_4; // @[Frontend.scala 234:66]
  assign taken_predictBranch_1 = s2_btb_resp_bits_bht_value & _taken_predictBranch_T_5; // @[Frontend.scala 234:41]
  assign taken_rviJump_1 = taken_rviBits_1[6:0] == 7'h6f; // @[Frontend.scala 215:34]
  assign _taken_predictJump_T_2 = taken_prevRVI_1 & taken_rviJump_1; // @[Frontend.scala 233:33]
  assign taken_rvcJump_1 = 16'ha001 == _taken_rvcBranch_T_4; // @[Frontend.scala 221:26]
  assign _taken_predictJump_T_3 = taken_valid_1 & taken_rvcJump_1; // @[Frontend.scala 233:53]
  assign taken_predictJump_1 = _taken_predictJump_T_2 | _taken_predictJump_T_3; // @[Frontend.scala 233:44]
  assign _taken_T_46 = taken_predictBranch_1 | taken_predictJump_1; // @[Frontend.scala 261:44]
  assign _taken_T_47 = s2_valid & _taken_T_46; // @[Frontend.scala 261:26]
  assign _s2_base_pc_T_1 = ~s2_pc | 40'h3; // @[Frontend.scala 201:31]
  assign s2_base_pc = ~_s2_base_pc_T_1; // @[Frontend.scala 201:22]
  assign taken_pc_1 = s2_base_pc | 40'h2; // @[Frontend.scala 262:33]
  assign _taken_npc_T_6 = taken_pc_1 - 40'h2; // @[Frontend.scala 265:36]
  assign _taken_npc_T_8 = taken_prevRVI_1 ? _taken_npc_T_6 : taken_pc_1; // @[Frontend.scala 265:57]
  assign taken_rviImm_sign_2 = taken_rviBits_1[31]; // @[RocketCore.scala 1037:53]
  assign taken_rviImm_hi_hi_hi_2 = taken_rviBits_1[31]; // @[Cat.scala 30:58]
  assign taken_rviImm_hi_hi_lo_2 = {11{taken_rviImm_sign_2}}; // @[Cat.scala 30:58]
  assign taken_rviImm_hi_lo_hi_2 = taken_rviBits_1[19:12]; // @[Cat.scala 30:58]
  assign taken_rviImm_hi_lo_lo_2 = taken_rviBits_1[20]; // @[Cat.scala 30:58]
  assign taken_rviImm_lo_hi_hi_2 = taken_rviBits_1[30:25]; // @[RocketCore.scala 1043:66]
  assign taken_rviImm_lo_hi_lo_2 = taken_rviBits_1[24:21]; // @[RocketCore.scala 1046:52]
  assign _taken_rviImm_T_7 = {taken_rviImm_hi_hi_hi_2,taken_rviImm_hi_hi_lo_2,taken_rviImm_hi_lo_hi_2,taken_rviImm_hi_lo_lo_2,taken_rviImm_lo_hi_hi_2,taken_rviImm_lo_hi_lo_2,1'h0}; // @[RocketCore.scala 1051:53]
  assign taken_rviImm_hi_lo_hi_3 = {8{taken_rviImm_sign_2}}; // @[Cat.scala 30:58]
  assign taken_rviImm_hi_lo_lo_3 = taken_rviBits_1[7]; // @[Cat.scala 30:58]
  assign _taken_rviImm_T_9 = {taken_rviImm_hi_hi_hi_2,taken_rviImm_hi_hi_lo_2,taken_rviImm_hi_lo_hi_3,taken_rviImm_hi_lo_lo_3,taken_rviImm_lo_hi_hi_2,taken_rviBits_1[11:8],1'h0}; // @[RocketCore.scala 1051:53]
  assign taken_rviImm_1 = taken_rviBits_1[3] ? $signed(_taken_rviImm_T_7) : $signed(_taken_rviImm_T_9); // @[Frontend.scala 227:23]
  assign taken_rvcImm_hi_hi_hi_2 = taken_bits_1[12] ? 5'h1f : 5'h0; // @[Bitwise.scala 72:12]
  assign taken_rvcImm_hi_hi_lo_2 = taken_bits_1[6:5]; // @[RVC.scala 45:35]
  assign taken_rvcImm_hi_lo_2 = taken_bits_1[2]; // @[RVC.scala 45:43]
  assign taken_rvcImm_lo_hi_hi_2 = taken_bits_1[11:10]; // @[RVC.scala 45:49]
  assign taken_rvcImm_lo_hi_lo_2 = taken_bits_1[4:3]; // @[RVC.scala 45:59]
  assign _taken_rvcImm_T_13 = {taken_rvcImm_hi_hi_hi_2,taken_rvcImm_hi_hi_lo_2,taken_rvcImm_hi_lo_2,taken_rvcImm_lo_hi_hi_2,taken_rvcImm_lo_hi_lo_2,1'h0}; // @[Frontend.scala 222:66]
  assign taken_rvcImm_hi_hi_hi_hi_1 = taken_bits_1[12] ? 10'h3ff : 10'h0; // @[Bitwise.scala 72:12]
  assign taken_rvcImm_hi_hi_hi_lo_1 = taken_bits_1[8]; // @[RVC.scala 44:36]
  assign taken_rvcImm_hi_hi_lo_3 = taken_bits_1[10:9]; // @[RVC.scala 44:42]
  assign taken_rvcImm_hi_lo_hi_1 = taken_bits_1[6]; // @[RVC.scala 44:51]
  assign taken_rvcImm_hi_lo_lo_1 = taken_bits_1[7]; // @[RVC.scala 44:57]
  assign taken_rvcImm_lo_hi_lo_3 = taken_bits_1[11]; // @[RVC.scala 44:69]
  assign taken_rvcImm_lo_lo_hi_1 = taken_bits_1[5:3]; // @[RVC.scala 44:76]
  assign _taken_rvcImm_T_17 = {taken_rvcImm_hi_hi_hi_hi_1,taken_rvcImm_hi_hi_hi_lo_1,taken_rvcImm_hi_hi_lo_3,taken_rvcImm_hi_lo_hi_1,taken_rvcImm_hi_lo_lo_1,taken_rvcImm_hi_lo_2,taken_rvcImm_lo_hi_lo_3,taken_rvcImm_lo_lo_hi_1,1'h0}; // @[Frontend.scala 222:106]
  assign taken_rvcImm_1 = taken_bits_1[14] ? $signed({{8{_taken_rvcImm_T_13[12]}},_taken_rvcImm_T_13}) : $signed(_taken_rvcImm_T_17); // @[Frontend.scala 222:23]
  assign _taken_npc_T_9 = taken_prevRVI_1 ? $signed(taken_rviImm_1) : $signed({{11{taken_rvcImm_1[20]}},taken_rvcImm_1}); // @[Frontend.scala 265:69]
  assign _GEN_127 = {{8{_taken_npc_T_9[31]}},_taken_npc_T_9}; // @[Frontend.scala 265:64]
  assign _taken_predicted_npc_T_1 = $signed(_taken_npc_T_8) + $signed(_GEN_127); // @[Frontend.scala 266:34]
  assign _taken_predictBranch_T = taken_prevRVI & taken_rviBranch; // @[Frontend.scala 234:53]
  assign _taken_predictBranch_T_1 = taken_valid & taken_rvcBranch; // @[Frontend.scala 234:75]
  assign _taken_predictBranch_T_2 = _taken_predictBranch_T | _taken_predictBranch_T_1; // @[Frontend.scala 234:66]
  assign taken_predictBranch = s2_btb_resp_bits_bht_value & _taken_predictBranch_T_2; // @[Frontend.scala 234:41]
  assign _taken_predictJump_T = taken_prevRVI & taken_rviJump; // @[Frontend.scala 233:33]
  assign _taken_predictJump_T_1 = taken_valid & taken_rvcJump; // @[Frontend.scala 233:53]
  assign taken_predictJump = _taken_predictJump_T | _taken_predictJump_T_1; // @[Frontend.scala 233:44]
  assign _taken_T_17 = taken_predictBranch | taken_predictJump; // @[Frontend.scala 261:44]
  assign _taken_T_18 = s2_valid & _taken_T_17; // @[Frontend.scala 261:26]
  assign _taken_npc_T = ~_s2_base_pc_T_1; // @[Frontend.scala 264:32]
  assign taken_rviImm_sign = taken_rviBits[31]; // @[RocketCore.scala 1037:53]
  assign taken_rviImm_hi_hi_hi = taken_rviBits[31]; // @[Cat.scala 30:58]
  assign taken_rviImm_hi_hi_lo = {11{taken_rviImm_sign}}; // @[Cat.scala 30:58]
  assign taken_rviImm_hi_lo_hi = taken_rviBits[19:12]; // @[Cat.scala 30:58]
  assign taken_rviImm_hi_lo_lo = taken_rviBits[20]; // @[Cat.scala 30:58]
  assign taken_rviImm_lo_hi_hi = taken_rviBits[30:25]; // @[RocketCore.scala 1043:66]
  assign taken_rviImm_lo_hi_lo = taken_rviBits[24:21]; // @[RocketCore.scala 1046:52]
  assign _taken_rviImm_T_2 = {taken_rviImm_hi_hi_hi,taken_rviImm_hi_hi_lo,taken_rviImm_hi_lo_hi,taken_rviImm_hi_lo_lo,taken_rviImm_lo_hi_hi,taken_rviImm_lo_hi_lo,1'h0}; // @[RocketCore.scala 1051:53]
  assign taken_rviImm_hi_lo_hi_1 = {8{taken_rviImm_sign}}; // @[Cat.scala 30:58]
  assign taken_rviImm_hi_lo_lo_1 = taken_rviBits[7]; // @[Cat.scala 30:58]
  assign _taken_rviImm_T_4 = {taken_rviImm_hi_hi_hi,taken_rviImm_hi_hi_lo,taken_rviImm_hi_lo_hi_1,taken_rviImm_hi_lo_lo_1,taken_rviImm_lo_hi_hi,taken_rviBits[11:8],1'h0}; // @[RocketCore.scala 1051:53]
  assign taken_rviImm = taken_rviBits[3] ? $signed(_taken_rviImm_T_2) : $signed(_taken_rviImm_T_4); // @[Frontend.scala 227:23]
  assign _taken_npc_T_1 = $signed(taken_rviImm) - 32'sh2; // @[Frontend.scala 264:61]
  assign taken_rvcImm_hi_hi_hi = taken_bits[12] ? 5'h1f : 5'h0; // @[Bitwise.scala 72:12]
  assign taken_rvcImm_hi_hi_lo = taken_bits[6:5]; // @[RVC.scala 45:35]
  assign taken_rvcImm_hi_lo = taken_bits[2]; // @[RVC.scala 45:43]
  assign taken_rvcImm_lo_hi_hi = taken_bits[11:10]; // @[RVC.scala 45:49]
  assign taken_rvcImm_lo_hi_lo = taken_bits[4:3]; // @[RVC.scala 45:59]
  assign _taken_rvcImm_T_4 = {taken_rvcImm_hi_hi_hi,taken_rvcImm_hi_hi_lo,taken_rvcImm_hi_lo,taken_rvcImm_lo_hi_hi,taken_rvcImm_lo_hi_lo,1'h0}; // @[Frontend.scala 222:66]
  assign taken_rvcImm_hi_hi_hi_hi = taken_bits[12] ? 10'h3ff : 10'h0; // @[Bitwise.scala 72:12]
  assign taken_rvcImm_hi_hi_hi_lo = taken_bits[8]; // @[RVC.scala 44:36]
  assign taken_rvcImm_hi_hi_lo_1 = taken_bits[10:9]; // @[RVC.scala 44:42]
  assign taken_rvcImm_hi_lo_hi = taken_bits[6]; // @[RVC.scala 44:51]
  assign taken_rvcImm_hi_lo_lo = taken_bits[7]; // @[RVC.scala 44:57]
  assign taken_rvcImm_lo_hi_lo_1 = taken_bits[11]; // @[RVC.scala 44:69]
  assign taken_rvcImm_lo_lo_hi = taken_bits[5:3]; // @[RVC.scala 44:76]
  assign _taken_rvcImm_T_8 = {taken_rvcImm_hi_hi_hi_hi,taken_rvcImm_hi_hi_hi_lo,taken_rvcImm_hi_hi_lo_1,taken_rvcImm_hi_lo_hi,taken_rvcImm_hi_lo_lo,taken_rvcImm_hi_lo,taken_rvcImm_lo_hi_lo_1,taken_rvcImm_lo_lo_hi,1'h0}; // @[Frontend.scala 222:106]
  assign taken_rvcImm = taken_bits[14] ? $signed({{8{_taken_rvcImm_T_4[12]}},_taken_rvcImm_T_4}) : $signed(_taken_rvcImm_T_8); // @[Frontend.scala 222:23]
  assign _taken_npc_T_2 = taken_prevRVI ? $signed(_taken_npc_T_1) : $signed({{12{taken_rvcImm[20]}},taken_rvcImm}); // @[Frontend.scala 264:44]
  assign _GEN_128 = {{7{_taken_npc_T_2[32]}},_taken_npc_T_2}; // @[Frontend.scala 264:39]
  assign _taken_predicted_npc_T = $signed(_taken_npc_T) + $signed(_GEN_128); // @[Frontend.scala 266:34]
  assign predicted_taken = btb_io_resp_valid & btb_io_resp_bits_taken; // @[Frontend.scala 192:29]
  assign predicted_npc_hi = btb_io_resp_bits_target[38]; // @[package.scala 123:38]
  assign _predicted_npc_T = {predicted_npc_hi,btb_io_resp_bits_target}; // @[Cat.scala 30:58]
  assign _GEN_28 = predicted_taken ? _predicted_npc_T : ntpc; // @[Frontend.scala 192:56]
  assign _GEN_43 = _taken_T_18 ? _taken_predicted_npc_T : _GEN_28; // @[Frontend.scala 261:61]
  assign _GEN_46 = s2_btb_taken ? _GEN_28 : _GEN_43; // @[Frontend.scala 254:30]
  assign _GEN_79 = _taken_T_47 ? _taken_predicted_npc_T_1 : _GEN_46; // @[Frontend.scala 261:61]
  assign _GEN_82 = s2_btb_taken ? _GEN_46 : _GEN_79; // @[Frontend.scala 254:30]
  assign _GEN_99 = taken_idx ? _GEN_82 : _GEN_46; // @[Frontend.scala 245:25]
  assign predicted_npc = useRAS ? {{1'd0}, btb_io_ras_head_bits} : _GEN_99; // @[Frontend.scala 305:19]
  assign npc = s2_replay ? s2_pc : predicted_npc; // @[Frontend.scala 128:16]
  assign _s0_speculative_T_1 = s2_valid & ~s2_speculative; // @[Frontend.scala 134:53]
  assign _s0_speculative_T_2 = s1_speculative | _s0_speculative_T_1; // @[Frontend.scala 134:41]
  assign s0_speculative = _s0_speculative_T_2 | predicted_taken; // @[Frontend.scala 134:72]
  assign _taken_taken_T_9 = taken_rviJump_1 | taken_rviJALR_1; // @[Frontend.scala 230:29]
  assign _taken_taken_T_10 = taken_rviBranch_1 & s2_btb_resp_bits_bht_value; // @[Frontend.scala 230:53]
  assign _taken_taken_T_11 = _taken_taken_T_9 | _taken_taken_T_10; // @[Frontend.scala 230:40]
  assign _taken_taken_T_12 = taken_prevRVI_1 & _taken_taken_T_11; // @[Frontend.scala 230:17]
  assign _taken_rvcJALR_T_5 = 16'h9002 == _taken_rvcJR_T_4; // @[Frontend.scala 225:26]
  assign taken_rvcJALR_1 = _taken_rvcJALR_T_5 & _taken_rvcJR_T_7; // @[Frontend.scala 225:49]
  assign _taken_taken_T_13 = taken_rvcJump_1 | taken_rvcJALR_1; // @[Frontend.scala 231:27]
  assign _taken_taken_T_14 = _taken_taken_T_13 | taken_rvcJR_1; // @[Frontend.scala 231:38]
  assign _taken_taken_T_15 = taken_rvcBranch_1 & s2_btb_resp_bits_bht_value; // @[Frontend.scala 231:60]
  assign _taken_taken_T_16 = _taken_taken_T_14 | _taken_taken_T_15; // @[Frontend.scala 231:47]
  assign _taken_taken_T_17 = taken_valid_1 & _taken_taken_T_16; // @[Frontend.scala 231:15]
  assign taken_taken_1 = _taken_taken_T_12 | _taken_taken_T_17; // @[Frontend.scala 230:71]
  assign taken = taken_taken | taken_taken_1; // @[Frontend.scala 286:19]
  assign _GEN_116 = _s2_replay_T | io_cpu_req_valid; // @[Frontend.scala 316:33]
  assign _GEN_120 = taken ? _GEN_116 : io_cpu_req_valid; // @[Frontend.scala 312:20]
  assign s2_redirect = s2_btb_taken ? io_cpu_req_valid : _GEN_120; // @[Frontend.scala 311:26]
  assign _GEN_0 = ~s2_replay & ~s2_redirect; // @[Frontend.scala 140:21]
  assign _icache_io_s1_kill_T = s2_redirect | tlb_io_resp_miss; // @[Frontend.scala 160:36]
  assign s2_can_speculatively_refill = s2_tlb_resp_cacheable & ~io_ptw_customCSRs_csrs_0_value[3]; // @[Frontend.scala 161:59]
  assign _icache_io_s2_kill_T_1 = s2_speculative & ~s2_can_speculatively_refill; // @[Frontend.scala 162:39]
  assign _fq_io_enq_valid_T = fq_io_enq_valid_REG & s2_valid; // @[Frontend.scala 165:40]
  assign _fq_io_enq_valid_T_2 = ~s2_tlb_resp_miss & icache_io_s2_kill; // @[Frontend.scala 165:98]
  assign _fq_io_enq_valid_T_3 = icache_io_resp_valid | _fq_io_enq_valid_T_2; // @[Frontend.scala 165:77]
  assign _io_cpu_npc_T = io_cpu_req_valid ? io_cpu_req_bits_pc : npc; // @[Frontend.scala 167:28]
  assign _io_cpu_npc_T_2 = ~_io_cpu_npc_T | 40'h1; // @[Frontend.scala 341:33]
  assign _fq_io_enq_bits_mask_T_1 = 3'h3 << s2_pc[1]; // @[Frontend.scala 170:52]
  assign _fq_io_enq_bits_replay_T_1 = icache_io_s2_kill & ~icache_io_resp_valid; // @[Frontend.scala 171:76]
  assign _fq_io_enq_bits_replay_T_3 = _fq_io_enq_bits_replay_T_1 & ~s2_xcpt; // @[Frontend.scala 171:101]
  assign _fq_io_enq_bits_replay_T_4 = icache_io_resp_bits_replay | _fq_io_enq_bits_replay_T_3; // @[Frontend.scala 171:55]
  assign _T_13 = s2_speculative & io_ptw_customCSRs_csrs_0_value[3]; // @[Frontend.scala 175:27]
  assign _T_15 = _T_13 & ~icache_io_s2_kill; // @[Frontend.scala 175:110]
  assign _T_18 = ~_T_15 | reset; // @[Frontend.scala 175:9]
  assign _T_20 = icache_io_resp_valid & icache_io_resp_bits_ae; // @[Frontend.scala 176:30]
  assign fetch_bubble_likely = ~fq_io_mask[1]; // @[Frontend.scala 293:33]
  assign _btb_io_btb_update_valid_T_2 = _s2_replay_T & ~wrong_path; // @[Frontend.scala 294:51]
  assign _btb_io_btb_update_valid_T_3 = _btb_io_btb_update_valid_T_2 & fetch_bubble_likely; // @[Frontend.scala 294:66]
  assign _taken_T_53 = taken_predictBranch_1 & s2_btb_resp_bits_bht_value; // @[Frontend.scala 273:52]
  assign _taken_T_54 = _taken_T_53 | taken_predictJump_1; // @[Frontend.scala 273:91]
  assign _taken_T_55 = _taken_T_54 | taken_predictReturn_1; // @[Frontend.scala 273:106]
  assign _taken_T_56 = ~s2_btb_resp_valid & _taken_T_55; // @[Frontend.scala 273:34]
  assign _taken_T_24 = taken_predictBranch & s2_btb_resp_bits_bht_value; // @[Frontend.scala 273:52]
  assign _taken_T_25 = _taken_T_24 | taken_predictJump; // @[Frontend.scala 273:91]
  assign _taken_T_26 = _taken_T_25 | taken_predictReturn; // @[Frontend.scala 273:106]
  assign _taken_T_27 = ~s2_btb_resp_valid & _taken_T_26; // @[Frontend.scala 273:34]
  assign _GEN_92 = _taken_T_56 | _taken_T_27; // @[Frontend.scala 273:125]
  assign updateBTB = taken_idx ? _GEN_92 : _taken_T_27; // @[Frontend.scala 245:25]
  assign _btb_io_btb_update_valid_T_4 = _btb_io_btb_update_valid_T_3 & updateBTB; // @[Frontend.scala 294:89]
  assign _btb_io_btb_update_bits_br_pc_T = {taken_idx, 1'h0}; // @[Frontend.scala 298:63]
  assign _GEN_129 = {{38'd0}, _btb_io_btb_update_bits_br_pc_T}; // @[Frontend.scala 298:50]
  assign _btb_io_btb_update_bits_br_pc_T_1 = s2_base_pc | _GEN_129; // @[Frontend.scala 298:50]
  assign _GEN_36 = io_cpu_btb_update_valid ? {{1'd0}, io_cpu_btb_update_bits_br_pc} : _btb_io_btb_update_bits_br_pc_T_1; // @[Frontend.scala 292:37]
  assign _GEN_37 = io_cpu_btb_update_valid ? {{1'd0}, io_cpu_btb_update_bits_pc} : s2_base_pc; // @[Frontend.scala 292:37]
  assign after_idx = taken_idx ? 2'h2 : 2'h1; // @[Frontend.scala 245:25]
  assign _btb_io_ras_update_bits_returnAddr_T = {after_idx, 1'h0}; // @[Frontend.scala 302:66]
  assign _GEN_130 = {{37'd0}, _btb_io_ras_update_bits_returnAddr_T}; // @[Frontend.scala 302:53]
  assign _btb_io_ras_update_bits_returnAddr_T_2 = s2_base_pc + _GEN_130; // @[Frontend.scala 302:53]
  assign _taken_rviCall_T = taken_rviJALR | taken_rviJump; // @[Frontend.scala 218:30]
  assign taken_rviCall = _taken_rviCall_T & taken_rviBits[7]; // @[Frontend.scala 218:42]
  assign _taken_T = s2_valid & s2_btb_resp_valid; // @[Frontend.scala 236:22]
  assign _taken_T_2 = _taken_T & ~s2_btb_resp_bits_bridx; // @[Frontend.scala 236:43]
  assign _taken_T_3 = _taken_T_2 & taken_valid; // @[Frontend.scala 236:77]
  assign _taken_T_5 = _taken_T_3 & ~_taken_prevRVI_T_4; // @[Frontend.scala 236:86]
  assign _GEN_39 = _taken_T_5 | _fq_io_enq_bits_replay_T_4; // @[Frontend.scala 236:95]
  assign _GEN_40 = _taken_T_5 | wrong_path; // @[Frontend.scala 236:95]
  assign _taken_btb_io_ras_update_valid_T_3 = taken_rviCall | taken_rviReturn; // @[Frontend.scala 248:92]
  assign _taken_btb_io_ras_update_valid_T_4 = taken_prevRVI & _taken_btb_io_ras_update_valid_T_3; // @[Frontend.scala 248:80]
  assign _taken_btb_io_ras_update_valid_T_5 = taken_rvcJALR | taken_rvcReturn; // @[Frontend.scala 248:127]
  assign _taken_btb_io_ras_update_valid_T_6 = taken_valid & _taken_btb_io_ras_update_valid_T_5; // @[Frontend.scala 248:115]
  assign _taken_btb_io_ras_update_valid_T_7 = _taken_btb_io_ras_update_valid_T_4 | _taken_btb_io_ras_update_valid_T_6; // @[Frontend.scala 248:106]
  assign _taken_btb_io_ras_update_valid_T_8 = _btb_io_btb_update_valid_T_2 & _taken_btb_io_ras_update_valid_T_7; // @[Frontend.scala 248:68]
  assign _taken_btb_io_ras_update_bits_cfiType_T = taken_prevRVI ? taken_rviReturn : taken_rvcReturn; // @[Frontend.scala 249:50]
  assign _taken_btb_io_ras_update_bits_cfiType_T_1 = taken_prevRVI ? taken_rviCall : taken_rvcJALR; // @[Frontend.scala 250:50]
  assign _taken_btb_io_ras_update_bits_cfiType_T_2 = taken_prevRVI ? taken_rviBranch : taken_rvcBranch; // @[Frontend.scala 251:50]
  assign _taken_btb_io_ras_update_bits_cfiType_T_5 = _taken_btb_io_ras_update_bits_cfiType_T_2 ? 1'h0 : 1'h1; // @[Frontend.scala 251:46]
  assign _taken_btb_io_ras_update_bits_cfiType_T_6 = _taken_btb_io_ras_update_bits_cfiType_T_1 ? 2'h2 : {{1'd0}, _taken_btb_io_ras_update_bits_cfiType_T_5}; // @[Frontend.scala 250:46]
  assign _taken_btb_io_ras_update_bits_cfiType_T_7 = _taken_btb_io_ras_update_bits_cfiType_T ? 2'h3 : _taken_btb_io_ras_update_bits_cfiType_T_6; // @[Frontend.scala 249:46]
  assign _taken_T_9 = _s2_replay_T & taken_taken; // @[Frontend.scala 255:34]
  assign _taken_T_11 = _taken_T_9 & ~taken_predictBranch; // @[Frontend.scala 255:43]
  assign _taken_T_13 = _taken_T_11 & ~taken_predictJump; // @[Frontend.scala 255:61]
  assign _taken_T_15 = _taken_T_13 & ~taken_predictReturn; // @[Frontend.scala 255:77]
  assign _GEN_41 = _taken_T_15 | _GEN_40; // @[Frontend.scala 255:96]
  assign _GEN_44 = s2_btb_taken ? _GEN_40 : _GEN_41; // @[Frontend.scala 254:30]
  assign _GEN_47 = _taken_predictBranch_T_2 & _btb_io_btb_update_valid_T_2; // @[Frontend.scala 269:59]
  assign taken_rvc_1 = taken_bits_1[1:0] != 2'h3; // @[Frontend.scala 208:45]
  assign _taken_rviCall_T_2 = taken_rviJALR_1 | taken_rviJump_1; // @[Frontend.scala 218:30]
  assign taken_rviCall_1 = _taken_rviCall_T_2 & taken_rviBits_1[7]; // @[Frontend.scala 218:42]
  assign _taken_T_31 = _taken_T & s2_btb_resp_bits_bridx; // @[Frontend.scala 236:43]
  assign _taken_T_32 = _taken_T_31 & taken_valid_1; // @[Frontend.scala 236:77]
  assign _taken_T_34 = _taken_T_32 & ~taken_rvc_1; // @[Frontend.scala 236:86]
  assign _GEN_76 = _taken_T_34 | _GEN_44; // @[Frontend.scala 236:95]
  assign _taken_btb_io_ras_update_valid_T_12 = taken_rviCall_1 | taken_rviReturn_1; // @[Frontend.scala 248:92]
  assign _taken_btb_io_ras_update_valid_T_13 = taken_prevRVI_1 & _taken_btb_io_ras_update_valid_T_12; // @[Frontend.scala 248:80]
  assign _taken_btb_io_ras_update_valid_T_14 = taken_rvcJALR_1 | taken_rvcReturn_1; // @[Frontend.scala 248:127]
  assign _taken_btb_io_ras_update_valid_T_15 = taken_valid_1 & _taken_btb_io_ras_update_valid_T_14; // @[Frontend.scala 248:115]
  assign _taken_btb_io_ras_update_valid_T_16 = _taken_btb_io_ras_update_valid_T_13 | _taken_btb_io_ras_update_valid_T_15; // @[Frontend.scala 248:106]
  assign _taken_btb_io_ras_update_valid_T_17 = _btb_io_btb_update_valid_T_2 & _taken_btb_io_ras_update_valid_T_16; // @[Frontend.scala 248:68]
  assign _taken_btb_io_ras_update_bits_cfiType_T_8 = taken_prevRVI_1 ? taken_rviReturn_1 : taken_rvcReturn_1; // @[Frontend.scala 249:50]
  assign _taken_btb_io_ras_update_bits_cfiType_T_9 = taken_prevRVI_1 ? taken_rviCall_1 : taken_rvcJALR_1; // @[Frontend.scala 250:50]
  assign _taken_btb_io_ras_update_bits_cfiType_T_10 = taken_prevRVI_1 ? taken_rviBranch_1 : taken_rvcBranch_1; // @[Frontend.scala 251:50]
  assign _taken_btb_io_ras_update_bits_cfiType_T_13 = _taken_btb_io_ras_update_bits_cfiType_T_10 ? 1'h0 : 1'h1; // @[Frontend.scala 251:46]
  assign _taken_btb_io_ras_update_bits_cfiType_T_14 = _taken_btb_io_ras_update_bits_cfiType_T_9 ? 2'h2 : {{1'd0}, _taken_btb_io_ras_update_bits_cfiType_T_13}; // @[Frontend.scala 250:46]
  assign _taken_btb_io_ras_update_bits_cfiType_T_15 = _taken_btb_io_ras_update_bits_cfiType_T_8 ? 2'h3 : _taken_btb_io_ras_update_bits_cfiType_T_14; // @[Frontend.scala 249:46]
  assign _taken_T_38 = _s2_replay_T & taken_taken_1; // @[Frontend.scala 255:34]
  assign _taken_T_40 = _taken_T_38 & ~taken_predictBranch_1; // @[Frontend.scala 255:43]
  assign _taken_T_42 = _taken_T_40 & ~taken_predictJump_1; // @[Frontend.scala 255:61]
  assign _taken_T_44 = _taken_T_42 & ~taken_predictReturn_1; // @[Frontend.scala 255:77]
  assign _GEN_77 = _taken_T_44 | _GEN_76; // @[Frontend.scala 255:96]
  assign _GEN_83 = _taken_predictBranch_T_5 ? _btb_io_btb_update_valid_T_2 : _GEN_47; // @[Frontend.scala 269:59]
  assign _taken_T_59 = taken_valid_1 & taken_idx; // @[Frontend.scala 281:23]
  assign _taken_T_61 = _taken_T_59 & ~taken_rvc_1; // @[Frontend.scala 281:37]
  assign _taken_lo_T = taken_bits_1 | 16'h3; // @[Frontend.scala 283:37]
  assign _T_25 = s2_btb_taken | taken; // @[Frontend.scala 308:45]
  assign _T_26 = _s2_replay_T & _T_25; // @[Frontend.scala 308:28]
  assign _GEN_117 = taken ? taken_idx : s2_btb_resp_bits_bridx; // @[Frontend.scala 312:20]
  assign _GEN_118 = taken | s2_btb_taken; // @[Frontend.scala 312:20]
  assign _GEN_119 = taken ? 5'h1c : s2_btb_resp_bits_entry; // @[Frontend.scala 312:20]
  assign _T_31 = ~s2_partial_insn_valid | fq_io_enq_bits_mask[0]; // @[Frontend.scala 320:35]
  assign _T_33 = _T_31 | reset; // @[Frontend.scala 320:11]
  assign auto_icache_master_out_a_valid = icache_auto_master_out_a_valid; // @[LazyModule.scala 311:12]
  assign auto_icache_master_out_a_bits_address = icache_auto_master_out_a_bits_address; // @[LazyModule.scala 311:12]
  assign io_cpu_resp_valid = fq_io_deq_valid; // @[Frontend.scala 325:15]
  assign io_cpu_resp_bits_btb_taken = fq_io_deq_bits_btb_taken; // @[Frontend.scala 325:15]
  assign io_cpu_resp_bits_btb_bridx = fq_io_deq_bits_btb_bridx; // @[Frontend.scala 325:15]
  assign io_cpu_resp_bits_btb_entry = fq_io_deq_bits_btb_entry; // @[Frontend.scala 325:15]
  assign io_cpu_resp_bits_btb_bht_history = fq_io_deq_bits_btb_bht_history; // @[Frontend.scala 325:15]
  assign io_cpu_resp_bits_pc = fq_io_deq_bits_pc; // @[Frontend.scala 325:15]
  assign io_cpu_resp_bits_data = fq_io_deq_bits_data; // @[Frontend.scala 325:15]
  assign io_cpu_resp_bits_xcpt_pf_inst = fq_io_deq_bits_xcpt_pf_inst; // @[Frontend.scala 325:15]
  assign io_cpu_resp_bits_xcpt_ae_inst = fq_io_deq_bits_xcpt_ae_inst; // @[Frontend.scala 325:15]
  assign io_cpu_resp_bits_replay = fq_io_deq_bits_replay; // @[Frontend.scala 325:15]
  assign io_cpu_npc = ~_io_cpu_npc_T_2; // @[Frontend.scala 167:14]
  assign io_ptw_req_valid = tlb_io_ptw_req_valid; // @[Frontend.scala 147:10]
  assign io_ptw_req_bits_valid = tlb_io_ptw_req_bits_valid; // @[Frontend.scala 147:10]
  assign io_ptw_req_bits_bits_addr = tlb_io_ptw_req_bits_bits_addr; // @[Frontend.scala 147:10]
  assign icache_clock = gated_clock; // @[Frontend.scala 94:16]
  assign icache_reset = reset;
  assign icache_auto_master_out_a_ready = auto_icache_master_out_a_ready; // @[LazyModule.scala 311:12]
  assign icache_auto_master_out_d_valid = auto_icache_master_out_d_valid; // @[LazyModule.scala 311:12]
  assign icache_auto_master_out_d_bits_opcode = auto_icache_master_out_d_bits_opcode; // @[LazyModule.scala 311:12]
  assign icache_auto_master_out_d_bits_size = auto_icache_master_out_d_bits_size; // @[LazyModule.scala 311:12]
  assign icache_auto_master_out_d_bits_data = auto_icache_master_out_d_bits_data; // @[LazyModule.scala 311:12]
  assign icache_auto_master_out_d_bits_corrupt = auto_icache_master_out_d_bits_corrupt; // @[LazyModule.scala 311:12]
  assign icache_io_req_valid = io_cpu_req_valid | s0_fq_has_space; // @[Frontend.scala 155:23]
  assign icache_io_req_bits_addr = io_cpu_npc[38:0]; // @[Frontend.scala 156:27]
  assign icache_io_s1_paddr = tlb_io_resp_paddr; // @[Frontend.scala 158:22]
  assign icache_io_s1_kill = _icache_io_s1_kill_T | s2_replay; // @[Frontend.scala 160:21]
  assign icache_io_s2_kill = _icache_io_s2_kill_T_1 | s2_xcpt; // @[Frontend.scala 162:21]
  assign icache_io_invalidate = io_cpu_flush_icache; // @[Frontend.scala 157:24]
  assign fq_clock = gated_clock;
  assign fq_reset = reset | io_cpu_req_valid;
  assign fq_io_enq_valid = _fq_io_enq_valid_T & _fq_io_enq_valid_T_3; // @[Frontend.scala 165:19]
  assign fq_io_enq_bits_btb_taken = s2_btb_taken ? s2_btb_taken : _GEN_118; // @[Frontend.scala 172:22 Frontend.scala 173:28 Frontend.scala 314:34]
  assign fq_io_enq_bits_btb_bridx = s2_btb_taken ? s2_btb_resp_bits_bridx : _GEN_117; // @[Frontend.scala 172:22 Frontend.scala 313:34]
  assign fq_io_enq_bits_btb_entry = s2_btb_taken ? s2_btb_resp_bits_entry : _GEN_119; // @[Frontend.scala 172:22 Frontend.scala 315:34]
  assign fq_io_enq_bits_btb_bht_history = s2_btb_resp_bits_bht_history; // @[Frontend.scala 172:22]
  assign fq_io_enq_bits_pc = s2_pc; // @[Frontend.scala 166:21]
  assign fq_io_enq_bits_data = icache_io_resp_bits_data; // @[Frontend.scala 169:23]
  assign fq_io_enq_bits_mask = _fq_io_enq_bits_mask_T_1[1:0]; // @[Frontend.scala 170:23]
  assign fq_io_enq_bits_xcpt_pf_inst = s2_tlb_resp_pf_inst; // @[Frontend.scala 174:23]
  assign fq_io_enq_bits_xcpt_ae_inst = _T_20 | s2_tlb_resp_ae_inst; // @[Frontend.scala 174:23 Frontend.scala 176:87]
  assign fq_io_enq_bits_replay = _taken_T_34 | _GEN_39; // @[Frontend.scala 171:25 Frontend.scala 240:31 Frontend.scala 240:31]
  assign fq_io_deq_ready = io_cpu_resp_ready; // @[Frontend.scala 325:15]
  assign tlb_clock = gated_clock;
  assign tlb_reset = reset;
  assign tlb_io_req_valid = s1_valid & ~s2_replay; // @[Frontend.scala 148:20]
  assign tlb_io_req_bits_vaddr = s1_pc; // @[Frontend.scala 149:25]
  assign tlb_io_sfence_valid = io_cpu_sfence_valid; // @[Frontend.scala 152:17]
  assign tlb_io_sfence_bits_rs1 = io_cpu_sfence_bits_rs1; // @[Frontend.scala 152:17]
  assign tlb_io_sfence_bits_rs2 = io_cpu_sfence_bits_rs2; // @[Frontend.scala 152:17]
  assign tlb_io_sfence_bits_addr = io_cpu_sfence_bits_addr; // @[Frontend.scala 152:17]
  assign tlb_io_ptw_req_ready = io_ptw_req_ready; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_resp_valid = io_ptw_resp_valid; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_resp_bits_ae = io_ptw_resp_bits_ae; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_resp_bits_pte_ppn = io_ptw_resp_bits_pte_ppn; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_resp_bits_pte_d = io_ptw_resp_bits_pte_d; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_resp_bits_pte_a = io_ptw_resp_bits_pte_a; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_resp_bits_pte_g = io_ptw_resp_bits_pte_g; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_resp_bits_pte_u = io_ptw_resp_bits_pte_u; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_resp_bits_pte_x = io_ptw_resp_bits_pte_x; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_resp_bits_pte_w = io_ptw_resp_bits_pte_w; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_resp_bits_pte_r = io_ptw_resp_bits_pte_r; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_resp_bits_pte_v = io_ptw_resp_bits_pte_v; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_resp_bits_level = io_ptw_resp_bits_level; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_resp_bits_homogeneous = io_ptw_resp_bits_homogeneous; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_ptbr_mode = io_ptw_ptbr_mode; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_status_debug = io_ptw_status_debug; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_status_prv = io_ptw_status_prv; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_0_cfg_l = io_ptw_pmp_0_cfg_l; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_0_cfg_a = io_ptw_pmp_0_cfg_a; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_0_cfg_x = io_ptw_pmp_0_cfg_x; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_0_cfg_w = io_ptw_pmp_0_cfg_w; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_0_cfg_r = io_ptw_pmp_0_cfg_r; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_0_addr = io_ptw_pmp_0_addr; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_0_mask = io_ptw_pmp_0_mask; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_1_cfg_l = io_ptw_pmp_1_cfg_l; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_1_cfg_a = io_ptw_pmp_1_cfg_a; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_1_cfg_x = io_ptw_pmp_1_cfg_x; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_1_cfg_w = io_ptw_pmp_1_cfg_w; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_1_cfg_r = io_ptw_pmp_1_cfg_r; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_1_addr = io_ptw_pmp_1_addr; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_1_mask = io_ptw_pmp_1_mask; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_2_cfg_l = io_ptw_pmp_2_cfg_l; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_2_cfg_a = io_ptw_pmp_2_cfg_a; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_2_cfg_x = io_ptw_pmp_2_cfg_x; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_2_cfg_w = io_ptw_pmp_2_cfg_w; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_2_cfg_r = io_ptw_pmp_2_cfg_r; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_2_addr = io_ptw_pmp_2_addr; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_2_mask = io_ptw_pmp_2_mask; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_3_cfg_l = io_ptw_pmp_3_cfg_l; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_3_cfg_a = io_ptw_pmp_3_cfg_a; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_3_cfg_x = io_ptw_pmp_3_cfg_x; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_3_cfg_w = io_ptw_pmp_3_cfg_w; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_3_cfg_r = io_ptw_pmp_3_cfg_r; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_3_addr = io_ptw_pmp_3_addr; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_3_mask = io_ptw_pmp_3_mask; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_4_cfg_l = io_ptw_pmp_4_cfg_l; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_4_cfg_a = io_ptw_pmp_4_cfg_a; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_4_cfg_x = io_ptw_pmp_4_cfg_x; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_4_cfg_w = io_ptw_pmp_4_cfg_w; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_4_cfg_r = io_ptw_pmp_4_cfg_r; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_4_addr = io_ptw_pmp_4_addr; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_4_mask = io_ptw_pmp_4_mask; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_5_cfg_l = io_ptw_pmp_5_cfg_l; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_5_cfg_a = io_ptw_pmp_5_cfg_a; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_5_cfg_x = io_ptw_pmp_5_cfg_x; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_5_cfg_w = io_ptw_pmp_5_cfg_w; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_5_cfg_r = io_ptw_pmp_5_cfg_r; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_5_addr = io_ptw_pmp_5_addr; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_5_mask = io_ptw_pmp_5_mask; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_6_cfg_l = io_ptw_pmp_6_cfg_l; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_6_cfg_a = io_ptw_pmp_6_cfg_a; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_6_cfg_x = io_ptw_pmp_6_cfg_x; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_6_cfg_w = io_ptw_pmp_6_cfg_w; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_6_cfg_r = io_ptw_pmp_6_cfg_r; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_6_addr = io_ptw_pmp_6_addr; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_6_mask = io_ptw_pmp_6_mask; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_7_cfg_l = io_ptw_pmp_7_cfg_l; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_7_cfg_a = io_ptw_pmp_7_cfg_a; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_7_cfg_x = io_ptw_pmp_7_cfg_x; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_7_cfg_w = io_ptw_pmp_7_cfg_w; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_7_cfg_r = io_ptw_pmp_7_cfg_r; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_7_addr = io_ptw_pmp_7_addr; // @[Frontend.scala 147:10]
  assign tlb_io_ptw_pmp_7_mask = io_ptw_pmp_7_mask; // @[Frontend.scala 147:10]
  assign tlb_io_kill = ~s2_valid; // @[Frontend.scala 153:15]
  assign btb_clock = gated_clock;
  assign btb_reset = reset;
  assign btb_io_req_bits_addr = s1_pc[38:0]; // @[Frontend.scala 182:26]
  assign btb_io_btb_update_valid = io_cpu_btb_update_valid ? io_cpu_btb_update_valid : _btb_io_btb_update_valid_T_4; // @[Frontend.scala 183:23 Frontend.scala 294:31]
  assign btb_io_btb_update_bits_prediction_entry = io_cpu_btb_update_valid ? io_cpu_btb_update_bits_prediction_entry : 5'h1c; // @[Frontend.scala 183:23 Frontend.scala 295:47]
  assign btb_io_btb_update_bits_pc = _GEN_37[38:0]; // @[Frontend.scala 183:23 Frontend.scala 299:33]
  assign btb_io_btb_update_bits_isValid = ~io_cpu_btb_update_valid | io_cpu_btb_update_bits_isValid; // @[Frontend.scala 183:23 Frontend.scala 296:38]
  assign btb_io_btb_update_bits_br_pc = _GEN_36[38:0]; // @[Frontend.scala 183:23 Frontend.scala 298:36]
  assign btb_io_btb_update_bits_cfiType = io_cpu_btb_update_valid ? io_cpu_btb_update_bits_cfiType : btb_io_ras_update_bits_cfiType; // @[Frontend.scala 183:23 Frontend.scala 297:38]
  assign btb_io_bht_update_valid = io_cpu_bht_update_valid; // @[Frontend.scala 184:23 Frontend.scala 199:50]
  assign btb_io_bht_update_bits_prediction_history = io_cpu_bht_update_bits_prediction_history; // @[Frontend.scala 184:23]
  assign btb_io_bht_update_bits_pc = io_cpu_bht_update_bits_pc; // @[Frontend.scala 184:23]
  assign btb_io_bht_update_bits_branch = io_cpu_bht_update_bits_branch; // @[Frontend.scala 184:23]
  assign btb_io_bht_update_bits_taken = io_cpu_bht_update_bits_taken; // @[Frontend.scala 184:23]
  assign btb_io_bht_update_bits_mispredict = io_cpu_bht_update_bits_mispredict; // @[Frontend.scala 184:23]
  assign btb_io_bht_advance_valid = taken_idx ? _GEN_83 : _GEN_47; // @[Frontend.scala 186:30 Frontend.scala 270:36 Frontend.scala 270:36]
  assign btb_io_bht_advance_bits_bht_value = s2_btb_resp_bits_bht_value; // @[Frontend.scala 271:35 Frontend.scala 271:35]
  assign btb_io_ras_update_valid = taken_idx ? _taken_btb_io_ras_update_valid_T_17 : _taken_btb_io_ras_update_valid_T_8; // @[Frontend.scala 185:29 Frontend.scala 248:33 Frontend.scala 248:33]
  assign btb_io_ras_update_bits_cfiType = taken_idx ? _taken_btb_io_ras_update_bits_cfiType_T_15 : _taken_btb_io_ras_update_bits_cfiType_T_7; // @[Frontend.scala 249:40 Frontend.scala 249:40]
  assign btb_io_ras_update_bits_returnAddr = _btb_io_ras_update_bits_returnAddr_T_2[38:0]; // @[Frontend.scala 302:39]
  assign btb_io_flush = _taken_T_34 | _taken_T_5; // @[Frontend.scala 180:18 Frontend.scala 198:54 Frontend.scala 239:22 Frontend.scala 239:22]
  assign Frontend_cov_read_addr = Frontend_state;
  assign Frontend_cov_read_data = Frontend_cov[Frontend_cov_read_addr]; // @[Coverage map for Frontend]
  assign Frontend_cov_write_data = 1'h1;
  assign Frontend_cov_write_addr = Frontend_state;
  assign Frontend_cov_write_mask = 1'h1;
  assign Frontend_cov_write_en = 1'h1;
  assign s2_partial_insn_valid_shl = s2_partial_insn_valid;
  assign s2_partial_insn_valid_pad = {5'h0,s2_partial_insn_valid_shl};
  assign s2_btb_resp_valid_shl = {s2_btb_resp_valid, 1'h0};
  assign s2_btb_resp_valid_pad = {4'h0,s2_btb_resp_valid_shl};
  assign s2_replay_REG_shl = {s2_replay_REG, 2'h0};
  assign s2_replay_REG_pad = {3'h0,s2_replay_REG_shl};
  assign s2_btb_resp_bits_bht_value_shl = {s2_btb_resp_bits_bht_value, 3'h0};
  assign s2_btb_resp_bits_bht_value_pad = {2'h0,s2_btb_resp_bits_bht_value_shl};
  assign s2_valid_shl = {s2_valid, 4'h0};
  assign s2_valid_pad = {1'h0,s2_valid_shl};
  assign s2_btb_resp_bits_taken_shl = {s2_btb_resp_bits_taken, 5'h0};
  assign s2_btb_resp_bits_taken_pad = s2_btb_resp_bits_taken_shl;
  assign Frontend_xor4 = s2_btb_resp_valid_pad ^ s2_replay_REG_pad;
  assign Frontend_xor1 = s2_partial_insn_valid_pad ^ Frontend_xor4;
  assign Frontend_xor6 = s2_valid_pad ^ s2_btb_resp_bits_taken_pad;
  assign Frontend_xor2 = s2_btb_resp_bits_bht_value_pad ^ Frontend_xor6;
  assign Frontend_xor0 = Frontend_xor1 ^ Frontend_xor2;
  assign icache_sum = Frontend_covSum + icache_io_covSum;
  assign fq_sum = icache_sum + fq_io_covSum;
  assign tlb_sum = fq_sum + tlb_io_covSum;
  assign btb_sum = tlb_sum + btb_io_covSum;
  assign io_covSum = btb_sum;
  assign stopEn0 = ~_T_9;
  assign stopEn1 = ~_T_18;
  assign stopEn2 = ~_T_33;
  assign icache_metaAssert_wire = icache_metaAssert;
  assign fq_metaAssert_wire = fq_metaAssert;
  assign tlb_metaAssert_wire = tlb_metaAssert;
  assign btb_metaAssert_wire = btb_metaAssert;
  assign Frontend_or4 = stopEn1 | stopEn2;
  assign Frontend_or1 = stopEn0 | Frontend_or4;
  assign Frontend_or5 = icache_metaAssert_wire | fq_metaAssert_wire;
  assign Frontend_or6 = tlb_metaAssert_wire | btb_metaAssert_wire;
  assign Frontend_or2 = Frontend_or5 | Frontend_or6;
  assign Frontend_or0 = Frontend_or1 | Frontend_or2;
  assign metaAssert = Frontend_or0;
  assign icache_metaReset = metaReset | icache_halt;
  assign fq_metaReset = metaReset | fq_halt;
  assign tlb_metaReset = metaReset | tlb_halt;
  assign btb_metaReset = metaReset | btb_halt;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s1_valid = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  s2_valid = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {2{`RANDOM}};
  s1_pc = _RAND_2[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  s1_speculative = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {2{`RANDOM}};
  s2_pc = _RAND_4[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  s2_btb_resp_valid = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  s2_btb_resp_bits_taken = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  s2_btb_resp_bits_bridx = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  s2_btb_resp_bits_entry = _RAND_8[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  s2_btb_resp_bits_bht_history = _RAND_9[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  s2_btb_resp_bits_bht_value = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  s2_tlb_resp_miss = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  s2_tlb_resp_pf_inst = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  s2_tlb_resp_ae_inst = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  s2_tlb_resp_cacheable = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  s2_speculative = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  s2_partial_insn_valid = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  s2_partial_insn = _RAND_17[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  wrong_path = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  s2_replay_REG = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  fq_io_enq_valid_REG = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  Frontend_state = _RAND_21[5:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    Frontend_cov[initvar] = _RAND_22[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  Frontend_covSum = _RAND_23[29:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge gated_clock) begin
    if (metaReset) begin
      s1_valid <= 1'h0;
    end else begin
      s1_valid <= io_cpu_req_valid | s0_fq_has_space;
    end
    if (metaReset) begin
      s2_valid <= 1'h0;
    end else if (reset) begin
      s2_valid <= 1'h0;
    end else begin
      s2_valid <= _GEN_0;
    end
    if (metaReset) begin
      s1_pc <= 40'h0;
    end else begin
      s1_pc <= io_cpu_npc;
    end
    if (metaReset) begin
      s1_speculative <= 1'h0;
    end else if (io_cpu_req_valid) begin
      s1_speculative <= io_cpu_req_bits_speculative;
    end else if (s2_replay) begin
      s1_speculative <= s2_speculative;
    end else begin
      s1_speculative <= s0_speculative;
    end
    if (metaReset) begin
      s2_pc <= 40'h0;
    end else if (reset) begin
      s2_pc <= {{8'd0}, ~_s2_pc_T_1};
    end else if (~s2_replay) begin
      s2_pc <= s1_pc;
    end
    if (metaReset) begin
      s2_btb_resp_valid <= 1'h0;
    end else if (~s2_replay) begin
      s2_btb_resp_valid <= btb_io_resp_valid;
    end
    if (metaReset) begin
      s2_btb_resp_bits_taken <= 1'h0;
    end else if (~s2_replay) begin
      s2_btb_resp_bits_taken <= btb_io_resp_bits_taken;
    end
    if (metaReset) begin
      s2_btb_resp_bits_bridx <= 1'h0;
    end else if (~s2_replay) begin
      s2_btb_resp_bits_bridx <= btb_io_resp_bits_bridx;
    end
    if (metaReset) begin
      s2_btb_resp_bits_entry <= 5'h0;
    end else if (~s2_replay) begin
      s2_btb_resp_bits_entry <= btb_io_resp_bits_entry;
    end
    if (metaReset) begin
      s2_btb_resp_bits_bht_history <= 8'h0;
    end else if (~s2_replay) begin
      s2_btb_resp_bits_bht_history <= btb_io_resp_bits_bht_history;
    end
    if (metaReset) begin
      s2_btb_resp_bits_bht_value <= 1'h0;
    end else if (~s2_replay) begin
      s2_btb_resp_bits_bht_value <= btb_io_resp_bits_bht_value;
    end
    if (metaReset) begin
      s2_tlb_resp_miss <= 1'h0;
    end else if (~s2_replay) begin
      s2_tlb_resp_miss <= tlb_io_resp_miss;
    end
    if (metaReset) begin
      s2_tlb_resp_pf_inst <= 1'h0;
    end else if (~s2_replay) begin
      s2_tlb_resp_pf_inst <= tlb_io_resp_pf_inst;
    end
    if (metaReset) begin
      s2_tlb_resp_ae_inst <= 1'h0;
    end else if (~s2_replay) begin
      s2_tlb_resp_ae_inst <= tlb_io_resp_ae_inst;
    end
    if (metaReset) begin
      s2_tlb_resp_cacheable <= 1'h0;
    end else if (~s2_replay) begin
      s2_tlb_resp_cacheable <= tlb_io_resp_cacheable;
    end
    if (metaReset) begin
      s2_speculative <= 1'h0;
    end else if (reset) begin
      s2_speculative <= 1'h0;
    end else if (~s2_replay) begin
      s2_speculative <= s1_speculative;
    end
    if (metaReset) begin
      s2_partial_insn_valid <= 1'h0;
    end else if (reset) begin
      s2_partial_insn_valid <= 1'h0;
    end else if (s2_redirect) begin
      s2_partial_insn_valid <= 1'h0;
    end else if (_T_26) begin
      s2_partial_insn_valid <= 1'h0;
    end else if (_s2_replay_T) begin
      s2_partial_insn_valid <= _taken_T_61;
    end
    if (metaReset) begin
      s2_partial_insn <= 16'h0;
    end else if (_s2_replay_T) begin
      if (_taken_T_61) begin
        s2_partial_insn <= _taken_lo_T;
      end
    end
    if (metaReset) begin
      wrong_path <= 1'h0;
    end else if (reset) begin
      wrong_path <= 1'h0;
    end else if (io_cpu_req_valid) begin
      wrong_path <= 1'h0;
    end else if (taken_idx) begin
      if (~s2_btb_taken) begin
        wrong_path <= _GEN_77;
      end else begin
        wrong_path <= _GEN_76;
      end
    end else begin
      wrong_path <= _GEN_76;
    end
    if (metaReset) begin
      s2_replay_REG <= 1'h0;
    end else begin
      s2_replay_REG <= reset | _s2_replay_T_4;
    end
    if (metaReset) begin
      fq_io_enq_valid_REG <= 1'h0;
    end else begin
      fq_io_enq_valid_REG <= s1_valid;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_9) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Frontend.scala:89 assert(!(io.cpu.req.valid || io.cpu.sfence.valid || io.cpu.flush_icache || io.cpu.bht_update.valid || io.cpu.btb_update.valid) || io.cpu.might_request)\n"); // @[Frontend.scala 89:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_9) begin
          $fatal; // @[Frontend.scala 89:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_18) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Frontend.scala:175 assert(!(s2_speculative && io.ptw.customCSRs.asInstanceOf[RocketCustomCSRs].disableSpeculativeICacheRefill && !icache.io.s2_kill))\n"); // @[Frontend.scala 175:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_18) begin
          $fatal; // @[Frontend.scala 175:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_33) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Frontend.scala:320 assert(!s2_partial_insn_valid || fq.io.enq.bits.mask(0))\n"); // @[Frontend.scala 320:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_33) begin
          $fatal; // @[Frontend.scala 320:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    Frontend_state <= Frontend_xor0;
    if (!(Frontend_cov_read_data)) begin
      Frontend_covSum <= Frontend_covSum + 1'h1;
    end
  end
  always @(posedge gated_clock) begin
    if(Frontend_cov_write_en & Frontend_cov_write_mask) begin
      Frontend_cov[Frontend_cov_write_addr] <= Frontend_cov_write_data; // @[Coverage map for Frontend]
    end
  end
endmodule
module FPU(
  input         clock,
  input         reset,
  input  [31:0] io_inst,
  input  [63:0] io_fromint_data,
  input  [2:0]  io_fcsr_rm,
  output        io_fcsr_flags_valid,
  output [4:0]  io_fcsr_flags_bits,
  output [63:0] io_store_data,
  output [63:0] io_toint_data,
  input         io_dmem_resp_val,
  input  [2:0]  io_dmem_resp_type,
  input  [4:0]  io_dmem_resp_tag,
  input  [63:0] io_dmem_resp_data,
  input         io_valid,
  output        io_fcsr_rdy,
  output        io_nack_mem,
  output        io_illegal_rm,
  input         io_killx,
  input         io_killm,
  output        io_dec_wen,
  output        io_dec_ren1,
  output        io_dec_ren2,
  output        io_dec_ren3,
  output        io_sboard_set,
  output        io_sboard_clr,
  output [4:0]  io_sboard_clra,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset,
  input         fpiu_halt,
  input         ifpu_halt,
  input         sfma_halt,
  input         fpmu_halt,
  input         divSqrt_1_halt,
  input         dfma_halt,
  input         divSqrt_halt
);
  wire [31:0] fp_decoder_io_inst; // @[FPU.scala 742:26]
  wire  fp_decoder_io_sigs_wen; // @[FPU.scala 742:26]
  wire  fp_decoder_io_sigs_ren1; // @[FPU.scala 742:26]
  wire  fp_decoder_io_sigs_ren2; // @[FPU.scala 742:26]
  wire  fp_decoder_io_sigs_ren3; // @[FPU.scala 742:26]
  wire  fp_decoder_io_sigs_swap12; // @[FPU.scala 742:26]
  wire  fp_decoder_io_sigs_swap23; // @[FPU.scala 742:26]
  wire [1:0] fp_decoder_io_sigs_typeTagIn; // @[FPU.scala 742:26]
  wire [1:0] fp_decoder_io_sigs_typeTagOut; // @[FPU.scala 742:26]
  wire  fp_decoder_io_sigs_fromint; // @[FPU.scala 742:26]
  wire  fp_decoder_io_sigs_toint; // @[FPU.scala 742:26]
  wire  fp_decoder_io_sigs_fastpipe; // @[FPU.scala 742:26]
  wire  fp_decoder_io_sigs_fma; // @[FPU.scala 742:26]
  wire  fp_decoder_io_sigs_div; // @[FPU.scala 742:26]
  wire  fp_decoder_io_sigs_sqrt; // @[FPU.scala 742:26]
  wire  fp_decoder_io_sigs_wflags; // @[FPU.scala 742:26]
  wire [29:0] fp_decoder_io_covSum; // @[FPU.scala 742:26]
  wire  fp_decoder_metaAssert; // @[FPU.scala 742:26]
  reg [64:0] regfile [0:31]; // @[FPU.scala 796:20]
  reg [95:0] _RAND_0;
  wire [64:0] regfile_ex_rs_0_data; // @[FPU.scala 796:20]
  wire [4:0] regfile_ex_rs_0_addr; // @[FPU.scala 796:20]
  wire [64:0] regfile_ex_rs_1_data; // @[FPU.scala 796:20]
  wire [4:0] regfile_ex_rs_1_addr; // @[FPU.scala 796:20]
  wire [64:0] regfile_ex_rs_2_data; // @[FPU.scala 796:20]
  wire [4:0] regfile_ex_rs_2_addr; // @[FPU.scala 796:20]
  wire [64:0] regfile_MPORT_data; // @[FPU.scala 796:20]
  wire [4:0] regfile_MPORT_addr; // @[FPU.scala 796:20]
  wire  regfile_MPORT_mask; // @[FPU.scala 796:20]
  wire  regfile_MPORT_en; // @[FPU.scala 796:20]
  wire [64:0] regfile_MPORT_1_data; // @[FPU.scala 796:20]
  wire [4:0] regfile_MPORT_1_addr; // @[FPU.scala 796:20]
  wire  regfile_MPORT_1_mask; // @[FPU.scala 796:20]
  wire  regfile_MPORT_1_en; // @[FPU.scala 796:20]
  wire  sfma_clock; // @[FPU.scala 844:20]
  wire  sfma_reset; // @[FPU.scala 844:20]
  wire  sfma_io_in_valid; // @[FPU.scala 844:20]
  wire  sfma_io_in_bits_ren3; // @[FPU.scala 844:20]
  wire  sfma_io_in_bits_swap23; // @[FPU.scala 844:20]
  wire [2:0] sfma_io_in_bits_rm; // @[FPU.scala 844:20]
  wire [1:0] sfma_io_in_bits_fmaCmd; // @[FPU.scala 844:20]
  wire [64:0] sfma_io_in_bits_in1; // @[FPU.scala 844:20]
  wire [64:0] sfma_io_in_bits_in2; // @[FPU.scala 844:20]
  wire [64:0] sfma_io_in_bits_in3; // @[FPU.scala 844:20]
  wire [64:0] sfma_io_out_bits_data; // @[FPU.scala 844:20]
  wire [4:0] sfma_io_out_bits_exc; // @[FPU.scala 844:20]
  wire [29:0] sfma_io_covSum; // @[FPU.scala 844:20]
  wire  sfma_metaAssert; // @[FPU.scala 844:20]
  wire  sfma_metaReset; // @[FPU.scala 844:20]
  wire  sfma_fma_halt; // @[FPU.scala 844:20]
  wire  fpiu_clock; // @[FPU.scala 848:20]
  wire  fpiu_io_in_valid; // @[FPU.scala 848:20]
  wire  fpiu_io_in_bits_ren2; // @[FPU.scala 848:20]
  wire [1:0] fpiu_io_in_bits_typeTagIn; // @[FPU.scala 848:20]
  wire [1:0] fpiu_io_in_bits_typeTagOut; // @[FPU.scala 848:20]
  wire  fpiu_io_in_bits_wflags; // @[FPU.scala 848:20]
  wire [2:0] fpiu_io_in_bits_rm; // @[FPU.scala 848:20]
  wire [1:0] fpiu_io_in_bits_typ; // @[FPU.scala 848:20]
  wire [1:0] fpiu_io_in_bits_fmt; // @[FPU.scala 848:20]
  wire [64:0] fpiu_io_in_bits_in1; // @[FPU.scala 848:20]
  wire [64:0] fpiu_io_in_bits_in2; // @[FPU.scala 848:20]
  wire [2:0] fpiu_io_out_bits_in_rm; // @[FPU.scala 848:20]
  wire [64:0] fpiu_io_out_bits_in_in1; // @[FPU.scala 848:20]
  wire [64:0] fpiu_io_out_bits_in_in2; // @[FPU.scala 848:20]
  wire  fpiu_io_out_bits_lt; // @[FPU.scala 848:20]
  wire [63:0] fpiu_io_out_bits_store; // @[FPU.scala 848:20]
  wire [63:0] fpiu_io_out_bits_toint; // @[FPU.scala 848:20]
  wire [4:0] fpiu_io_out_bits_exc; // @[FPU.scala 848:20]
  wire [29:0] fpiu_io_covSum; // @[FPU.scala 848:20]
  wire  fpiu_metaAssert; // @[FPU.scala 848:20]
  wire  fpiu_metaReset; // @[FPU.scala 848:20]
  wire  ifpu_clock; // @[FPU.scala 858:20]
  wire  ifpu_reset; // @[FPU.scala 858:20]
  wire  ifpu_io_in_valid; // @[FPU.scala 858:20]
  wire [1:0] ifpu_io_in_bits_typeTagIn; // @[FPU.scala 858:20]
  wire  ifpu_io_in_bits_wflags; // @[FPU.scala 858:20]
  wire [2:0] ifpu_io_in_bits_rm; // @[FPU.scala 858:20]
  wire [1:0] ifpu_io_in_bits_typ; // @[FPU.scala 858:20]
  wire [63:0] ifpu_io_in_bits_in1; // @[FPU.scala 858:20]
  wire [64:0] ifpu_io_out_bits_data; // @[FPU.scala 858:20]
  wire [4:0] ifpu_io_out_bits_exc; // @[FPU.scala 858:20]
  wire [29:0] ifpu_io_covSum; // @[FPU.scala 858:20]
  wire  ifpu_metaAssert; // @[FPU.scala 858:20]
  wire  ifpu_metaReset; // @[FPU.scala 858:20]
  wire  fpmu_clock; // @[FPU.scala 863:20]
  wire  fpmu_reset; // @[FPU.scala 863:20]
  wire  fpmu_io_in_valid; // @[FPU.scala 863:20]
  wire  fpmu_io_in_bits_ren2; // @[FPU.scala 863:20]
  wire [1:0] fpmu_io_in_bits_typeTagOut; // @[FPU.scala 863:20]
  wire  fpmu_io_in_bits_wflags; // @[FPU.scala 863:20]
  wire [2:0] fpmu_io_in_bits_rm; // @[FPU.scala 863:20]
  wire [64:0] fpmu_io_in_bits_in1; // @[FPU.scala 863:20]
  wire [64:0] fpmu_io_in_bits_in2; // @[FPU.scala 863:20]
  wire [64:0] fpmu_io_out_bits_data; // @[FPU.scala 863:20]
  wire [4:0] fpmu_io_out_bits_exc; // @[FPU.scala 863:20]
  wire  fpmu_io_lt; // @[FPU.scala 863:20]
  wire [29:0] fpmu_io_covSum; // @[FPU.scala 863:20]
  wire  fpmu_metaAssert; // @[FPU.scala 863:20]
  wire  fpmu_metaReset; // @[FPU.scala 863:20]
  wire  dfma_clock; // @[FPU.scala 882:28]
  wire  dfma_reset; // @[FPU.scala 882:28]
  wire  dfma_io_in_valid; // @[FPU.scala 882:28]
  wire  dfma_io_in_bits_ren3; // @[FPU.scala 882:28]
  wire  dfma_io_in_bits_swap23; // @[FPU.scala 882:28]
  wire [2:0] dfma_io_in_bits_rm; // @[FPU.scala 882:28]
  wire [1:0] dfma_io_in_bits_fmaCmd; // @[FPU.scala 882:28]
  wire [64:0] dfma_io_in_bits_in1; // @[FPU.scala 882:28]
  wire [64:0] dfma_io_in_bits_in2; // @[FPU.scala 882:28]
  wire [64:0] dfma_io_in_bits_in3; // @[FPU.scala 882:28]
  wire [64:0] dfma_io_out_bits_data; // @[FPU.scala 882:28]
  wire [4:0] dfma_io_out_bits_exc; // @[FPU.scala 882:28]
  wire [29:0] dfma_io_covSum; // @[FPU.scala 882:28]
  wire  dfma_metaAssert; // @[FPU.scala 882:28]
  wire  dfma_metaReset; // @[FPU.scala 882:28]
  wire  dfma_fma_halt; // @[FPU.scala 882:28]
  wire  divSqrt_clock; // @[FPU.scala 986:55]
  wire  divSqrt_reset; // @[FPU.scala 986:55]
  wire  divSqrt_io_inReady; // @[FPU.scala 986:55]
  wire  divSqrt_io_inValid; // @[FPU.scala 986:55]
  wire  divSqrt_io_sqrtOp; // @[FPU.scala 986:55]
  wire [32:0] divSqrt_io_a; // @[FPU.scala 986:55]
  wire [32:0] divSqrt_io_b; // @[FPU.scala 986:55]
  wire [2:0] divSqrt_io_roundingMode; // @[FPU.scala 986:55]
  wire  divSqrt_io_outValid_div; // @[FPU.scala 986:55]
  wire  divSqrt_io_outValid_sqrt; // @[FPU.scala 986:55]
  wire [32:0] divSqrt_io_out; // @[FPU.scala 986:55]
  wire [4:0] divSqrt_io_exceptionFlags; // @[FPU.scala 986:55]
  wire [29:0] divSqrt_io_covSum; // @[FPU.scala 986:55]
  wire  divSqrt_metaAssert; // @[FPU.scala 986:55]
  wire  divSqrt_metaReset; // @[FPU.scala 986:55]
  wire  divSqrt_divSqrtRecFNToRaw_halt; // @[FPU.scala 986:55]
  wire  divSqrt_1_clock; // @[FPU.scala 986:55]
  wire  divSqrt_1_reset; // @[FPU.scala 986:55]
  wire  divSqrt_1_io_inReady; // @[FPU.scala 986:55]
  wire  divSqrt_1_io_inValid; // @[FPU.scala 986:55]
  wire  divSqrt_1_io_sqrtOp; // @[FPU.scala 986:55]
  wire [64:0] divSqrt_1_io_a; // @[FPU.scala 986:55]
  wire [64:0] divSqrt_1_io_b; // @[FPU.scala 986:55]
  wire [2:0] divSqrt_1_io_roundingMode; // @[FPU.scala 986:55]
  wire  divSqrt_1_io_outValid_div; // @[FPU.scala 986:55]
  wire  divSqrt_1_io_outValid_sqrt; // @[FPU.scala 986:55]
  wire [64:0] divSqrt_1_io_out; // @[FPU.scala 986:55]
  wire [4:0] divSqrt_1_io_exceptionFlags; // @[FPU.scala 986:55]
  wire [29:0] divSqrt_1_io_covSum; // @[FPU.scala 986:55]
  wire  divSqrt_1_metaAssert; // @[FPU.scala 986:55]
  wire  divSqrt_1_metaReset; // @[FPU.scala 986:55]
  wire  divSqrt_1_divSqrtRecFNToRaw_halt; // @[FPU.scala 986:55]
  reg  ex_reg_valid; // @[FPU.scala 746:25]
  reg [31:0] _RAND_1;
  reg [31:0] ex_reg_inst; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg  ex_reg_ctrl_ren2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg  ex_reg_ctrl_ren3; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg  ex_reg_ctrl_swap23; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg [1:0] ex_reg_ctrl_typeTagIn; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg [1:0] ex_reg_ctrl_typeTagOut; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7;
  reg  ex_reg_ctrl_fromint; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8;
  reg  ex_reg_ctrl_toint; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  reg  ex_reg_ctrl_fastpipe; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10;
  reg  ex_reg_ctrl_fma; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11;
  reg  ex_reg_ctrl_div; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12;
  reg  ex_reg_ctrl_sqrt; // @[Reg.scala 15:16]
  reg [31:0] _RAND_13;
  reg  ex_reg_ctrl_wflags; // @[Reg.scala 15:16]
  reg [31:0] _RAND_14;
  reg [4:0] ex_ra_0; // @[FPU.scala 749:31]
  reg [31:0] _RAND_15;
  reg [4:0] ex_ra_1; // @[FPU.scala 749:31]
  reg [31:0] _RAND_16;
  reg [4:0] ex_ra_2; // @[FPU.scala 749:31]
  reg [31:0] _RAND_17;
  reg  load_wb; // @[FPU.scala 752:20]
  reg [31:0] _RAND_18;
  wire [1:0] _load_wb_typeTag_T_2; // @[FPU.scala 753:58]
  reg [1:0] load_wb_typeTag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_19;
  reg [63:0] load_wb_data; // @[Reg.scala 15:16]
  reg [63:0] _RAND_20;
  reg [4:0] load_wb_tag; // @[Reg.scala 15:16]
  reg [31:0] _RAND_21;
  reg  mem_reg_valid; // @[FPU.scala 763:30]
  reg [31:0] _RAND_22;
  wire  killm; // @[FPU.scala 764:25]
  wire  _killx_T; // @[FPU.scala 768:41]
  wire  killx; // @[FPU.scala 768:24]
  wire  _mem_reg_valid_T_1; // @[FPU.scala 769:33]
  reg [31:0] mem_reg_inst; // @[Reg.scala 15:16]
  reg [31:0] _RAND_23;
  wire  wb_reg_valid_x7; // @[FPU.scala 771:45]
  reg  wb_reg_valid; // @[FPU.scala 771:25]
  reg [31:0] _RAND_24;
  reg [1:0] mem_ctrl_typeTagOut; // @[Reg.scala 15:16]
  reg [31:0] _RAND_25;
  reg  mem_ctrl_fromint; // @[Reg.scala 15:16]
  reg [31:0] _RAND_26;
  reg  mem_ctrl_toint; // @[Reg.scala 15:16]
  reg [31:0] _RAND_27;
  reg  mem_ctrl_fastpipe; // @[Reg.scala 15:16]
  reg [31:0] _RAND_28;
  reg  mem_ctrl_fma; // @[Reg.scala 15:16]
  reg [31:0] _RAND_29;
  reg  mem_ctrl_div; // @[Reg.scala 15:16]
  reg [31:0] _RAND_30;
  reg  mem_ctrl_sqrt; // @[Reg.scala 15:16]
  reg [31:0] _RAND_31;
  reg  mem_ctrl_wflags; // @[Reg.scala 15:16]
  reg [31:0] _RAND_32;
  reg  wb_ctrl_toint; // @[Reg.scala 15:16]
  reg [31:0] _RAND_33;
  wire  wdata_truncIdx; // @[package.scala 31:49]
  wire [63:0] _wdata_T_1; // @[package.scala 32:76]
  wire [63:0] _wdata_T_2; // @[FPU.scala 426:23]
  wire  wdata_rawIn_sign; // @[rawFloatFromFN.scala 46:22]
  wire [10:0] wdata_rawIn_expIn; // @[rawFloatFromFN.scala 47:23]
  wire [51:0] wdata_rawIn_fractIn; // @[rawFloatFromFN.scala 48:25]
  wire  wdata_rawIn_isZeroExpIn; // @[rawFloatFromFN.scala 50:34]
  wire  wdata_rawIn_isZeroFractIn; // @[rawFloatFromFN.scala 51:38]
  wire [5:0] _wdata_rawIn_normDist_T_52; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_53; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_54; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_55; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_56; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_57; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_58; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_59; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_60; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_61; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_62; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_63; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_64; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_65; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_66; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_67; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_68; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_69; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_70; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_71; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_72; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_73; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_74; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_75; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_76; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_77; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_78; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_79; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_80; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_81; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_82; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_83; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_84; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_85; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_86; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_87; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_88; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_89; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_90; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_91; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_92; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_93; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_94; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_95; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_96; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_97; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_98; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_99; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_100; // @[Mux.scala 47:69]
  wire [5:0] _wdata_rawIn_normDist_T_101; // @[Mux.scala 47:69]
  wire [5:0] wdata_rawIn_normDist; // @[Mux.scala 47:69]
  wire [114:0] _GEN_168; // @[rawFloatFromFN.scala 54:36]
  wire [114:0] _wdata_rawIn_subnormFract_T; // @[rawFloatFromFN.scala 54:36]
  wire [51:0] wdata_rawIn_subnormFract; // @[rawFloatFromFN.scala 54:64]
  wire [11:0] _GEN_169; // @[rawFloatFromFN.scala 57:26]
  wire [11:0] _wdata_rawIn_adjustedExp_T; // @[rawFloatFromFN.scala 57:26]
  wire [11:0] _wdata_rawIn_adjustedExp_T_1; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _wdata_rawIn_adjustedExp_T_2; // @[rawFloatFromFN.scala 60:27]
  wire [10:0] _GEN_170; // @[rawFloatFromFN.scala 60:22]
  wire [10:0] _wdata_rawIn_adjustedExp_T_3; // @[rawFloatFromFN.scala 60:22]
  wire [11:0] _GEN_171; // @[rawFloatFromFN.scala 59:15]
  wire [11:0] wdata_rawIn_adjustedExp; // @[rawFloatFromFN.scala 59:15]
  wire  wdata_rawIn_isZero; // @[rawFloatFromFN.scala 62:34]
  wire  wdata_rawIn_isSpecial; // @[rawFloatFromFN.scala 63:62]
  wire  wdata_rawIn__isNaN; // @[rawFloatFromFN.scala 66:33]
  wire [12:0] wdata_rawIn__sExp; // @[rawFloatFromFN.scala 70:48]
  wire  wdata_rawIn_out_sig_hi_lo; // @[rawFloatFromFN.scala 72:29]
  wire [51:0] wdata_rawIn_out_sig_lo; // @[rawFloatFromFN.scala 72:42]
  wire [53:0] wdata_rawIn__sig; // @[Cat.scala 30:58]
  wire [2:0] _wdata_T_4; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_172; // @[recFNFromFN.scala 48:79]
  wire [2:0] wdata_hi_lo; // @[recFNFromFN.scala 48:79]
  wire [8:0] wdata_lo_hi; // @[recFNFromFN.scala 50:23]
  wire [51:0] wdata_lo_lo; // @[recFNFromFN.scala 51:22]
  wire [64:0] _wdata_T_6; // @[Cat.scala 30:58]
  wire  wdata_rawIn_sign_1; // @[rawFloatFromFN.scala 46:22]
  wire [7:0] wdata_rawIn_expIn_1; // @[rawFloatFromFN.scala 47:23]
  wire [22:0] wdata_rawIn_fractIn_1; // @[rawFloatFromFN.scala 48:25]
  wire  wdata_rawIn_isZeroExpIn_1; // @[rawFloatFromFN.scala 50:34]
  wire  wdata_rawIn_isZeroFractIn_1; // @[rawFloatFromFN.scala 51:38]
  wire [4:0] _wdata_rawIn_normDist_T_125; // @[Mux.scala 47:69]
  wire [4:0] _wdata_rawIn_normDist_T_126; // @[Mux.scala 47:69]
  wire [4:0] _wdata_rawIn_normDist_T_127; // @[Mux.scala 47:69]
  wire [4:0] _wdata_rawIn_normDist_T_128; // @[Mux.scala 47:69]
  wire [4:0] _wdata_rawIn_normDist_T_129; // @[Mux.scala 47:69]
  wire [4:0] _wdata_rawIn_normDist_T_130; // @[Mux.scala 47:69]
  wire [4:0] _wdata_rawIn_normDist_T_131; // @[Mux.scala 47:69]
  wire [4:0] _wdata_rawIn_normDist_T_132; // @[Mux.scala 47:69]
  wire [4:0] _wdata_rawIn_normDist_T_133; // @[Mux.scala 47:69]
  wire [4:0] _wdata_rawIn_normDist_T_134; // @[Mux.scala 47:69]
  wire [4:0] _wdata_rawIn_normDist_T_135; // @[Mux.scala 47:69]
  wire [4:0] _wdata_rawIn_normDist_T_136; // @[Mux.scala 47:69]
  wire [4:0] _wdata_rawIn_normDist_T_137; // @[Mux.scala 47:69]
  wire [4:0] _wdata_rawIn_normDist_T_138; // @[Mux.scala 47:69]
  wire [4:0] _wdata_rawIn_normDist_T_139; // @[Mux.scala 47:69]
  wire [4:0] _wdata_rawIn_normDist_T_140; // @[Mux.scala 47:69]
  wire [4:0] _wdata_rawIn_normDist_T_141; // @[Mux.scala 47:69]
  wire [4:0] _wdata_rawIn_normDist_T_142; // @[Mux.scala 47:69]
  wire [4:0] _wdata_rawIn_normDist_T_143; // @[Mux.scala 47:69]
  wire [4:0] _wdata_rawIn_normDist_T_144; // @[Mux.scala 47:69]
  wire [4:0] _wdata_rawIn_normDist_T_145; // @[Mux.scala 47:69]
  wire [4:0] wdata_rawIn_normDist_1; // @[Mux.scala 47:69]
  wire [53:0] _GEN_173; // @[rawFloatFromFN.scala 54:36]
  wire [53:0] _wdata_rawIn_subnormFract_T_2; // @[rawFloatFromFN.scala 54:36]
  wire [22:0] wdata_rawIn_subnormFract_1; // @[rawFloatFromFN.scala 54:64]
  wire [8:0] _GEN_174; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _wdata_rawIn_adjustedExp_T_5; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _wdata_rawIn_adjustedExp_T_6; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _wdata_rawIn_adjustedExp_T_7; // @[rawFloatFromFN.scala 60:27]
  wire [7:0] _GEN_175; // @[rawFloatFromFN.scala 60:22]
  wire [7:0] _wdata_rawIn_adjustedExp_T_8; // @[rawFloatFromFN.scala 60:22]
  wire [8:0] _GEN_176; // @[rawFloatFromFN.scala 59:15]
  wire [8:0] wdata_rawIn_adjustedExp_1; // @[rawFloatFromFN.scala 59:15]
  wire  wdata_rawIn_isZero_1; // @[rawFloatFromFN.scala 62:34]
  wire  wdata_rawIn_isSpecial_1; // @[rawFloatFromFN.scala 63:62]
  wire  wdata_rawIn_1_isNaN; // @[rawFloatFromFN.scala 66:33]
  wire [9:0] wdata_rawIn_1_sExp; // @[rawFloatFromFN.scala 70:48]
  wire  wdata_rawIn_out_sig_hi_lo_1; // @[rawFloatFromFN.scala 72:29]
  wire [22:0] wdata_rawIn_out_sig_lo_1; // @[rawFloatFromFN.scala 72:42]
  wire [24:0] wdata_rawIn_1_sig; // @[Cat.scala 30:58]
  wire [2:0] _wdata_T_8; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_177; // @[recFNFromFN.scala 48:79]
  wire [2:0] wdata_hi_lo_1; // @[recFNFromFN.scala 48:79]
  wire [5:0] wdata_lo_hi_1; // @[recFNFromFN.scala 50:23]
  wire [22:0] wdata_lo_lo_1; // @[recFNFromFN.scala 51:22]
  wire [32:0] _wdata_T_10; // @[Cat.scala 30:58]
  wire [3:0] wdata_swizzledNaN_hi_hi_hi; // @[FPU.scala 332:8]
  wire  wdata_swizzledNaN_hi_hi_lo; // @[FPU.scala 333:42]
  wire [6:0] wdata_swizzledNaN_hi_lo_hi; // @[FPU.scala 334:8]
  wire  wdata_swizzledNaN_hi_lo_lo; // @[FPU.scala 335:8]
  wire  wdata_swizzledNaN_lo_hi_lo; // @[FPU.scala 337:8]
  wire [30:0] wdata_swizzledNaN_lo_lo; // @[FPU.scala 338:8]
  wire [64:0] wdata_swizzledNaN; // @[Cat.scala 30:58]
  wire  _wdata_T_12; // @[FPU.scala 243:56]
  wire [64:0] wdata; // @[FPU.scala 339:8]
  wire  _curOK_T_1; // @[FPU.scala 243:56]
  wire  _curOK_T_5; // @[FPU.scala 380:96]
  wire  _curOK_T_6; // @[FPU.scala 380:55]
  wire  curOK; // @[FPU.scala 380:31]
  wire  _T_2; // @[FPU.scala 800:11]
  wire [5:0] _GEN_178; // @[FPU.scala 802:57]
  wire [5:0] _T_5; // @[FPU.scala 802:57]
  wire  _T_11; // @[FPU.scala 817:29]
  wire  _ex_rm_T_1; // @[FPU.scala 821:38]
  wire  _sfma_io_in_valid_T; // @[FPU.scala 845:33]
  wire  _sfma_io_in_valid_T_1; // @[FPU.scala 845:70]
  wire  sfma_io_in_bits_req_in1_unswizzled_hi_hi; // @[FPU.scala 352:14]
  wire  sfma_io_in_bits_req_in1_unswizzled_hi_lo; // @[FPU.scala 353:14]
  wire [30:0] sfma_io_in_bits_req_in1_unswizzled_lo; // @[FPU.scala 354:14]
  wire [32:0] sfma_io_in_bits_req_in1_floats_0; // @[Cat.scala 30:58]
  wire  sfma_io_in_bits_req_in1_isbox; // @[FPU.scala 327:84]
  wire [32:0] _sfma_io_in_bits_req_in1_T; // @[FPU.scala 367:31]
  wire [32:0] _sfma_io_in_bits_req_in1_T_1; // @[FPU.scala 367:26]
  wire  sfma_io_in_bits_req_in2_unswizzled_hi_hi; // @[FPU.scala 352:14]
  wire  sfma_io_in_bits_req_in2_unswizzled_hi_lo; // @[FPU.scala 353:14]
  wire [30:0] sfma_io_in_bits_req_in2_unswizzled_lo; // @[FPU.scala 354:14]
  wire [32:0] sfma_io_in_bits_req_in2_floats_0; // @[Cat.scala 30:58]
  wire  sfma_io_in_bits_req_in2_isbox; // @[FPU.scala 327:84]
  wire [32:0] _sfma_io_in_bits_req_in2_T; // @[FPU.scala 367:31]
  wire [32:0] _sfma_io_in_bits_req_in2_T_1; // @[FPU.scala 367:26]
  wire  sfma_io_in_bits_req_in3_unswizzled_hi_hi; // @[FPU.scala 352:14]
  wire  sfma_io_in_bits_req_in3_unswizzled_hi_lo; // @[FPU.scala 353:14]
  wire [30:0] sfma_io_in_bits_req_in3_unswizzled_lo; // @[FPU.scala 354:14]
  wire [32:0] sfma_io_in_bits_req_in3_floats_0; // @[Cat.scala 30:58]
  wire  sfma_io_in_bits_req_in3_isbox; // @[FPU.scala 327:84]
  wire [32:0] _sfma_io_in_bits_req_in3_T; // @[FPU.scala 367:31]
  wire [32:0] _sfma_io_in_bits_req_in3_T_1; // @[FPU.scala 367:26]
  wire  _sfma_io_in_bits_req_fmaCmd_T_3; // @[FPU.scala 833:53]
  wire [1:0] _GEN_179; // @[FPU.scala 833:36]
  wire  _fpiu_io_in_valid_T; // @[FPU.scala 849:51]
  wire  _fpiu_io_in_valid_T_1; // @[FPU.scala 849:66]
  wire  _fpiu_io_in_valid_T_2; // @[FPU.scala 849:103]
  wire  _fpiu_io_in_valid_T_3; // @[FPU.scala 849:82]
  wire  fpiu_io_in_bits_req_in1_hi_hi; // @[FPU.scala 268:17]
  wire [22:0] fpiu_io_in_bits_req_in1_fractIn; // @[FPU.scala 269:20]
  wire [8:0] fpiu_io_in_bits_req_in1_expIn; // @[FPU.scala 270:18]
  wire [75:0] _fpiu_io_in_bits_req_in1_fractOut_T; // @[FPU.scala 271:28]
  wire [51:0] fpiu_io_in_bits_req_in1_lo; // @[FPU.scala 271:38]
  wire [2:0] fpiu_io_in_bits_req_in1_expOut_hi; // @[FPU.scala 273:26]
  wire [11:0] _GEN_180; // @[FPU.scala 274:31]
  wire [11:0] _fpiu_io_in_bits_req_in1_expOut_commonCase_T_1; // @[FPU.scala 274:31]
  wire [11:0] fpiu_io_in_bits_req_in1_expOut_commonCase; // @[FPU.scala 274:48]
  wire  _fpiu_io_in_bits_req_in1_expOut_T; // @[FPU.scala 275:19]
  wire  _fpiu_io_in_bits_req_in1_expOut_T_1; // @[FPU.scala 275:36]
  wire  _fpiu_io_in_bits_req_in1_expOut_T_2; // @[FPU.scala 275:25]
  wire [8:0] fpiu_io_in_bits_req_in1_expOut_lo; // @[FPU.scala 275:65]
  wire [11:0] _fpiu_io_in_bits_req_in1_expOut_T_3; // @[Cat.scala 30:58]
  wire [11:0] fpiu_io_in_bits_req_in1_hi_lo; // @[FPU.scala 275:10]
  wire [64:0] fpiu_io_in_bits_req_in1_floats_0; // @[Cat.scala 30:58]
  wire  fpiu_io_in_bits_req_in1_truncIdx; // @[package.scala 31:49]
  wire  _fpiu_io_in_bits_req_in1_T_1; // @[package.scala 32:76]
  wire [64:0] _fpiu_io_in_bits_req_in1_T_3; // @[package.scala 32:76]
  wire  fpiu_io_in_bits_req_in2_hi_hi; // @[FPU.scala 268:17]
  wire [22:0] fpiu_io_in_bits_req_in2_fractIn; // @[FPU.scala 269:20]
  wire [8:0] fpiu_io_in_bits_req_in2_expIn; // @[FPU.scala 270:18]
  wire [75:0] _fpiu_io_in_bits_req_in2_fractOut_T; // @[FPU.scala 271:28]
  wire [51:0] fpiu_io_in_bits_req_in2_lo; // @[FPU.scala 271:38]
  wire [2:0] fpiu_io_in_bits_req_in2_expOut_hi; // @[FPU.scala 273:26]
  wire [11:0] _GEN_181; // @[FPU.scala 274:31]
  wire [11:0] _fpiu_io_in_bits_req_in2_expOut_commonCase_T_1; // @[FPU.scala 274:31]
  wire [11:0] fpiu_io_in_bits_req_in2_expOut_commonCase; // @[FPU.scala 274:48]
  wire  _fpiu_io_in_bits_req_in2_expOut_T; // @[FPU.scala 275:19]
  wire  _fpiu_io_in_bits_req_in2_expOut_T_1; // @[FPU.scala 275:36]
  wire  _fpiu_io_in_bits_req_in2_expOut_T_2; // @[FPU.scala 275:25]
  wire [8:0] fpiu_io_in_bits_req_in2_expOut_lo; // @[FPU.scala 275:65]
  wire [11:0] _fpiu_io_in_bits_req_in2_expOut_T_3; // @[Cat.scala 30:58]
  wire [11:0] fpiu_io_in_bits_req_in2_hi_lo; // @[FPU.scala 275:10]
  wire [64:0] fpiu_io_in_bits_req_in2_floats_0; // @[Cat.scala 30:58]
  wire  _fpiu_io_in_bits_req_in2_T_1; // @[package.scala 32:76]
  wire [64:0] _fpiu_io_in_bits_req_in2_T_3; // @[package.scala 32:76]
  wire [64:0] _ifpu_io_in_bits_in1_T; // @[FPU.scala 861:29]
  reg [4:0] divSqrt_waddr; // @[FPU.scala 870:26]
  reg [31:0] _RAND_34;
  wire  _dfma_io_in_valid_T_1; // @[FPU.scala 883:78]
  wire  _memLatencyMask_T_2; // @[FPU.scala 880:72]
  wire  _memLatencyMask_T_3; // @[FPU.scala 880:56]
  wire [1:0] _memLatencyMask_T_4; // @[FPU.scala 895:23]
  wire  _memLatencyMask_T_5; // @[FPU.scala 885:78]
  wire  _memLatencyMask_T_6; // @[FPU.scala 885:62]
  wire [2:0] _memLatencyMask_T_7; // @[FPU.scala 895:23]
  wire  _memLatencyMask_T_8; // @[FPU.scala 895:78]
  wire [1:0] _GEN_188; // @[FPU.scala 895:78]
  wire [1:0] _memLatencyMask_T_9; // @[FPU.scala 895:78]
  wire [2:0] _GEN_189; // @[FPU.scala 895:78]
  wire [2:0] memLatencyMask; // @[FPU.scala 895:78]
  reg [2:0] wen; // @[FPU.scala 909:16]
  reg [31:0] _RAND_35;
  reg [4:0] wbInfo_0_rd; // @[FPU.scala 910:19]
  reg [31:0] _RAND_36;
  reg  wbInfo_0_typeTag; // @[FPU.scala 910:19]
  reg [31:0] _RAND_37;
  reg [1:0] wbInfo_0_pipeid; // @[FPU.scala 910:19]
  reg [31:0] _RAND_38;
  reg [4:0] wbInfo_1_rd; // @[FPU.scala 910:19]
  reg [31:0] _RAND_39;
  reg  wbInfo_1_typeTag; // @[FPU.scala 910:19]
  reg [31:0] _RAND_40;
  reg [1:0] wbInfo_1_pipeid; // @[FPU.scala 910:19]
  reg [31:0] _RAND_41;
  reg [4:0] wbInfo_2_rd; // @[FPU.scala 910:19]
  reg [31:0] _RAND_42;
  reg  wbInfo_2_typeTag; // @[FPU.scala 910:19]
  reg [31:0] _RAND_43;
  reg [1:0] wbInfo_2_pipeid; // @[FPU.scala 910:19]
  reg [31:0] _RAND_44;
  wire  _mem_wen_T; // @[FPU.scala 911:48]
  wire  _mem_wen_T_1; // @[FPU.scala 911:69]
  wire  mem_wen; // @[FPU.scala 911:31]
  wire [1:0] _write_port_busy_T; // @[FPU.scala 895:23]
  wire [1:0] _write_port_busy_T_1; // @[FPU.scala 895:23]
  wire  _write_port_busy_T_3; // @[FPU.scala 880:56]
  wire [2:0] _write_port_busy_T_4; // @[FPU.scala 895:23]
  wire  _write_port_busy_T_6; // @[FPU.scala 885:62]
  wire [3:0] _write_port_busy_T_7; // @[FPU.scala 895:23]
  wire [1:0] _write_port_busy_T_8; // @[FPU.scala 895:78]
  wire [2:0] _GEN_190; // @[FPU.scala 895:78]
  wire [2:0] _write_port_busy_T_9; // @[FPU.scala 895:78]
  wire [3:0] _GEN_191; // @[FPU.scala 895:78]
  wire [3:0] _write_port_busy_T_10; // @[FPU.scala 895:78]
  wire [3:0] _GEN_192; // @[FPU.scala 912:62]
  wire [3:0] _write_port_busy_T_11; // @[FPU.scala 912:62]
  wire  _write_port_busy_T_12; // @[FPU.scala 912:89]
  wire  _write_port_busy_T_13; // @[FPU.scala 912:43]
  wire [2:0] _write_port_busy_T_14; // @[FPU.scala 895:23]
  wire [2:0] _write_port_busy_T_15; // @[FPU.scala 895:23]
  wire [3:0] _write_port_busy_T_18; // @[FPU.scala 895:23]
  wire [4:0] _write_port_busy_T_21; // @[FPU.scala 895:23]
  wire [2:0] _write_port_busy_T_22; // @[FPU.scala 895:78]
  wire [3:0] _GEN_193; // @[FPU.scala 895:78]
  wire [3:0] _write_port_busy_T_23; // @[FPU.scala 895:78]
  wire [4:0] _GEN_194; // @[FPU.scala 895:78]
  wire [4:0] _write_port_busy_T_24; // @[FPU.scala 895:78]
  wire [4:0] _GEN_195; // @[FPU.scala 912:101]
  wire [4:0] _write_port_busy_T_25; // @[FPU.scala 912:101]
  wire  _write_port_busy_T_26; // @[FPU.scala 912:128]
  wire  _write_port_busy_T_27; // @[FPU.scala 912:93]
  reg  write_port_busy; // @[Reg.scala 15:16]
  reg [31:0] _RAND_45;
  wire  _GEN_114; // @[FPU.scala 916:21]
  wire  _GEN_118; // @[FPU.scala 916:21]
  wire [2:0] _GEN_196; // @[FPU.scala 921:23]
  wire [2:0] _wen_T_2; // @[FPU.scala 921:23]
  wire  _T_20; // @[FPU.scala 924:30]
  wire [1:0] _wbInfo_0_pipeid_T_7; // @[FPU.scala 897:63]
  wire [1:0] _GEN_197; // @[FPU.scala 897:108]
  wire [1:0] _wbInfo_0_pipeid_T_9; // @[FPU.scala 897:108]
  wire [1:0] _wbInfo_0_pipeid_T_10; // @[FPU.scala 897:108]
  wire [1:0] _GEN_123; // @[FPU.scala 924:52]
  wire  _T_23; // @[FPU.scala 924:30]
  wire [1:0] _GEN_127; // @[FPU.scala 924:52]
  wire  _T_26; // @[FPU.scala 924:30]
  wire [1:0] _GEN_131; // @[FPU.scala 924:52]
  wire [1:0] _GEN_136; // @[FPU.scala 919:18]
  wire [1:0] _GEN_140; // @[FPU.scala 919:18]
  wire [1:0] _GEN_144; // @[FPU.scala 919:18]
  wire  divSqrt_typeTag; // @[FPU.scala 996:37]
  reg  divSqrt_killed; // @[FPU.scala 975:33]
  reg [31:0] _RAND_46;
  wire  _T_52; // @[FPU.scala 996:37]
  wire  _GEN_158; // @[FPU.scala 996:66]
  wire  divSqrt_wen; // @[FPU.scala 996:66]
  wire [4:0] waddr; // @[FPU.scala 933:18]
  wire  wtypeTag; // @[FPU.scala 934:21]
  wire  _wdata_T_13; // @[package.scala 32:86]
  wire [64:0] _wdata_T_14; // @[package.scala 32:76]
  wire  _wdata_T_15; // @[package.scala 32:86]
  wire [64:0] _wdata_T_16; // @[package.scala 32:76]
  wire  _wdata_T_17; // @[package.scala 32:86]
  wire [64:0] _wdata_T_18; // @[package.scala 32:76]
  wire  _divSqrt_wdata_T_1; // @[FPU.scala 243:56]
  wire [64:0] divSqrt_wdata_maskedNaN; // @[FPU.scala 408:25]
  wire [64:0] _divSqrt_wdata_T_2; // @[FPU.scala 409:10]
  wire [32:0] _GEN_159; // @[FPU.scala 996:66]
  wire [64:0] divSqrt_wdata; // @[FPU.scala 996:66]
  wire [64:0] _wdata_T_19; // @[FPU.scala 935:22]
  wire  wdata_opts_bigger_swizzledNaN_hi_hi_lo; // @[FPU.scala 333:42]
  wire  wdata_opts_bigger_swizzledNaN_hi_lo_lo; // @[FPU.scala 335:8]
  wire  wdata_opts_bigger_swizzledNaN_lo_hi_lo; // @[FPU.scala 337:8]
  wire [30:0] wdata_opts_bigger_swizzledNaN_lo_lo; // @[FPU.scala 338:8]
  wire [64:0] wdata_opts_bigger_swizzledNaN; // @[Cat.scala 30:58]
  wire  _wdata_opts_bigger_T; // @[FPU.scala 243:56]
  wire [64:0] wdata_opts_bigger; // @[FPU.scala 339:8]
  wire [64:0] wdata_1; // @[package.scala 32:76]
  wire [4:0] _wexc_T_1; // @[package.scala 32:76]
  wire [4:0] _wexc_T_3; // @[package.scala 32:76]
  wire [4:0] wexc; // @[package.scala 32:76]
  wire  frfWriteBundle_1_wrenf; // @[FPU.scala 937:35]
  wire  unswizzled_hi_hi_1; // @[FPU.scala 376:10]
  wire  unswizzled_hi_lo_1; // @[FPU.scala 377:10]
  wire [30:0] unswizzled_lo_1; // @[FPU.scala 378:10]
  wire [32:0] unswizzled_1; // @[Cat.scala 30:58]
  wire  _curOK_T_8; // @[FPU.scala 243:56]
  wire  _curOK_T_12; // @[FPU.scala 380:96]
  wire  _curOK_T_13; // @[FPU.scala 380:55]
  wire  curOK_1; // @[FPU.scala 380:31]
  wire  _T_33; // @[FPU.scala 938:11]
  wire [5:0] _GEN_200; // @[FPU.scala 941:45]
  wire [5:0] _T_36; // @[FPU.scala 941:45]
  wire [11:0] unrecoded_rawIn_exp; // @[rawFloatFromRecFN.scala 50:21]
  wire  unrecoded_rawIn_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  unrecoded_rawIn_isSpecial; // @[rawFloatFromRecFN.scala 52:54]
  wire  unrecoded_rawIn__isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  unrecoded_rawIn__isInf; // @[rawFloatFromRecFN.scala 56:33]
  wire  unrecoded_rawIn__sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [12:0] unrecoded_rawIn__sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire  unrecoded_rawIn_out_sig_hi_lo; // @[rawFloatFromRecFN.scala 60:39]
  wire [51:0] unrecoded_rawIn_out_sig_lo; // @[rawFloatFromRecFN.scala 60:51]
  wire [53:0] unrecoded_rawIn__sig; // @[Cat.scala 30:58]
  wire  unrecoded_isSubnormal; // @[fNFromRecFN.scala 50:39]
  wire [5:0] unrecoded_denormShiftDist; // @[fNFromRecFN.scala 51:39]
  wire [52:0] _unrecoded_denormFract_T_1; // @[fNFromRecFN.scala 52:42]
  wire [51:0] unrecoded_denormFract; // @[fNFromRecFN.scala 52:60]
  wire [10:0] _unrecoded_expOut_T_2; // @[fNFromRecFN.scala 57:45]
  wire [10:0] _unrecoded_expOut_T_3; // @[fNFromRecFN.scala 55:16]
  wire  _unrecoded_expOut_T_4; // @[fNFromRecFN.scala 59:44]
  wire [10:0] _unrecoded_expOut_T_6; // @[Bitwise.scala 72:12]
  wire [10:0] unrecoded_hi_lo; // @[fNFromRecFN.scala 59:15]
  wire [51:0] _unrecoded_fractOut_T_1; // @[fNFromRecFN.scala 63:20]
  wire [51:0] unrecoded_lo; // @[fNFromRecFN.scala 61:16]
  wire [63:0] unrecoded; // @[Cat.scala 30:58]
  wire [8:0] prevUnrecoded_rawIn_exp; // @[rawFloatFromRecFN.scala 50:21]
  wire  prevUnrecoded_rawIn_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  prevUnrecoded_rawIn_isSpecial; // @[rawFloatFromRecFN.scala 52:54]
  wire  prevUnrecoded_rawIn__isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  prevUnrecoded_rawIn__isInf; // @[rawFloatFromRecFN.scala 56:33]
  wire  prevUnrecoded_rawIn__sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [9:0] prevUnrecoded_rawIn__sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire  prevUnrecoded_rawIn_out_sig_hi_lo; // @[rawFloatFromRecFN.scala 60:39]
  wire [22:0] prevUnrecoded_rawIn_out_sig_lo; // @[rawFloatFromRecFN.scala 60:51]
  wire [24:0] prevUnrecoded_rawIn__sig; // @[Cat.scala 30:58]
  wire  prevUnrecoded_isSubnormal; // @[fNFromRecFN.scala 50:39]
  wire [4:0] prevUnrecoded_denormShiftDist; // @[fNFromRecFN.scala 51:39]
  wire [23:0] _prevUnrecoded_denormFract_T_1; // @[fNFromRecFN.scala 52:42]
  wire [22:0] prevUnrecoded_denormFract; // @[fNFromRecFN.scala 52:60]
  wire [7:0] _prevUnrecoded_expOut_T_2; // @[fNFromRecFN.scala 57:45]
  wire [7:0] _prevUnrecoded_expOut_T_3; // @[fNFromRecFN.scala 55:16]
  wire  _prevUnrecoded_expOut_T_4; // @[fNFromRecFN.scala 59:44]
  wire [7:0] _prevUnrecoded_expOut_T_6; // @[Bitwise.scala 72:12]
  wire [7:0] prevUnrecoded_hi_lo; // @[fNFromRecFN.scala 59:15]
  wire [22:0] _prevUnrecoded_fractOut_T_1; // @[fNFromRecFN.scala 63:20]
  wire [22:0] prevUnrecoded_lo; // @[fNFromRecFN.scala 61:16]
  wire [31:0] prevUnrecoded; // @[Cat.scala 30:58]
  wire [31:0] hi; // @[FPU.scala 441:21]
  wire [31:0] lo; // @[FPU.scala 441:44]
  wire [63:0] _T_40; // @[Cat.scala 30:58]
  wire  wb_toint_valid; // @[FPU.scala 953:37]
  reg [4:0] wb_toint_exc; // @[Reg.scala 15:16]
  reg [31:0] _RAND_47;
  wire  _io_fcsr_flags_valid_T; // @[FPU.scala 955:41]
  wire [4:0] _io_fcsr_flags_bits_T; // @[FPU.scala 957:8]
  wire [4:0] _GEN_160; // @[FPU.scala 996:66]
  wire [4:0] divSqrt_flags; // @[FPU.scala 996:66]
  wire [4:0] _io_fcsr_flags_bits_T_1; // @[FPU.scala 958:8]
  wire [4:0] _io_fcsr_flags_bits_T_2; // @[FPU.scala 957:48]
  wire [4:0] _io_fcsr_flags_bits_T_4; // @[FPU.scala 959:8]
  wire  _divSqrt_write_port_busy_T; // @[FPU.scala 961:47]
  wire  _divSqrt_write_port_busy_T_1; // @[FPU.scala 961:72]
  wire  divSqrt_write_port_busy; // @[FPU.scala 961:65]
  wire  _io_fcsr_rdy_T; // @[FPU.scala 962:33]
  wire  _io_fcsr_rdy_T_1; // @[FPU.scala 962:68]
  wire  _io_fcsr_rdy_T_2; // @[FPU.scala 962:51]
  wire  _io_fcsr_rdy_T_4; // @[FPU.scala 962:87]
  wire  _io_fcsr_rdy_T_6; // @[FPU.scala 962:120]
  wire  _GEN_162; // @[FPU.scala 994:34]
  wire  divSqrt_inFlight; // @[FPU.scala 1004:27]
  wire  _io_fcsr_rdy_T_7; // @[FPU.scala 962:131]
  wire  _io_nack_mem_T; // @[FPU.scala 963:34]
  wire  _io_sboard_set_x27_T_3; // @[FPU.scala 966:96]
  reg  io_sboard_set_REG; // @[FPU.scala 966:55]
  reg [31:0] _RAND_48;
  wire  _io_sboard_clr_T_4; // @[FPU.scala 967:60]
  wire  _io_illegal_rm_T_1; // @[package.scala 15:47]
  wire  _io_illegal_rm_T_2; // @[package.scala 15:47]
  wire  _io_illegal_rm_T_3; // @[package.scala 72:59]
  wire  _io_illegal_rm_T_5; // @[FPU.scala 971:67]
  wire  _io_illegal_rm_T_6; // @[FPU.scala 971:87]
  wire  _io_illegal_rm_T_7; // @[FPU.scala 971:73]
  wire  _divSqrt_inValid_T_1; // @[FPU.scala 974:41]
  wire  divSqrt_inValid; // @[FPU.scala 974:76]
  wire  _divSqrt_killed_T; // @[FPU.scala 975:50]
  wire  divSqrt_io_a_hi_hi; // @[FPU.scala 268:17]
  wire [51:0] divSqrt_io_a_fractIn; // @[FPU.scala 269:20]
  wire [11:0] divSqrt_io_a_expIn; // @[FPU.scala 270:18]
  wire [75:0] _divSqrt_io_a_fractOut_T; // @[FPU.scala 271:28]
  wire [22:0] divSqrt_io_a_lo; // @[FPU.scala 271:38]
  wire [2:0] divSqrt_io_a_expOut_hi; // @[FPU.scala 273:26]
  wire [11:0] _divSqrt_io_a_expOut_commonCase_T_1; // @[FPU.scala 274:31]
  wire [11:0] divSqrt_io_a_expOut_commonCase; // @[FPU.scala 274:48]
  wire  _divSqrt_io_a_expOut_T; // @[FPU.scala 275:19]
  wire  _divSqrt_io_a_expOut_T_1; // @[FPU.scala 275:36]
  wire  _divSqrt_io_a_expOut_T_2; // @[FPU.scala 275:25]
  wire [5:0] divSqrt_io_a_expOut_lo; // @[FPU.scala 275:65]
  wire [8:0] _divSqrt_io_a_expOut_T_3; // @[Cat.scala 30:58]
  wire [8:0] divSqrt_io_a_hi_lo; // @[FPU.scala 275:10]
  wire [9:0] divSqrt_io_a_hi; // @[Cat.scala 30:58]
  wire  divSqrt_io_b_hi_hi; // @[FPU.scala 268:17]
  wire [51:0] divSqrt_io_b_fractIn; // @[FPU.scala 269:20]
  wire [11:0] divSqrt_io_b_expIn; // @[FPU.scala 270:18]
  wire [75:0] _divSqrt_io_b_fractOut_T; // @[FPU.scala 271:28]
  wire [22:0] divSqrt_io_b_lo; // @[FPU.scala 271:38]
  wire [2:0] divSqrt_io_b_expOut_hi; // @[FPU.scala 273:26]
  wire [11:0] _divSqrt_io_b_expOut_commonCase_T_1; // @[FPU.scala 274:31]
  wire [11:0] divSqrt_io_b_expOut_commonCase; // @[FPU.scala 274:48]
  wire  _divSqrt_io_b_expOut_T; // @[FPU.scala 275:19]
  wire  _divSqrt_io_b_expOut_T_1; // @[FPU.scala 275:36]
  wire  _divSqrt_io_b_expOut_T_2; // @[FPU.scala 275:25]
  wire [5:0] divSqrt_io_b_expOut_lo; // @[FPU.scala 275:65]
  wire [8:0] _divSqrt_io_b_expOut_T_3; // @[Cat.scala 30:58]
  wire [8:0] divSqrt_io_b_hi_lo; // @[FPU.scala 275:10]
  wire [9:0] divSqrt_io_b_hi; // @[Cat.scala 30:58]
  reg [19:0] FPU_state; // @[Register tracking FPU state]
  reg [31:0] _RAND_49;
  reg  FPU_cov [0:1048575]; // @[Coverage map for FPU]
  reg [31:0] _RAND_50;
  wire  FPU_cov_read_data; // @[Coverage map for FPU]
  wire [19:0] FPU_cov_read_addr; // @[Coverage map for FPU]
  wire  FPU_cov_write_data; // @[Coverage map for FPU]
  wire [19:0] FPU_cov_write_addr; // @[Coverage map for FPU]
  wire  FPU_cov_write_mask; // @[Coverage map for FPU]
  wire  FPU_cov_write_en; // @[Coverage map for FPU]
  reg [29:0] FPU_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_51;
  wire [16:0] wbInfo_0_typeTag_shl;
  wire [19:0] wbInfo_0_typeTag_pad;
  wire [2:0] wb_reg_valid_shl;
  wire [19:0] wb_reg_valid_pad;
  wire [7:0] mem_ctrl_sqrt_shl;
  wire [19:0] mem_ctrl_sqrt_pad;
  wire [19:0] divSqrt_killed_shl;
  wire [19:0] divSqrt_killed_pad;
  wire [8:0] ex_reg_ctrl_typeTagIn_shl;
  wire [19:0] ex_reg_ctrl_typeTagIn_pad;
  wire [2:0] ex_reg_ctrl_fromint_shl;
  wire [19:0] ex_reg_ctrl_fromint_pad;
  wire [8:0] mem_ctrl_typeTagOut_shl;
  wire [19:0] mem_ctrl_typeTagOut_pad;
  wire [7:0] wen_shl;
  wire [19:0] wen_pad;
  wire [11:0] wb_ctrl_toint_shl;
  wire [19:0] wb_ctrl_toint_pad;
  wire [18:0] ex_reg_ctrl_fastpipe_shl;
  wire [19:0] ex_reg_ctrl_fastpipe_pad;
  wire [14:0] write_port_busy_shl;
  wire [19:0] write_port_busy_pad;
  wire [5:0] mem_ctrl_fastpipe_shl;
  wire [19:0] mem_ctrl_fastpipe_pad;
  wire [14:0] ex_reg_ctrl_typeTagOut_shl;
  wire [19:0] ex_reg_ctrl_typeTagOut_pad;
  wire [17:0] mem_reg_valid_shl;
  wire [19:0] mem_reg_valid_pad;
  wire [13:0] mem_ctrl_div_shl;
  wire [19:0] mem_ctrl_div_pad;
  wire [11:0] wbInfo_0_pipeid_shl;
  wire [19:0] wbInfo_0_pipeid_pad;
  wire [1:0] mem_ctrl_toint_shl;
  wire [19:0] mem_ctrl_toint_pad;
  wire [4:0] ex_reg_ctrl_fma_shl;
  wire [19:0] ex_reg_ctrl_fma_pad;
  wire [3:0] ex_reg_valid_shl;
  wire [19:0] ex_reg_valid_pad;
  wire [10:0] mem_ctrl_fromint_shl;
  wire [19:0] mem_ctrl_fromint_pad;
  wire [2:0] mem_ctrl_fma_shl;
  wire [19:0] mem_ctrl_fma_pad;
  wire [19:0] FPU_xor7;
  wire [19:0] FPU_xor18;
  wire [19:0] FPU_xor8;
  wire [19:0] FPU_xor3;
  wire [19:0] FPU_xor9;
  wire [19:0] FPU_xor22;
  wire [19:0] FPU_xor10;
  wire [19:0] FPU_xor4;
  wire [19:0] FPU_xor1;
  wire [19:0] FPU_xor11;
  wire [19:0] FPU_xor26;
  wire [19:0] FPU_xor12;
  wire [19:0] FPU_xor5;
  wire [19:0] FPU_xor28;
  wire [19:0] FPU_xor13;
  wire [19:0] FPU_xor30;
  wire [19:0] FPU_xor14;
  wire [19:0] FPU_xor6;
  wire [19:0] FPU_xor2;
  wire [19:0] FPU_xor0;
  wire [29:0] fpiu_sum;
  wire [29:0] fp_decoder_sum;
  wire [29:0] ifpu_sum;
  wire [29:0] sfma_sum;
  wire [29:0] fpmu_sum;
  wire [29:0] divSqrt_1_sum;
  wire [29:0] dfma_sum;
  wire [29:0] divSqrt_sum;
  wire  stopEn0;
  wire  stopEn1;
  wire  ifpu_metaAssert_wire;
  wire  fpmu_metaAssert_wire;
  wire  fp_decoder_metaAssert_wire;
  wire  fpiu_metaAssert_wire;
  wire  divSqrt_1_metaAssert_wire;
  wire  divSqrt_metaAssert_wire;
  wire  dfma_metaAssert_wire;
  wire  sfma_metaAssert_wire;
  wire  FPU_or3;
  wire  FPU_or10;
  wire  FPU_or4;
  wire  FPU_or1;
  wire  FPU_or5;
  wire  FPU_or14;
  wire  FPU_or6;
  wire  FPU_or2;
  wire  FPU_or0;
  reg  FPU_metaAssert;
  reg [31:0] _RAND_52;
  FPUDecoder fp_decoder ( // @[FPU.scala 742:26]
    .io_inst(fp_decoder_io_inst),
    .io_sigs_wen(fp_decoder_io_sigs_wen),
    .io_sigs_ren1(fp_decoder_io_sigs_ren1),
    .io_sigs_ren2(fp_decoder_io_sigs_ren2),
    .io_sigs_ren3(fp_decoder_io_sigs_ren3),
    .io_sigs_swap12(fp_decoder_io_sigs_swap12),
    .io_sigs_swap23(fp_decoder_io_sigs_swap23),
    .io_sigs_typeTagIn(fp_decoder_io_sigs_typeTagIn),
    .io_sigs_typeTagOut(fp_decoder_io_sigs_typeTagOut),
    .io_sigs_fromint(fp_decoder_io_sigs_fromint),
    .io_sigs_toint(fp_decoder_io_sigs_toint),
    .io_sigs_fastpipe(fp_decoder_io_sigs_fastpipe),
    .io_sigs_fma(fp_decoder_io_sigs_fma),
    .io_sigs_div(fp_decoder_io_sigs_div),
    .io_sigs_sqrt(fp_decoder_io_sigs_sqrt),
    .io_sigs_wflags(fp_decoder_io_sigs_wflags),
    .io_covSum(fp_decoder_io_covSum),
    .metaAssert(fp_decoder_metaAssert)
  );
  FPUFMAPipe sfma ( // @[FPU.scala 844:20]
    .clock(sfma_clock),
    .reset(sfma_reset),
    .io_in_valid(sfma_io_in_valid),
    .io_in_bits_ren3(sfma_io_in_bits_ren3),
    .io_in_bits_swap23(sfma_io_in_bits_swap23),
    .io_in_bits_rm(sfma_io_in_bits_rm),
    .io_in_bits_fmaCmd(sfma_io_in_bits_fmaCmd),
    .io_in_bits_in1(sfma_io_in_bits_in1),
    .io_in_bits_in2(sfma_io_in_bits_in2),
    .io_in_bits_in3(sfma_io_in_bits_in3),
    .io_out_bits_data(sfma_io_out_bits_data),
    .io_out_bits_exc(sfma_io_out_bits_exc),
    .io_covSum(sfma_io_covSum),
    .metaAssert(sfma_metaAssert),
    .metaReset(sfma_metaReset),
    .fma_halt(sfma_fma_halt)
  );
  FPToInt fpiu ( // @[FPU.scala 848:20]
    .clock(fpiu_clock),
    .io_in_valid(fpiu_io_in_valid),
    .io_in_bits_ren2(fpiu_io_in_bits_ren2),
    .io_in_bits_typeTagIn(fpiu_io_in_bits_typeTagIn),
    .io_in_bits_typeTagOut(fpiu_io_in_bits_typeTagOut),
    .io_in_bits_wflags(fpiu_io_in_bits_wflags),
    .io_in_bits_rm(fpiu_io_in_bits_rm),
    .io_in_bits_typ(fpiu_io_in_bits_typ),
    .io_in_bits_fmt(fpiu_io_in_bits_fmt),
    .io_in_bits_in1(fpiu_io_in_bits_in1),
    .io_in_bits_in2(fpiu_io_in_bits_in2),
    .io_out_bits_in_rm(fpiu_io_out_bits_in_rm),
    .io_out_bits_in_in1(fpiu_io_out_bits_in_in1),
    .io_out_bits_in_in2(fpiu_io_out_bits_in_in2),
    .io_out_bits_lt(fpiu_io_out_bits_lt),
    .io_out_bits_store(fpiu_io_out_bits_store),
    .io_out_bits_toint(fpiu_io_out_bits_toint),
    .io_out_bits_exc(fpiu_io_out_bits_exc),
    .io_covSum(fpiu_io_covSum),
    .metaAssert(fpiu_metaAssert),
    .metaReset(fpiu_metaReset)
  );
  IntToFP ifpu ( // @[FPU.scala 858:20]
    .clock(ifpu_clock),
    .reset(ifpu_reset),
    .io_in_valid(ifpu_io_in_valid),
    .io_in_bits_typeTagIn(ifpu_io_in_bits_typeTagIn),
    .io_in_bits_wflags(ifpu_io_in_bits_wflags),
    .io_in_bits_rm(ifpu_io_in_bits_rm),
    .io_in_bits_typ(ifpu_io_in_bits_typ),
    .io_in_bits_in1(ifpu_io_in_bits_in1),
    .io_out_bits_data(ifpu_io_out_bits_data),
    .io_out_bits_exc(ifpu_io_out_bits_exc),
    .io_covSum(ifpu_io_covSum),
    .metaAssert(ifpu_metaAssert),
    .metaReset(ifpu_metaReset)
  );
  FPToFP fpmu ( // @[FPU.scala 863:20]
    .clock(fpmu_clock),
    .reset(fpmu_reset),
    .io_in_valid(fpmu_io_in_valid),
    .io_in_bits_ren2(fpmu_io_in_bits_ren2),
    .io_in_bits_typeTagOut(fpmu_io_in_bits_typeTagOut),
    .io_in_bits_wflags(fpmu_io_in_bits_wflags),
    .io_in_bits_rm(fpmu_io_in_bits_rm),
    .io_in_bits_in1(fpmu_io_in_bits_in1),
    .io_in_bits_in2(fpmu_io_in_bits_in2),
    .io_out_bits_data(fpmu_io_out_bits_data),
    .io_out_bits_exc(fpmu_io_out_bits_exc),
    .io_lt(fpmu_io_lt),
    .io_covSum(fpmu_io_covSum),
    .metaAssert(fpmu_metaAssert),
    .metaReset(fpmu_metaReset)
  );
  FPUFMAPipe_1 dfma ( // @[FPU.scala 882:28]
    .clock(dfma_clock),
    .reset(dfma_reset),
    .io_in_valid(dfma_io_in_valid),
    .io_in_bits_ren3(dfma_io_in_bits_ren3),
    .io_in_bits_swap23(dfma_io_in_bits_swap23),
    .io_in_bits_rm(dfma_io_in_bits_rm),
    .io_in_bits_fmaCmd(dfma_io_in_bits_fmaCmd),
    .io_in_bits_in1(dfma_io_in_bits_in1),
    .io_in_bits_in2(dfma_io_in_bits_in2),
    .io_in_bits_in3(dfma_io_in_bits_in3),
    .io_out_bits_data(dfma_io_out_bits_data),
    .io_out_bits_exc(dfma_io_out_bits_exc),
    .io_covSum(dfma_io_covSum),
    .metaAssert(dfma_metaAssert),
    .metaReset(dfma_metaReset),
    .fma_halt(dfma_fma_halt)
  );
  DivSqrtRecFN_small divSqrt ( // @[FPU.scala 986:55]
    .clock(divSqrt_clock),
    .reset(divSqrt_reset),
    .io_inReady(divSqrt_io_inReady),
    .io_inValid(divSqrt_io_inValid),
    .io_sqrtOp(divSqrt_io_sqrtOp),
    .io_a(divSqrt_io_a),
    .io_b(divSqrt_io_b),
    .io_roundingMode(divSqrt_io_roundingMode),
    .io_outValid_div(divSqrt_io_outValid_div),
    .io_outValid_sqrt(divSqrt_io_outValid_sqrt),
    .io_out(divSqrt_io_out),
    .io_exceptionFlags(divSqrt_io_exceptionFlags),
    .io_covSum(divSqrt_io_covSum),
    .metaAssert(divSqrt_metaAssert),
    .metaReset(divSqrt_metaReset),
    .divSqrtRecFNToRaw_halt(divSqrt_divSqrtRecFNToRaw_halt)
  );
  DivSqrtRecFN_small_1 divSqrt_1 ( // @[FPU.scala 986:55]
    .clock(divSqrt_1_clock),
    .reset(divSqrt_1_reset),
    .io_inReady(divSqrt_1_io_inReady),
    .io_inValid(divSqrt_1_io_inValid),
    .io_sqrtOp(divSqrt_1_io_sqrtOp),
    .io_a(divSqrt_1_io_a),
    .io_b(divSqrt_1_io_b),
    .io_roundingMode(divSqrt_1_io_roundingMode),
    .io_outValid_div(divSqrt_1_io_outValid_div),
    .io_outValid_sqrt(divSqrt_1_io_outValid_sqrt),
    .io_out(divSqrt_1_io_out),
    .io_exceptionFlags(divSqrt_1_io_exceptionFlags),
    .io_covSum(divSqrt_1_io_covSum),
    .metaAssert(divSqrt_1_metaAssert),
    .metaReset(divSqrt_1_metaReset),
    .divSqrtRecFNToRaw_halt(divSqrt_1_divSqrtRecFNToRaw_halt)
  );
  assign regfile_ex_rs_0_addr = ex_ra_0;
  assign regfile_ex_rs_0_data = regfile[regfile_ex_rs_0_addr]; // @[FPU.scala 796:20]
  assign regfile_ex_rs_1_addr = ex_ra_1;
  assign regfile_ex_rs_1_data = regfile[regfile_ex_rs_1_addr]; // @[FPU.scala 796:20]
  assign regfile_ex_rs_2_addr = ex_ra_2;
  assign regfile_ex_rs_2_data = regfile[regfile_ex_rs_2_addr]; // @[FPU.scala 796:20]
  assign regfile_MPORT_data = _wdata_T_12 ? wdata_swizzledNaN : _wdata_T_6;
  assign regfile_MPORT_addr = load_wb_tag;
  assign regfile_MPORT_mask = 1'h1;
  assign regfile_MPORT_en = load_wb;
  assign regfile_MPORT_1_data = wtypeTag ? _wdata_T_19 : wdata_opts_bigger;
  assign regfile_MPORT_1_addr = divSqrt_wen ? divSqrt_waddr : wbInfo_0_rd;
  assign regfile_MPORT_1_mask = 1'h1;
  assign regfile_MPORT_1_en = wen[0] | divSqrt_wen;
  assign _load_wb_typeTag_T_2 = io_dmem_resp_type[1:0] - 2'h2; // @[FPU.scala 753:58]
  assign killm = io_killm | io_nack_mem; // @[FPU.scala 764:25]
  assign _killx_T = mem_reg_valid & killm; // @[FPU.scala 768:41]
  assign killx = io_killx | _killx_T; // @[FPU.scala 768:24]
  assign _mem_reg_valid_T_1 = ex_reg_valid & ~killx; // @[FPU.scala 769:33]
  assign wb_reg_valid_x7 = mem_reg_valid & ~killm; // @[FPU.scala 771:45]
  assign wdata_truncIdx = load_wb_typeTag[0]; // @[package.scala 31:49]
  assign _wdata_T_1 = wdata_truncIdx ? 64'h0 : 64'hffffffff00000000; // @[package.scala 32:76]
  assign _wdata_T_2 = _wdata_T_1 | load_wb_data; // @[FPU.scala 426:23]
  assign wdata_rawIn_sign = _wdata_T_2[63]; // @[rawFloatFromFN.scala 46:22]
  assign wdata_rawIn_expIn = _wdata_T_2[62:52]; // @[rawFloatFromFN.scala 47:23]
  assign wdata_rawIn_fractIn = _wdata_T_2[51:0]; // @[rawFloatFromFN.scala 48:25]
  assign wdata_rawIn_isZeroExpIn = wdata_rawIn_expIn == 11'h0; // @[rawFloatFromFN.scala 50:34]
  assign wdata_rawIn_isZeroFractIn = wdata_rawIn_fractIn == 52'h0; // @[rawFloatFromFN.scala 51:38]
  assign _wdata_rawIn_normDist_T_52 = wdata_rawIn_fractIn[1] ? 6'h32 : 6'h33; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_53 = wdata_rawIn_fractIn[2] ? 6'h31 : _wdata_rawIn_normDist_T_52; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_54 = wdata_rawIn_fractIn[3] ? 6'h30 : _wdata_rawIn_normDist_T_53; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_55 = wdata_rawIn_fractIn[4] ? 6'h2f : _wdata_rawIn_normDist_T_54; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_56 = wdata_rawIn_fractIn[5] ? 6'h2e : _wdata_rawIn_normDist_T_55; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_57 = wdata_rawIn_fractIn[6] ? 6'h2d : _wdata_rawIn_normDist_T_56; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_58 = wdata_rawIn_fractIn[7] ? 6'h2c : _wdata_rawIn_normDist_T_57; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_59 = wdata_rawIn_fractIn[8] ? 6'h2b : _wdata_rawIn_normDist_T_58; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_60 = wdata_rawIn_fractIn[9] ? 6'h2a : _wdata_rawIn_normDist_T_59; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_61 = wdata_rawIn_fractIn[10] ? 6'h29 : _wdata_rawIn_normDist_T_60; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_62 = wdata_rawIn_fractIn[11] ? 6'h28 : _wdata_rawIn_normDist_T_61; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_63 = wdata_rawIn_fractIn[12] ? 6'h27 : _wdata_rawIn_normDist_T_62; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_64 = wdata_rawIn_fractIn[13] ? 6'h26 : _wdata_rawIn_normDist_T_63; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_65 = wdata_rawIn_fractIn[14] ? 6'h25 : _wdata_rawIn_normDist_T_64; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_66 = wdata_rawIn_fractIn[15] ? 6'h24 : _wdata_rawIn_normDist_T_65; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_67 = wdata_rawIn_fractIn[16] ? 6'h23 : _wdata_rawIn_normDist_T_66; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_68 = wdata_rawIn_fractIn[17] ? 6'h22 : _wdata_rawIn_normDist_T_67; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_69 = wdata_rawIn_fractIn[18] ? 6'h21 : _wdata_rawIn_normDist_T_68; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_70 = wdata_rawIn_fractIn[19] ? 6'h20 : _wdata_rawIn_normDist_T_69; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_71 = wdata_rawIn_fractIn[20] ? 6'h1f : _wdata_rawIn_normDist_T_70; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_72 = wdata_rawIn_fractIn[21] ? 6'h1e : _wdata_rawIn_normDist_T_71; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_73 = wdata_rawIn_fractIn[22] ? 6'h1d : _wdata_rawIn_normDist_T_72; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_74 = wdata_rawIn_fractIn[23] ? 6'h1c : _wdata_rawIn_normDist_T_73; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_75 = wdata_rawIn_fractIn[24] ? 6'h1b : _wdata_rawIn_normDist_T_74; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_76 = wdata_rawIn_fractIn[25] ? 6'h1a : _wdata_rawIn_normDist_T_75; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_77 = wdata_rawIn_fractIn[26] ? 6'h19 : _wdata_rawIn_normDist_T_76; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_78 = wdata_rawIn_fractIn[27] ? 6'h18 : _wdata_rawIn_normDist_T_77; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_79 = wdata_rawIn_fractIn[28] ? 6'h17 : _wdata_rawIn_normDist_T_78; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_80 = wdata_rawIn_fractIn[29] ? 6'h16 : _wdata_rawIn_normDist_T_79; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_81 = wdata_rawIn_fractIn[30] ? 6'h15 : _wdata_rawIn_normDist_T_80; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_82 = wdata_rawIn_fractIn[31] ? 6'h14 : _wdata_rawIn_normDist_T_81; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_83 = wdata_rawIn_fractIn[32] ? 6'h13 : _wdata_rawIn_normDist_T_82; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_84 = wdata_rawIn_fractIn[33] ? 6'h12 : _wdata_rawIn_normDist_T_83; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_85 = wdata_rawIn_fractIn[34] ? 6'h11 : _wdata_rawIn_normDist_T_84; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_86 = wdata_rawIn_fractIn[35] ? 6'h10 : _wdata_rawIn_normDist_T_85; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_87 = wdata_rawIn_fractIn[36] ? 6'hf : _wdata_rawIn_normDist_T_86; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_88 = wdata_rawIn_fractIn[37] ? 6'he : _wdata_rawIn_normDist_T_87; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_89 = wdata_rawIn_fractIn[38] ? 6'hd : _wdata_rawIn_normDist_T_88; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_90 = wdata_rawIn_fractIn[39] ? 6'hc : _wdata_rawIn_normDist_T_89; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_91 = wdata_rawIn_fractIn[40] ? 6'hb : _wdata_rawIn_normDist_T_90; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_92 = wdata_rawIn_fractIn[41] ? 6'ha : _wdata_rawIn_normDist_T_91; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_93 = wdata_rawIn_fractIn[42] ? 6'h9 : _wdata_rawIn_normDist_T_92; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_94 = wdata_rawIn_fractIn[43] ? 6'h8 : _wdata_rawIn_normDist_T_93; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_95 = wdata_rawIn_fractIn[44] ? 6'h7 : _wdata_rawIn_normDist_T_94; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_96 = wdata_rawIn_fractIn[45] ? 6'h6 : _wdata_rawIn_normDist_T_95; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_97 = wdata_rawIn_fractIn[46] ? 6'h5 : _wdata_rawIn_normDist_T_96; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_98 = wdata_rawIn_fractIn[47] ? 6'h4 : _wdata_rawIn_normDist_T_97; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_99 = wdata_rawIn_fractIn[48] ? 6'h3 : _wdata_rawIn_normDist_T_98; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_100 = wdata_rawIn_fractIn[49] ? 6'h2 : _wdata_rawIn_normDist_T_99; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_101 = wdata_rawIn_fractIn[50] ? 6'h1 : _wdata_rawIn_normDist_T_100; // @[Mux.scala 47:69]
  assign wdata_rawIn_normDist = wdata_rawIn_fractIn[51] ? 6'h0 : _wdata_rawIn_normDist_T_101; // @[Mux.scala 47:69]
  assign _GEN_168 = {{63'd0}, wdata_rawIn_fractIn}; // @[rawFloatFromFN.scala 54:36]
  assign _wdata_rawIn_subnormFract_T = _GEN_168 << wdata_rawIn_normDist; // @[rawFloatFromFN.scala 54:36]
  assign wdata_rawIn_subnormFract = {_wdata_rawIn_subnormFract_T[50:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  assign _GEN_169 = {{6'd0}, wdata_rawIn_normDist}; // @[rawFloatFromFN.scala 57:26]
  assign _wdata_rawIn_adjustedExp_T = _GEN_169 ^ 12'hfff; // @[rawFloatFromFN.scala 57:26]
  assign _wdata_rawIn_adjustedExp_T_1 = wdata_rawIn_isZeroExpIn ? _wdata_rawIn_adjustedExp_T : {{1'd0}, wdata_rawIn_expIn}; // @[rawFloatFromFN.scala 56:16]
  assign _wdata_rawIn_adjustedExp_T_2 = wdata_rawIn_isZeroExpIn ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  assign _GEN_170 = {{9'd0}, _wdata_rawIn_adjustedExp_T_2}; // @[rawFloatFromFN.scala 60:22]
  assign _wdata_rawIn_adjustedExp_T_3 = 11'h400 | _GEN_170; // @[rawFloatFromFN.scala 60:22]
  assign _GEN_171 = {{1'd0}, _wdata_rawIn_adjustedExp_T_3}; // @[rawFloatFromFN.scala 59:15]
  assign wdata_rawIn_adjustedExp = _wdata_rawIn_adjustedExp_T_1 + _GEN_171; // @[rawFloatFromFN.scala 59:15]
  assign wdata_rawIn_isZero = wdata_rawIn_isZeroExpIn & wdata_rawIn_isZeroFractIn; // @[rawFloatFromFN.scala 62:34]
  assign wdata_rawIn_isSpecial = wdata_rawIn_adjustedExp[11:10] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  assign wdata_rawIn__isNaN = wdata_rawIn_isSpecial & ~wdata_rawIn_isZeroFractIn; // @[rawFloatFromFN.scala 66:33]
  assign wdata_rawIn__sExp = {1'b0,$signed(wdata_rawIn_adjustedExp)}; // @[rawFloatFromFN.scala 70:48]
  assign wdata_rawIn_out_sig_hi_lo = ~wdata_rawIn_isZero; // @[rawFloatFromFN.scala 72:29]
  assign wdata_rawIn_out_sig_lo = wdata_rawIn_isZeroExpIn ? wdata_rawIn_subnormFract : wdata_rawIn_fractIn; // @[rawFloatFromFN.scala 72:42]
  assign wdata_rawIn__sig = {1'h0,wdata_rawIn_out_sig_hi_lo,wdata_rawIn_out_sig_lo}; // @[Cat.scala 30:58]
  assign _wdata_T_4 = wdata_rawIn_isZero ? 3'h0 : wdata_rawIn__sExp[11:9]; // @[recFNFromFN.scala 48:16]
  assign _GEN_172 = {{2'd0}, wdata_rawIn__isNaN}; // @[recFNFromFN.scala 48:79]
  assign wdata_hi_lo = _wdata_T_4 | _GEN_172; // @[recFNFromFN.scala 48:79]
  assign wdata_lo_hi = wdata_rawIn__sExp[8:0]; // @[recFNFromFN.scala 50:23]
  assign wdata_lo_lo = wdata_rawIn__sig[51:0]; // @[recFNFromFN.scala 51:22]
  assign _wdata_T_6 = {wdata_rawIn_sign,wdata_hi_lo,wdata_lo_hi,wdata_lo_lo}; // @[Cat.scala 30:58]
  assign wdata_rawIn_sign_1 = _wdata_T_2[31]; // @[rawFloatFromFN.scala 46:22]
  assign wdata_rawIn_expIn_1 = _wdata_T_2[30:23]; // @[rawFloatFromFN.scala 47:23]
  assign wdata_rawIn_fractIn_1 = _wdata_T_2[22:0]; // @[rawFloatFromFN.scala 48:25]
  assign wdata_rawIn_isZeroExpIn_1 = wdata_rawIn_expIn_1 == 8'h0; // @[rawFloatFromFN.scala 50:34]
  assign wdata_rawIn_isZeroFractIn_1 = wdata_rawIn_fractIn_1 == 23'h0; // @[rawFloatFromFN.scala 51:38]
  assign _wdata_rawIn_normDist_T_125 = wdata_rawIn_fractIn_1[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_126 = wdata_rawIn_fractIn_1[2] ? 5'h14 : _wdata_rawIn_normDist_T_125; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_127 = wdata_rawIn_fractIn_1[3] ? 5'h13 : _wdata_rawIn_normDist_T_126; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_128 = wdata_rawIn_fractIn_1[4] ? 5'h12 : _wdata_rawIn_normDist_T_127; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_129 = wdata_rawIn_fractIn_1[5] ? 5'h11 : _wdata_rawIn_normDist_T_128; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_130 = wdata_rawIn_fractIn_1[6] ? 5'h10 : _wdata_rawIn_normDist_T_129; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_131 = wdata_rawIn_fractIn_1[7] ? 5'hf : _wdata_rawIn_normDist_T_130; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_132 = wdata_rawIn_fractIn_1[8] ? 5'he : _wdata_rawIn_normDist_T_131; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_133 = wdata_rawIn_fractIn_1[9] ? 5'hd : _wdata_rawIn_normDist_T_132; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_134 = wdata_rawIn_fractIn_1[10] ? 5'hc : _wdata_rawIn_normDist_T_133; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_135 = wdata_rawIn_fractIn_1[11] ? 5'hb : _wdata_rawIn_normDist_T_134; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_136 = wdata_rawIn_fractIn_1[12] ? 5'ha : _wdata_rawIn_normDist_T_135; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_137 = wdata_rawIn_fractIn_1[13] ? 5'h9 : _wdata_rawIn_normDist_T_136; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_138 = wdata_rawIn_fractIn_1[14] ? 5'h8 : _wdata_rawIn_normDist_T_137; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_139 = wdata_rawIn_fractIn_1[15] ? 5'h7 : _wdata_rawIn_normDist_T_138; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_140 = wdata_rawIn_fractIn_1[16] ? 5'h6 : _wdata_rawIn_normDist_T_139; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_141 = wdata_rawIn_fractIn_1[17] ? 5'h5 : _wdata_rawIn_normDist_T_140; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_142 = wdata_rawIn_fractIn_1[18] ? 5'h4 : _wdata_rawIn_normDist_T_141; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_143 = wdata_rawIn_fractIn_1[19] ? 5'h3 : _wdata_rawIn_normDist_T_142; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_144 = wdata_rawIn_fractIn_1[20] ? 5'h2 : _wdata_rawIn_normDist_T_143; // @[Mux.scala 47:69]
  assign _wdata_rawIn_normDist_T_145 = wdata_rawIn_fractIn_1[21] ? 5'h1 : _wdata_rawIn_normDist_T_144; // @[Mux.scala 47:69]
  assign wdata_rawIn_normDist_1 = wdata_rawIn_fractIn_1[22] ? 5'h0 : _wdata_rawIn_normDist_T_145; // @[Mux.scala 47:69]
  assign _GEN_173 = {{31'd0}, wdata_rawIn_fractIn_1}; // @[rawFloatFromFN.scala 54:36]
  assign _wdata_rawIn_subnormFract_T_2 = _GEN_173 << wdata_rawIn_normDist_1; // @[rawFloatFromFN.scala 54:36]
  assign wdata_rawIn_subnormFract_1 = {_wdata_rawIn_subnormFract_T_2[21:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  assign _GEN_174 = {{4'd0}, wdata_rawIn_normDist_1}; // @[rawFloatFromFN.scala 57:26]
  assign _wdata_rawIn_adjustedExp_T_5 = _GEN_174 ^ 9'h1ff; // @[rawFloatFromFN.scala 57:26]
  assign _wdata_rawIn_adjustedExp_T_6 = wdata_rawIn_isZeroExpIn_1 ? _wdata_rawIn_adjustedExp_T_5 : {{1'd0}, wdata_rawIn_expIn_1}; // @[rawFloatFromFN.scala 56:16]
  assign _wdata_rawIn_adjustedExp_T_7 = wdata_rawIn_isZeroExpIn_1 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  assign _GEN_175 = {{6'd0}, _wdata_rawIn_adjustedExp_T_7}; // @[rawFloatFromFN.scala 60:22]
  assign _wdata_rawIn_adjustedExp_T_8 = 8'h80 | _GEN_175; // @[rawFloatFromFN.scala 60:22]
  assign _GEN_176 = {{1'd0}, _wdata_rawIn_adjustedExp_T_8}; // @[rawFloatFromFN.scala 59:15]
  assign wdata_rawIn_adjustedExp_1 = _wdata_rawIn_adjustedExp_T_6 + _GEN_176; // @[rawFloatFromFN.scala 59:15]
  assign wdata_rawIn_isZero_1 = wdata_rawIn_isZeroExpIn_1 & wdata_rawIn_isZeroFractIn_1; // @[rawFloatFromFN.scala 62:34]
  assign wdata_rawIn_isSpecial_1 = wdata_rawIn_adjustedExp_1[8:7] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  assign wdata_rawIn_1_isNaN = wdata_rawIn_isSpecial_1 & ~wdata_rawIn_isZeroFractIn_1; // @[rawFloatFromFN.scala 66:33]
  assign wdata_rawIn_1_sExp = {1'b0,$signed(wdata_rawIn_adjustedExp_1)}; // @[rawFloatFromFN.scala 70:48]
  assign wdata_rawIn_out_sig_hi_lo_1 = ~wdata_rawIn_isZero_1; // @[rawFloatFromFN.scala 72:29]
  assign wdata_rawIn_out_sig_lo_1 = wdata_rawIn_isZeroExpIn_1 ? wdata_rawIn_subnormFract_1 : wdata_rawIn_fractIn_1; // @[rawFloatFromFN.scala 72:42]
  assign wdata_rawIn_1_sig = {1'h0,wdata_rawIn_out_sig_hi_lo_1,wdata_rawIn_out_sig_lo_1}; // @[Cat.scala 30:58]
  assign _wdata_T_8 = wdata_rawIn_isZero_1 ? 3'h0 : wdata_rawIn_1_sExp[8:6]; // @[recFNFromFN.scala 48:16]
  assign _GEN_177 = {{2'd0}, wdata_rawIn_1_isNaN}; // @[recFNFromFN.scala 48:79]
  assign wdata_hi_lo_1 = _wdata_T_8 | _GEN_177; // @[recFNFromFN.scala 48:79]
  assign wdata_lo_hi_1 = wdata_rawIn_1_sExp[5:0]; // @[recFNFromFN.scala 50:23]
  assign wdata_lo_lo_1 = wdata_rawIn_1_sig[22:0]; // @[recFNFromFN.scala 51:22]
  assign _wdata_T_10 = {wdata_rawIn_sign_1,wdata_hi_lo_1,wdata_lo_hi_1,wdata_lo_lo_1}; // @[Cat.scala 30:58]
  assign wdata_swizzledNaN_hi_hi_hi = _wdata_T_6[64:61]; // @[FPU.scala 332:8]
  assign wdata_swizzledNaN_hi_hi_lo = &_wdata_T_6[51:32]; // @[FPU.scala 333:42]
  assign wdata_swizzledNaN_hi_lo_hi = _wdata_T_6[59:53]; // @[FPU.scala 334:8]
  assign wdata_swizzledNaN_hi_lo_lo = _wdata_T_10[31]; // @[FPU.scala 335:8]
  assign wdata_swizzledNaN_lo_hi_lo = _wdata_T_10[32]; // @[FPU.scala 337:8]
  assign wdata_swizzledNaN_lo_lo = _wdata_T_10[30:0]; // @[FPU.scala 338:8]
  assign wdata_swizzledNaN = {wdata_swizzledNaN_hi_hi_hi,wdata_swizzledNaN_hi_hi_lo,wdata_swizzledNaN_hi_lo_hi,wdata_swizzledNaN_hi_lo_lo,_wdata_T_6[51:32],wdata_swizzledNaN_lo_hi_lo,wdata_swizzledNaN_lo_lo}; // @[Cat.scala 30:58]
  assign _wdata_T_12 = &_wdata_T_6[63:61]; // @[FPU.scala 243:56]
  assign wdata = _wdata_T_12 ? wdata_swizzledNaN : _wdata_T_6; // @[FPU.scala 339:8]
  assign _curOK_T_1 = &wdata[63:61]; // @[FPU.scala 243:56]
  assign _curOK_T_5 = &wdata[51:32]; // @[FPU.scala 380:96]
  assign _curOK_T_6 = wdata[60] == _curOK_T_5; // @[FPU.scala 380:55]
  assign curOK = ~_curOK_T_1 | _curOK_T_6; // @[FPU.scala 380:31]
  assign _T_2 = curOK | reset; // @[FPU.scala 800:11]
  assign _GEN_178 = {{1'd0}, load_wb_tag}; // @[FPU.scala 802:57]
  assign _T_5 = _GEN_178 + 6'h20; // @[FPU.scala 802:57]
  assign _T_11 = ~fp_decoder_io_sigs_swap12 & ~fp_decoder_io_sigs_swap23; // @[FPU.scala 817:29]
  assign _ex_rm_T_1 = ex_reg_inst[14:12] == 3'h7; // @[FPU.scala 821:38]
  assign _sfma_io_in_valid_T = ex_reg_valid & ex_reg_ctrl_fma; // @[FPU.scala 845:33]
  assign _sfma_io_in_valid_T_1 = ex_reg_ctrl_typeTagOut == 2'h0; // @[FPU.scala 845:70]
  assign sfma_io_in_bits_req_in1_unswizzled_hi_hi = regfile_ex_rs_0_data[31]; // @[FPU.scala 352:14]
  assign sfma_io_in_bits_req_in1_unswizzled_hi_lo = regfile_ex_rs_0_data[52]; // @[FPU.scala 353:14]
  assign sfma_io_in_bits_req_in1_unswizzled_lo = regfile_ex_rs_0_data[30:0]; // @[FPU.scala 354:14]
  assign sfma_io_in_bits_req_in1_floats_0 = {sfma_io_in_bits_req_in1_unswizzled_hi_hi,sfma_io_in_bits_req_in1_unswizzled_hi_lo,sfma_io_in_bits_req_in1_unswizzled_lo}; // @[Cat.scala 30:58]
  assign sfma_io_in_bits_req_in1_isbox = &regfile_ex_rs_0_data[64:60]; // @[FPU.scala 327:84]
  assign _sfma_io_in_bits_req_in1_T = sfma_io_in_bits_req_in1_isbox ? 33'h0 : 33'he0400000; // @[FPU.scala 367:31]
  assign _sfma_io_in_bits_req_in1_T_1 = sfma_io_in_bits_req_in1_floats_0 | _sfma_io_in_bits_req_in1_T; // @[FPU.scala 367:26]
  assign sfma_io_in_bits_req_in2_unswizzled_hi_hi = regfile_ex_rs_1_data[31]; // @[FPU.scala 352:14]
  assign sfma_io_in_bits_req_in2_unswizzled_hi_lo = regfile_ex_rs_1_data[52]; // @[FPU.scala 353:14]
  assign sfma_io_in_bits_req_in2_unswizzled_lo = regfile_ex_rs_1_data[30:0]; // @[FPU.scala 354:14]
  assign sfma_io_in_bits_req_in2_floats_0 = {sfma_io_in_bits_req_in2_unswizzled_hi_hi,sfma_io_in_bits_req_in2_unswizzled_hi_lo,sfma_io_in_bits_req_in2_unswizzled_lo}; // @[Cat.scala 30:58]
  assign sfma_io_in_bits_req_in2_isbox = &regfile_ex_rs_1_data[64:60]; // @[FPU.scala 327:84]
  assign _sfma_io_in_bits_req_in2_T = sfma_io_in_bits_req_in2_isbox ? 33'h0 : 33'he0400000; // @[FPU.scala 367:31]
  assign _sfma_io_in_bits_req_in2_T_1 = sfma_io_in_bits_req_in2_floats_0 | _sfma_io_in_bits_req_in2_T; // @[FPU.scala 367:26]
  assign sfma_io_in_bits_req_in3_unswizzled_hi_hi = regfile_ex_rs_2_data[31]; // @[FPU.scala 352:14]
  assign sfma_io_in_bits_req_in3_unswizzled_hi_lo = regfile_ex_rs_2_data[52]; // @[FPU.scala 353:14]
  assign sfma_io_in_bits_req_in3_unswizzled_lo = regfile_ex_rs_2_data[30:0]; // @[FPU.scala 354:14]
  assign sfma_io_in_bits_req_in3_floats_0 = {sfma_io_in_bits_req_in3_unswizzled_hi_hi,sfma_io_in_bits_req_in3_unswizzled_hi_lo,sfma_io_in_bits_req_in3_unswizzled_lo}; // @[Cat.scala 30:58]
  assign sfma_io_in_bits_req_in3_isbox = &regfile_ex_rs_2_data[64:60]; // @[FPU.scala 327:84]
  assign _sfma_io_in_bits_req_in3_T = sfma_io_in_bits_req_in3_isbox ? 33'h0 : 33'he0400000; // @[FPU.scala 367:31]
  assign _sfma_io_in_bits_req_in3_T_1 = sfma_io_in_bits_req_in3_floats_0 | _sfma_io_in_bits_req_in3_T; // @[FPU.scala 367:26]
  assign _sfma_io_in_bits_req_fmaCmd_T_3 = ~ex_reg_ctrl_ren3 & ex_reg_inst[27]; // @[FPU.scala 833:53]
  assign _GEN_179 = {{1'd0}, _sfma_io_in_bits_req_fmaCmd_T_3}; // @[FPU.scala 833:36]
  assign _fpiu_io_in_valid_T = ex_reg_ctrl_toint | ex_reg_ctrl_div; // @[FPU.scala 849:51]
  assign _fpiu_io_in_valid_T_1 = _fpiu_io_in_valid_T | ex_reg_ctrl_sqrt; // @[FPU.scala 849:66]
  assign _fpiu_io_in_valid_T_2 = ex_reg_ctrl_fastpipe & ex_reg_ctrl_wflags; // @[FPU.scala 849:103]
  assign _fpiu_io_in_valid_T_3 = _fpiu_io_in_valid_T_1 | _fpiu_io_in_valid_T_2; // @[FPU.scala 849:82]
  assign fpiu_io_in_bits_req_in1_hi_hi = sfma_io_in_bits_req_in1_floats_0[32]; // @[FPU.scala 268:17]
  assign fpiu_io_in_bits_req_in1_fractIn = sfma_io_in_bits_req_in1_floats_0[22:0]; // @[FPU.scala 269:20]
  assign fpiu_io_in_bits_req_in1_expIn = sfma_io_in_bits_req_in1_floats_0[31:23]; // @[FPU.scala 270:18]
  assign _fpiu_io_in_bits_req_in1_fractOut_T = {fpiu_io_in_bits_req_in1_fractIn, 53'h0}; // @[FPU.scala 271:28]
  assign fpiu_io_in_bits_req_in1_lo = _fpiu_io_in_bits_req_in1_fractOut_T[75:24]; // @[FPU.scala 271:38]
  assign fpiu_io_in_bits_req_in1_expOut_hi = fpiu_io_in_bits_req_in1_expIn[8:6]; // @[FPU.scala 273:26]
  assign _GEN_180 = {{3'd0}, fpiu_io_in_bits_req_in1_expIn}; // @[FPU.scala 274:31]
  assign _fpiu_io_in_bits_req_in1_expOut_commonCase_T_1 = _GEN_180 + 12'h800; // @[FPU.scala 274:31]
  assign fpiu_io_in_bits_req_in1_expOut_commonCase = _fpiu_io_in_bits_req_in1_expOut_commonCase_T_1 - 12'h100; // @[FPU.scala 274:48]
  assign _fpiu_io_in_bits_req_in1_expOut_T = fpiu_io_in_bits_req_in1_expOut_hi == 3'h0; // @[FPU.scala 275:19]
  assign _fpiu_io_in_bits_req_in1_expOut_T_1 = fpiu_io_in_bits_req_in1_expOut_hi >= 3'h6; // @[FPU.scala 275:36]
  assign _fpiu_io_in_bits_req_in1_expOut_T_2 = _fpiu_io_in_bits_req_in1_expOut_T | _fpiu_io_in_bits_req_in1_expOut_T_1; // @[FPU.scala 275:25]
  assign fpiu_io_in_bits_req_in1_expOut_lo = fpiu_io_in_bits_req_in1_expOut_commonCase[8:0]; // @[FPU.scala 275:65]
  assign _fpiu_io_in_bits_req_in1_expOut_T_3 = {fpiu_io_in_bits_req_in1_expOut_hi,fpiu_io_in_bits_req_in1_expOut_lo}; // @[Cat.scala 30:58]
  assign fpiu_io_in_bits_req_in1_hi_lo = _fpiu_io_in_bits_req_in1_expOut_T_2 ? _fpiu_io_in_bits_req_in1_expOut_T_3 : fpiu_io_in_bits_req_in1_expOut_commonCase; // @[FPU.scala 275:10]
  assign fpiu_io_in_bits_req_in1_floats_0 = {fpiu_io_in_bits_req_in1_hi_hi,fpiu_io_in_bits_req_in1_hi_lo,fpiu_io_in_bits_req_in1_lo}; // @[Cat.scala 30:58]
  assign fpiu_io_in_bits_req_in1_truncIdx = ex_reg_ctrl_typeTagIn[0]; // @[package.scala 31:49]
  assign _fpiu_io_in_bits_req_in1_T_1 = fpiu_io_in_bits_req_in1_truncIdx | sfma_io_in_bits_req_in1_isbox; // @[package.scala 32:76]
  assign _fpiu_io_in_bits_req_in1_T_3 = fpiu_io_in_bits_req_in1_truncIdx ? regfile_ex_rs_0_data : fpiu_io_in_bits_req_in1_floats_0; // @[package.scala 32:76]
  assign fpiu_io_in_bits_req_in2_hi_hi = sfma_io_in_bits_req_in2_floats_0[32]; // @[FPU.scala 268:17]
  assign fpiu_io_in_bits_req_in2_fractIn = sfma_io_in_bits_req_in2_floats_0[22:0]; // @[FPU.scala 269:20]
  assign fpiu_io_in_bits_req_in2_expIn = sfma_io_in_bits_req_in2_floats_0[31:23]; // @[FPU.scala 270:18]
  assign _fpiu_io_in_bits_req_in2_fractOut_T = {fpiu_io_in_bits_req_in2_fractIn, 53'h0}; // @[FPU.scala 271:28]
  assign fpiu_io_in_bits_req_in2_lo = _fpiu_io_in_bits_req_in2_fractOut_T[75:24]; // @[FPU.scala 271:38]
  assign fpiu_io_in_bits_req_in2_expOut_hi = fpiu_io_in_bits_req_in2_expIn[8:6]; // @[FPU.scala 273:26]
  assign _GEN_181 = {{3'd0}, fpiu_io_in_bits_req_in2_expIn}; // @[FPU.scala 274:31]
  assign _fpiu_io_in_bits_req_in2_expOut_commonCase_T_1 = _GEN_181 + 12'h800; // @[FPU.scala 274:31]
  assign fpiu_io_in_bits_req_in2_expOut_commonCase = _fpiu_io_in_bits_req_in2_expOut_commonCase_T_1 - 12'h100; // @[FPU.scala 274:48]
  assign _fpiu_io_in_bits_req_in2_expOut_T = fpiu_io_in_bits_req_in2_expOut_hi == 3'h0; // @[FPU.scala 275:19]
  assign _fpiu_io_in_bits_req_in2_expOut_T_1 = fpiu_io_in_bits_req_in2_expOut_hi >= 3'h6; // @[FPU.scala 275:36]
  assign _fpiu_io_in_bits_req_in2_expOut_T_2 = _fpiu_io_in_bits_req_in2_expOut_T | _fpiu_io_in_bits_req_in2_expOut_T_1; // @[FPU.scala 275:25]
  assign fpiu_io_in_bits_req_in2_expOut_lo = fpiu_io_in_bits_req_in2_expOut_commonCase[8:0]; // @[FPU.scala 275:65]
  assign _fpiu_io_in_bits_req_in2_expOut_T_3 = {fpiu_io_in_bits_req_in2_expOut_hi,fpiu_io_in_bits_req_in2_expOut_lo}; // @[Cat.scala 30:58]
  assign fpiu_io_in_bits_req_in2_hi_lo = _fpiu_io_in_bits_req_in2_expOut_T_2 ? _fpiu_io_in_bits_req_in2_expOut_T_3 : fpiu_io_in_bits_req_in2_expOut_commonCase; // @[FPU.scala 275:10]
  assign fpiu_io_in_bits_req_in2_floats_0 = {fpiu_io_in_bits_req_in2_hi_hi,fpiu_io_in_bits_req_in2_hi_lo,fpiu_io_in_bits_req_in2_lo}; // @[Cat.scala 30:58]
  assign _fpiu_io_in_bits_req_in2_T_1 = fpiu_io_in_bits_req_in1_truncIdx | sfma_io_in_bits_req_in2_isbox; // @[package.scala 32:76]
  assign _fpiu_io_in_bits_req_in2_T_3 = fpiu_io_in_bits_req_in1_truncIdx ? regfile_ex_rs_1_data : fpiu_io_in_bits_req_in2_floats_0; // @[package.scala 32:76]
  assign _ifpu_io_in_bits_in1_T = {{1'd0}, io_fromint_data}; // @[FPU.scala 861:29]
  assign _dfma_io_in_valid_T_1 = ex_reg_ctrl_typeTagOut == 2'h1; // @[FPU.scala 883:78]
  assign _memLatencyMask_T_2 = mem_ctrl_typeTagOut == 2'h0; // @[FPU.scala 880:72]
  assign _memLatencyMask_T_3 = mem_ctrl_fma & _memLatencyMask_T_2; // @[FPU.scala 880:56]
  assign _memLatencyMask_T_4 = _memLatencyMask_T_3 ? 2'h2 : 2'h0; // @[FPU.scala 895:23]
  assign _memLatencyMask_T_5 = mem_ctrl_typeTagOut == 2'h1; // @[FPU.scala 885:78]
  assign _memLatencyMask_T_6 = mem_ctrl_fma & _memLatencyMask_T_5; // @[FPU.scala 885:62]
  assign _memLatencyMask_T_7 = _memLatencyMask_T_6 ? 3'h4 : 3'h0; // @[FPU.scala 895:23]
  assign _memLatencyMask_T_8 = mem_ctrl_fastpipe | mem_ctrl_fromint; // @[FPU.scala 895:78]
  assign _GEN_188 = {{1'd0}, _memLatencyMask_T_8}; // @[FPU.scala 895:78]
  assign _memLatencyMask_T_9 = _GEN_188 | _memLatencyMask_T_4; // @[FPU.scala 895:78]
  assign _GEN_189 = {{1'd0}, _memLatencyMask_T_9}; // @[FPU.scala 895:78]
  assign memLatencyMask = _GEN_189 | _memLatencyMask_T_7; // @[FPU.scala 895:78]
  assign _mem_wen_T = mem_ctrl_fma | mem_ctrl_fastpipe; // @[FPU.scala 911:48]
  assign _mem_wen_T_1 = _mem_wen_T | mem_ctrl_fromint; // @[FPU.scala 911:69]
  assign mem_wen = mem_reg_valid & _mem_wen_T_1; // @[FPU.scala 911:31]
  assign _write_port_busy_T = ex_reg_ctrl_fastpipe ? 2'h2 : 2'h0; // @[FPU.scala 895:23]
  assign _write_port_busy_T_1 = ex_reg_ctrl_fromint ? 2'h2 : 2'h0; // @[FPU.scala 895:23]
  assign _write_port_busy_T_3 = ex_reg_ctrl_fma & _sfma_io_in_valid_T_1; // @[FPU.scala 880:56]
  assign _write_port_busy_T_4 = _write_port_busy_T_3 ? 3'h4 : 3'h0; // @[FPU.scala 895:23]
  assign _write_port_busy_T_6 = ex_reg_ctrl_fma & _dfma_io_in_valid_T_1; // @[FPU.scala 885:62]
  assign _write_port_busy_T_7 = _write_port_busy_T_6 ? 4'h8 : 4'h0; // @[FPU.scala 895:23]
  assign _write_port_busy_T_8 = _write_port_busy_T | _write_port_busy_T_1; // @[FPU.scala 895:78]
  assign _GEN_190 = {{1'd0}, _write_port_busy_T_8}; // @[FPU.scala 895:78]
  assign _write_port_busy_T_9 = _GEN_190 | _write_port_busy_T_4; // @[FPU.scala 895:78]
  assign _GEN_191 = {{1'd0}, _write_port_busy_T_9}; // @[FPU.scala 895:78]
  assign _write_port_busy_T_10 = _GEN_191 | _write_port_busy_T_7; // @[FPU.scala 895:78]
  assign _GEN_192 = {{1'd0}, memLatencyMask}; // @[FPU.scala 912:62]
  assign _write_port_busy_T_11 = _GEN_192 & _write_port_busy_T_10; // @[FPU.scala 912:62]
  assign _write_port_busy_T_12 = |_write_port_busy_T_11; // @[FPU.scala 912:89]
  assign _write_port_busy_T_13 = mem_wen & _write_port_busy_T_12; // @[FPU.scala 912:43]
  assign _write_port_busy_T_14 = ex_reg_ctrl_fastpipe ? 3'h4 : 3'h0; // @[FPU.scala 895:23]
  assign _write_port_busy_T_15 = ex_reg_ctrl_fromint ? 3'h4 : 3'h0; // @[FPU.scala 895:23]
  assign _write_port_busy_T_18 = _write_port_busy_T_3 ? 4'h8 : 4'h0; // @[FPU.scala 895:23]
  assign _write_port_busy_T_21 = _write_port_busy_T_6 ? 5'h10 : 5'h0; // @[FPU.scala 895:23]
  assign _write_port_busy_T_22 = _write_port_busy_T_14 | _write_port_busy_T_15; // @[FPU.scala 895:78]
  assign _GEN_193 = {{1'd0}, _write_port_busy_T_22}; // @[FPU.scala 895:78]
  assign _write_port_busy_T_23 = _GEN_193 | _write_port_busy_T_18; // @[FPU.scala 895:78]
  assign _GEN_194 = {{1'd0}, _write_port_busy_T_23}; // @[FPU.scala 895:78]
  assign _write_port_busy_T_24 = _GEN_194 | _write_port_busy_T_21; // @[FPU.scala 895:78]
  assign _GEN_195 = {{2'd0}, wen}; // @[FPU.scala 912:101]
  assign _write_port_busy_T_25 = _GEN_195 & _write_port_busy_T_24; // @[FPU.scala 912:101]
  assign _write_port_busy_T_26 = |_write_port_busy_T_25; // @[FPU.scala 912:128]
  assign _write_port_busy_T_27 = _write_port_busy_T_13 | _write_port_busy_T_26; // @[FPU.scala 912:93]
  assign _GEN_114 = wen[1] ? wbInfo_1_typeTag : wbInfo_0_typeTag; // @[FPU.scala 916:21]
  assign _GEN_118 = wen[2] ? wbInfo_2_typeTag : wbInfo_1_typeTag; // @[FPU.scala 916:21]
  assign _GEN_196 = {{1'd0}, wen[2:1]}; // @[FPU.scala 921:23]
  assign _wen_T_2 = _GEN_196 | memLatencyMask; // @[FPU.scala 921:23]
  assign _T_20 = ~write_port_busy & memLatencyMask[0]; // @[FPU.scala 924:30]
  assign _wbInfo_0_pipeid_T_7 = _memLatencyMask_T_6 ? 2'h3 : 2'h0; // @[FPU.scala 897:63]
  assign _GEN_197 = {{1'd0}, mem_ctrl_fromint}; // @[FPU.scala 897:108]
  assign _wbInfo_0_pipeid_T_9 = _GEN_197 | _memLatencyMask_T_4; // @[FPU.scala 897:108]
  assign _wbInfo_0_pipeid_T_10 = _wbInfo_0_pipeid_T_9 | _wbInfo_0_pipeid_T_7; // @[FPU.scala 897:108]
  assign _GEN_123 = _T_20 ? mem_ctrl_typeTagOut : {{1'd0}, _GEN_114}; // @[FPU.scala 924:52]
  assign _T_23 = ~write_port_busy & memLatencyMask[1]; // @[FPU.scala 924:30]
  assign _GEN_127 = _T_23 ? mem_ctrl_typeTagOut : {{1'd0}, _GEN_118}; // @[FPU.scala 924:52]
  assign _T_26 = ~write_port_busy & memLatencyMask[2]; // @[FPU.scala 924:30]
  assign _GEN_131 = _T_26 ? mem_ctrl_typeTagOut : {{1'd0}, wbInfo_2_typeTag}; // @[FPU.scala 924:52]
  assign _GEN_136 = mem_wen ? _GEN_123 : {{1'd0}, _GEN_114}; // @[FPU.scala 919:18]
  assign _GEN_140 = mem_wen ? _GEN_127 : {{1'd0}, _GEN_118}; // @[FPU.scala 919:18]
  assign _GEN_144 = mem_wen ? _GEN_131 : {{1'd0}, wbInfo_2_typeTag}; // @[FPU.scala 919:18]
  assign divSqrt_typeTag = divSqrt_1_io_outValid_div | divSqrt_1_io_outValid_sqrt; // @[FPU.scala 996:37]
  assign _T_52 = divSqrt_io_outValid_div | divSqrt_io_outValid_sqrt; // @[FPU.scala 996:37]
  assign _GEN_158 = _T_52 & ~divSqrt_killed; // @[FPU.scala 996:66]
  assign divSqrt_wen = divSqrt_typeTag ? ~divSqrt_killed : _GEN_158; // @[FPU.scala 996:66]
  assign waddr = divSqrt_wen ? divSqrt_waddr : wbInfo_0_rd; // @[FPU.scala 933:18]
  assign wtypeTag = divSqrt_wen ? divSqrt_typeTag : wbInfo_0_typeTag; // @[FPU.scala 934:21]
  assign _wdata_T_13 = wbInfo_0_pipeid == 2'h1; // @[package.scala 32:86]
  assign _wdata_T_14 = _wdata_T_13 ? ifpu_io_out_bits_data : fpmu_io_out_bits_data; // @[package.scala 32:76]
  assign _wdata_T_15 = wbInfo_0_pipeid == 2'h2; // @[package.scala 32:86]
  assign _wdata_T_16 = _wdata_T_15 ? sfma_io_out_bits_data : _wdata_T_14; // @[package.scala 32:76]
  assign _wdata_T_17 = wbInfo_0_pipeid == 2'h3; // @[package.scala 32:86]
  assign _wdata_T_18 = _wdata_T_17 ? dfma_io_out_bits_data : _wdata_T_16; // @[package.scala 32:76]
  assign _divSqrt_wdata_T_1 = &divSqrt_1_io_out[63:61]; // @[FPU.scala 243:56]
  assign divSqrt_wdata_maskedNaN = divSqrt_1_io_out & 65'h1efefffffffffffff; // @[FPU.scala 408:25]
  assign _divSqrt_wdata_T_2 = _divSqrt_wdata_T_1 ? divSqrt_wdata_maskedNaN : divSqrt_1_io_out; // @[FPU.scala 409:10]
  assign _GEN_159 = divSqrt_io_out; // @[FPU.scala 996:66]
  assign divSqrt_wdata = divSqrt_typeTag ? _divSqrt_wdata_T_2 : {{32'd0}, _GEN_159}; // @[FPU.scala 996:66]
  assign _wdata_T_19 = divSqrt_wen ? divSqrt_wdata : _wdata_T_18; // @[FPU.scala 935:22]
  assign wdata_opts_bigger_swizzledNaN_hi_hi_lo = &20'hfffff; // @[FPU.scala 333:42]
  assign wdata_opts_bigger_swizzledNaN_hi_lo_lo = _wdata_T_19[31]; // @[FPU.scala 335:8]
  assign wdata_opts_bigger_swizzledNaN_lo_hi_lo = _wdata_T_19[32]; // @[FPU.scala 337:8]
  assign wdata_opts_bigger_swizzledNaN_lo_lo = _wdata_T_19[30:0]; // @[FPU.scala 338:8]
  assign wdata_opts_bigger_swizzledNaN = {4'hf,wdata_opts_bigger_swizzledNaN_hi_hi_lo,7'h7f,wdata_opts_bigger_swizzledNaN_hi_lo_lo,20'hfffff,wdata_opts_bigger_swizzledNaN_lo_hi_lo,wdata_opts_bigger_swizzledNaN_lo_lo}; // @[Cat.scala 30:58]
  assign _wdata_opts_bigger_T = &3'h7; // @[FPU.scala 243:56]
  assign wdata_opts_bigger = _wdata_opts_bigger_T ? wdata_opts_bigger_swizzledNaN : 65'h1ffffffffffffffff; // @[FPU.scala 339:8]
  assign wdata_1 = wtypeTag ? _wdata_T_19 : wdata_opts_bigger; // @[package.scala 32:76]
  assign _wexc_T_1 = _wdata_T_13 ? ifpu_io_out_bits_exc : fpmu_io_out_bits_exc; // @[package.scala 32:76]
  assign _wexc_T_3 = _wdata_T_15 ? sfma_io_out_bits_exc : _wexc_T_1; // @[package.scala 32:76]
  assign wexc = _wdata_T_17 ? dfma_io_out_bits_exc : _wexc_T_3; // @[package.scala 32:76]
  assign frfWriteBundle_1_wrenf = wen[0] | divSqrt_wen; // @[FPU.scala 937:35]
  assign unswizzled_hi_hi_1 = wdata_1[31]; // @[FPU.scala 376:10]
  assign unswizzled_hi_lo_1 = wdata_1[52]; // @[FPU.scala 377:10]
  assign unswizzled_lo_1 = wdata_1[30:0]; // @[FPU.scala 378:10]
  assign unswizzled_1 = {unswizzled_hi_hi_1,unswizzled_hi_lo_1,unswizzled_lo_1}; // @[Cat.scala 30:58]
  assign _curOK_T_8 = &wdata_1[63:61]; // @[FPU.scala 243:56]
  assign _curOK_T_12 = &wdata_1[51:32]; // @[FPU.scala 380:96]
  assign _curOK_T_13 = wdata_1[60] == _curOK_T_12; // @[FPU.scala 380:55]
  assign curOK_1 = ~_curOK_T_8 | _curOK_T_13; // @[FPU.scala 380:31]
  assign _T_33 = curOK_1 | reset; // @[FPU.scala 938:11]
  assign _GEN_200 = {{1'd0}, waddr}; // @[FPU.scala 941:45]
  assign _T_36 = _GEN_200 + 6'h20; // @[FPU.scala 941:45]
  assign unrecoded_rawIn_exp = wdata_1[63:52]; // @[rawFloatFromRecFN.scala 50:21]
  assign unrecoded_rawIn_isZero = unrecoded_rawIn_exp[11:9] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign unrecoded_rawIn_isSpecial = unrecoded_rawIn_exp[11:10] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign unrecoded_rawIn__isNaN = unrecoded_rawIn_isSpecial & unrecoded_rawIn_exp[9]; // @[rawFloatFromRecFN.scala 55:33]
  assign unrecoded_rawIn__isInf = unrecoded_rawIn_isSpecial & ~unrecoded_rawIn_exp[9]; // @[rawFloatFromRecFN.scala 56:33]
  assign unrecoded_rawIn__sign = wdata_1[64]; // @[rawFloatFromRecFN.scala 58:25]
  assign unrecoded_rawIn__sExp = {1'b0,$signed(unrecoded_rawIn_exp)}; // @[rawFloatFromRecFN.scala 59:27]
  assign unrecoded_rawIn_out_sig_hi_lo = ~unrecoded_rawIn_isZero; // @[rawFloatFromRecFN.scala 60:39]
  assign unrecoded_rawIn_out_sig_lo = wdata_1[51:0]; // @[rawFloatFromRecFN.scala 60:51]
  assign unrecoded_rawIn__sig = {1'h0,unrecoded_rawIn_out_sig_hi_lo,unrecoded_rawIn_out_sig_lo}; // @[Cat.scala 30:58]
  assign unrecoded_isSubnormal = $signed(unrecoded_rawIn__sExp) < 13'sh402; // @[fNFromRecFN.scala 50:39]
  assign unrecoded_denormShiftDist = 6'h1 - unrecoded_rawIn__sExp[5:0]; // @[fNFromRecFN.scala 51:39]
  assign _unrecoded_denormFract_T_1 = unrecoded_rawIn__sig[53:1] >> unrecoded_denormShiftDist; // @[fNFromRecFN.scala 52:42]
  assign unrecoded_denormFract = _unrecoded_denormFract_T_1[51:0]; // @[fNFromRecFN.scala 52:60]
  assign _unrecoded_expOut_T_2 = unrecoded_rawIn__sExp[10:0] - 11'h401; // @[fNFromRecFN.scala 57:45]
  assign _unrecoded_expOut_T_3 = unrecoded_isSubnormal ? 11'h0 : _unrecoded_expOut_T_2; // @[fNFromRecFN.scala 55:16]
  assign _unrecoded_expOut_T_4 = unrecoded_rawIn__isNaN | unrecoded_rawIn__isInf; // @[fNFromRecFN.scala 59:44]
  assign _unrecoded_expOut_T_6 = _unrecoded_expOut_T_4 ? 11'h7ff : 11'h0; // @[Bitwise.scala 72:12]
  assign unrecoded_hi_lo = _unrecoded_expOut_T_3 | _unrecoded_expOut_T_6; // @[fNFromRecFN.scala 59:15]
  assign _unrecoded_fractOut_T_1 = unrecoded_rawIn__isInf ? 52'h0 : unrecoded_rawIn__sig[51:0]; // @[fNFromRecFN.scala 63:20]
  assign unrecoded_lo = unrecoded_isSubnormal ? unrecoded_denormFract : _unrecoded_fractOut_T_1; // @[fNFromRecFN.scala 61:16]
  assign unrecoded = {unrecoded_rawIn__sign,unrecoded_hi_lo,unrecoded_lo}; // @[Cat.scala 30:58]
  assign prevUnrecoded_rawIn_exp = unswizzled_1[31:23]; // @[rawFloatFromRecFN.scala 50:21]
  assign prevUnrecoded_rawIn_isZero = prevUnrecoded_rawIn_exp[8:6] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign prevUnrecoded_rawIn_isSpecial = prevUnrecoded_rawIn_exp[8:7] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign prevUnrecoded_rawIn__isNaN = prevUnrecoded_rawIn_isSpecial & prevUnrecoded_rawIn_exp[6]; // @[rawFloatFromRecFN.scala 55:33]
  assign prevUnrecoded_rawIn__isInf = prevUnrecoded_rawIn_isSpecial & ~prevUnrecoded_rawIn_exp[6]; // @[rawFloatFromRecFN.scala 56:33]
  assign prevUnrecoded_rawIn__sign = unswizzled_1[32]; // @[rawFloatFromRecFN.scala 58:25]
  assign prevUnrecoded_rawIn__sExp = {1'b0,$signed(prevUnrecoded_rawIn_exp)}; // @[rawFloatFromRecFN.scala 59:27]
  assign prevUnrecoded_rawIn_out_sig_hi_lo = ~prevUnrecoded_rawIn_isZero; // @[rawFloatFromRecFN.scala 60:39]
  assign prevUnrecoded_rawIn_out_sig_lo = unswizzled_1[22:0]; // @[rawFloatFromRecFN.scala 60:51]
  assign prevUnrecoded_rawIn__sig = {1'h0,prevUnrecoded_rawIn_out_sig_hi_lo,prevUnrecoded_rawIn_out_sig_lo}; // @[Cat.scala 30:58]
  assign prevUnrecoded_isSubnormal = $signed(prevUnrecoded_rawIn__sExp) < 10'sh82; // @[fNFromRecFN.scala 50:39]
  assign prevUnrecoded_denormShiftDist = 5'h1 - prevUnrecoded_rawIn__sExp[4:0]; // @[fNFromRecFN.scala 51:39]
  assign _prevUnrecoded_denormFract_T_1 = prevUnrecoded_rawIn__sig[24:1] >> prevUnrecoded_denormShiftDist; // @[fNFromRecFN.scala 52:42]
  assign prevUnrecoded_denormFract = _prevUnrecoded_denormFract_T_1[22:0]; // @[fNFromRecFN.scala 52:60]
  assign _prevUnrecoded_expOut_T_2 = prevUnrecoded_rawIn__sExp[7:0] - 8'h81; // @[fNFromRecFN.scala 57:45]
  assign _prevUnrecoded_expOut_T_3 = prevUnrecoded_isSubnormal ? 8'h0 : _prevUnrecoded_expOut_T_2; // @[fNFromRecFN.scala 55:16]
  assign _prevUnrecoded_expOut_T_4 = prevUnrecoded_rawIn__isNaN | prevUnrecoded_rawIn__isInf; // @[fNFromRecFN.scala 59:44]
  assign _prevUnrecoded_expOut_T_6 = _prevUnrecoded_expOut_T_4 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign prevUnrecoded_hi_lo = _prevUnrecoded_expOut_T_3 | _prevUnrecoded_expOut_T_6; // @[fNFromRecFN.scala 59:15]
  assign _prevUnrecoded_fractOut_T_1 = prevUnrecoded_rawIn__isInf ? 23'h0 : prevUnrecoded_rawIn__sig[22:0]; // @[fNFromRecFN.scala 63:20]
  assign prevUnrecoded_lo = prevUnrecoded_isSubnormal ? prevUnrecoded_denormFract : _prevUnrecoded_fractOut_T_1; // @[fNFromRecFN.scala 61:16]
  assign prevUnrecoded = {prevUnrecoded_rawIn__sign,prevUnrecoded_hi_lo,prevUnrecoded_lo}; // @[Cat.scala 30:58]
  assign hi = unrecoded[63:32]; // @[FPU.scala 441:21]
  assign lo = _curOK_T_8 ? prevUnrecoded : unrecoded[31:0]; // @[FPU.scala 441:44]
  assign _T_40 = {hi,lo}; // @[Cat.scala 30:58]
  assign wb_toint_valid = wb_reg_valid & wb_ctrl_toint; // @[FPU.scala 953:37]
  assign _io_fcsr_flags_valid_T = wb_toint_valid | divSqrt_wen; // @[FPU.scala 955:41]
  assign _io_fcsr_flags_bits_T = wb_toint_valid ? wb_toint_exc : 5'h0; // @[FPU.scala 957:8]
  assign _GEN_160 = divSqrt_io_exceptionFlags; // @[FPU.scala 996:66]
  assign divSqrt_flags = divSqrt_typeTag ? divSqrt_1_io_exceptionFlags : _GEN_160; // @[FPU.scala 996:66]
  assign _io_fcsr_flags_bits_T_1 = divSqrt_wen ? divSqrt_flags : 5'h0; // @[FPU.scala 958:8]
  assign _io_fcsr_flags_bits_T_2 = _io_fcsr_flags_bits_T | _io_fcsr_flags_bits_T_1; // @[FPU.scala 957:48]
  assign _io_fcsr_flags_bits_T_4 = wen[0] ? wexc : 5'h0; // @[FPU.scala 959:8]
  assign _divSqrt_write_port_busy_T = mem_ctrl_div | mem_ctrl_sqrt; // @[FPU.scala 961:47]
  assign _divSqrt_write_port_busy_T_1 = |wen; // @[FPU.scala 961:72]
  assign divSqrt_write_port_busy = _divSqrt_write_port_busy_T & _divSqrt_write_port_busy_T_1; // @[FPU.scala 961:65]
  assign _io_fcsr_rdy_T = ex_reg_valid & ex_reg_ctrl_wflags; // @[FPU.scala 962:33]
  assign _io_fcsr_rdy_T_1 = mem_reg_valid & mem_ctrl_wflags; // @[FPU.scala 962:68]
  assign _io_fcsr_rdy_T_2 = _io_fcsr_rdy_T | _io_fcsr_rdy_T_1; // @[FPU.scala 962:51]
  assign _io_fcsr_rdy_T_4 = _io_fcsr_rdy_T_2 | wb_toint_valid; // @[FPU.scala 962:87]
  assign _io_fcsr_rdy_T_6 = _io_fcsr_rdy_T_4 | _divSqrt_write_port_busy_T_1; // @[FPU.scala 962:120]
  assign _GEN_162 = ~divSqrt_1_io_inReady | ~divSqrt_io_inReady; // @[FPU.scala 994:34]
  assign divSqrt_inFlight = divSqrt_killed ? 1'h0 : _GEN_162; // @[FPU.scala 1004:27]
  assign _io_fcsr_rdy_T_7 = _io_fcsr_rdy_T_6 | divSqrt_inFlight; // @[FPU.scala 962:131]
  assign _io_nack_mem_T = write_port_busy | divSqrt_write_port_busy; // @[FPU.scala 963:34]
  assign _io_sboard_set_x27_T_3 = _memLatencyMask_T_6 | mem_ctrl_div; // @[FPU.scala 966:96]
  assign _io_sboard_clr_T_4 = wen[0] & _wdata_T_17; // @[FPU.scala 967:60]
  assign _io_illegal_rm_T_1 = io_inst[14:12] == 3'h5; // @[package.scala 15:47]
  assign _io_illegal_rm_T_2 = io_inst[14:12] == 3'h6; // @[package.scala 15:47]
  assign _io_illegal_rm_T_3 = _io_illegal_rm_T_1 | _io_illegal_rm_T_2; // @[package.scala 72:59]
  assign _io_illegal_rm_T_5 = io_inst[14:12] == 3'h7; // @[FPU.scala 971:67]
  assign _io_illegal_rm_T_6 = io_fcsr_rm >= 3'h5; // @[FPU.scala 971:87]
  assign _io_illegal_rm_T_7 = _io_illegal_rm_T_5 & _io_illegal_rm_T_6; // @[FPU.scala 971:73]
  assign _divSqrt_inValid_T_1 = mem_reg_valid & _divSqrt_write_port_busy_T; // @[FPU.scala 974:41]
  assign divSqrt_inValid = _divSqrt_inValid_T_1 & ~divSqrt_inFlight; // @[FPU.scala 974:76]
  assign _divSqrt_killed_T = divSqrt_inValid & killm; // @[FPU.scala 975:50]
  assign divSqrt_io_a_hi_hi = fpiu_io_out_bits_in_in1[64]; // @[FPU.scala 268:17]
  assign divSqrt_io_a_fractIn = fpiu_io_out_bits_in_in1[51:0]; // @[FPU.scala 269:20]
  assign divSqrt_io_a_expIn = fpiu_io_out_bits_in_in1[63:52]; // @[FPU.scala 270:18]
  assign _divSqrt_io_a_fractOut_T = {divSqrt_io_a_fractIn, 24'h0}; // @[FPU.scala 271:28]
  assign divSqrt_io_a_lo = _divSqrt_io_a_fractOut_T[75:53]; // @[FPU.scala 271:38]
  assign divSqrt_io_a_expOut_hi = divSqrt_io_a_expIn[11:9]; // @[FPU.scala 273:26]
  assign _divSqrt_io_a_expOut_commonCase_T_1 = divSqrt_io_a_expIn + 12'h100; // @[FPU.scala 274:31]
  assign divSqrt_io_a_expOut_commonCase = _divSqrt_io_a_expOut_commonCase_T_1 - 12'h800; // @[FPU.scala 274:48]
  assign _divSqrt_io_a_expOut_T = divSqrt_io_a_expOut_hi == 3'h0; // @[FPU.scala 275:19]
  assign _divSqrt_io_a_expOut_T_1 = divSqrt_io_a_expOut_hi >= 3'h6; // @[FPU.scala 275:36]
  assign _divSqrt_io_a_expOut_T_2 = _divSqrt_io_a_expOut_T | _divSqrt_io_a_expOut_T_1; // @[FPU.scala 275:25]
  assign divSqrt_io_a_expOut_lo = divSqrt_io_a_expOut_commonCase[5:0]; // @[FPU.scala 275:65]
  assign _divSqrt_io_a_expOut_T_3 = {divSqrt_io_a_expOut_hi,divSqrt_io_a_expOut_lo}; // @[Cat.scala 30:58]
  assign divSqrt_io_a_hi_lo = _divSqrt_io_a_expOut_T_2 ? _divSqrt_io_a_expOut_T_3 : divSqrt_io_a_expOut_commonCase[8:0]; // @[FPU.scala 275:10]
  assign divSqrt_io_a_hi = {divSqrt_io_a_hi_hi,divSqrt_io_a_hi_lo}; // @[Cat.scala 30:58]
  assign divSqrt_io_b_hi_hi = fpiu_io_out_bits_in_in2[64]; // @[FPU.scala 268:17]
  assign divSqrt_io_b_fractIn = fpiu_io_out_bits_in_in2[51:0]; // @[FPU.scala 269:20]
  assign divSqrt_io_b_expIn = fpiu_io_out_bits_in_in2[63:52]; // @[FPU.scala 270:18]
  assign _divSqrt_io_b_fractOut_T = {divSqrt_io_b_fractIn, 24'h0}; // @[FPU.scala 271:28]
  assign divSqrt_io_b_lo = _divSqrt_io_b_fractOut_T[75:53]; // @[FPU.scala 271:38]
  assign divSqrt_io_b_expOut_hi = divSqrt_io_b_expIn[11:9]; // @[FPU.scala 273:26]
  assign _divSqrt_io_b_expOut_commonCase_T_1 = divSqrt_io_b_expIn + 12'h100; // @[FPU.scala 274:31]
  assign divSqrt_io_b_expOut_commonCase = _divSqrt_io_b_expOut_commonCase_T_1 - 12'h800; // @[FPU.scala 274:48]
  assign _divSqrt_io_b_expOut_T = divSqrt_io_b_expOut_hi == 3'h0; // @[FPU.scala 275:19]
  assign _divSqrt_io_b_expOut_T_1 = divSqrt_io_b_expOut_hi >= 3'h6; // @[FPU.scala 275:36]
  assign _divSqrt_io_b_expOut_T_2 = _divSqrt_io_b_expOut_T | _divSqrt_io_b_expOut_T_1; // @[FPU.scala 275:25]
  assign divSqrt_io_b_expOut_lo = divSqrt_io_b_expOut_commonCase[5:0]; // @[FPU.scala 275:65]
  assign _divSqrt_io_b_expOut_T_3 = {divSqrt_io_b_expOut_hi,divSqrt_io_b_expOut_lo}; // @[Cat.scala 30:58]
  assign divSqrt_io_b_hi_lo = _divSqrt_io_b_expOut_T_2 ? _divSqrt_io_b_expOut_T_3 : divSqrt_io_b_expOut_commonCase[8:0]; // @[FPU.scala 275:10]
  assign divSqrt_io_b_hi = {divSqrt_io_b_hi_hi,divSqrt_io_b_hi_lo}; // @[Cat.scala 30:58]
  assign io_fcsr_flags_valid = _io_fcsr_flags_valid_T | wen[0]; // @[FPU.scala 955:23]
  assign io_fcsr_flags_bits = _io_fcsr_flags_bits_T_2 | _io_fcsr_flags_bits_T_4; // @[FPU.scala 956:22]
  assign io_store_data = fpiu_io_out_bits_store; // @[FPU.scala 851:17]
  assign io_toint_data = fpiu_io_out_bits_toint; // @[FPU.scala 852:17]
  assign io_fcsr_rdy = ~_io_fcsr_rdy_T_7; // @[FPU.scala 962:15]
  assign io_nack_mem = _io_nack_mem_T | divSqrt_inFlight; // @[FPU.scala 963:15]
  assign io_illegal_rm = _io_illegal_rm_T_3 | _io_illegal_rm_T_7; // @[FPU.scala 971:17]
  assign io_dec_wen = fp_decoder_io_sigs_wen; // @[FPU.scala 964:10]
  assign io_dec_ren1 = fp_decoder_io_sigs_ren1; // @[FPU.scala 964:10]
  assign io_dec_ren2 = fp_decoder_io_sigs_ren2; // @[FPU.scala 964:10]
  assign io_dec_ren3 = fp_decoder_io_sigs_ren3; // @[FPU.scala 964:10]
  assign io_sboard_set = wb_reg_valid & io_sboard_set_REG; // @[FPU.scala 966:17]
  assign io_sboard_clr = divSqrt_wen | _io_sboard_clr_T_4; // @[FPU.scala 967:17]
  assign io_sboard_clra = divSqrt_wen ? divSqrt_waddr : wbInfo_0_rd; // @[FPU.scala 968:18]
  assign fp_decoder_io_inst = io_inst; // @[FPU.scala 743:22]
  assign sfma_clock = clock;
  assign sfma_reset = reset;
  assign sfma_io_in_valid = _sfma_io_in_valid_T & _sfma_io_in_valid_T_1; // @[FPU.scala 845:20]
  assign sfma_io_in_bits_ren3 = ex_reg_ctrl_ren3; // @[FPU.scala 846:19]
  assign sfma_io_in_bits_swap23 = ex_reg_ctrl_swap23; // @[FPU.scala 846:19]
  assign sfma_io_in_bits_rm = _ex_rm_T_1 ? io_fcsr_rm : ex_reg_inst[14:12]; // @[FPU.scala 846:19]
  assign sfma_io_in_bits_fmaCmd = ex_reg_inst[3:2] | _GEN_179; // @[FPU.scala 846:19]
  assign sfma_io_in_bits_in1 = {{32'd0}, _sfma_io_in_bits_req_in1_T_1}; // @[FPU.scala 846:19]
  assign sfma_io_in_bits_in2 = {{32'd0}, _sfma_io_in_bits_req_in2_T_1}; // @[FPU.scala 846:19]
  assign sfma_io_in_bits_in3 = {{32'd0}, _sfma_io_in_bits_req_in3_T_1}; // @[FPU.scala 846:19]
  assign fpiu_clock = clock;
  assign fpiu_io_in_valid = ex_reg_valid & _fpiu_io_in_valid_T_3; // @[FPU.scala 849:20]
  assign fpiu_io_in_bits_ren2 = ex_reg_ctrl_ren2; // @[FPU.scala 850:19]
  assign fpiu_io_in_bits_typeTagIn = ex_reg_ctrl_typeTagIn; // @[FPU.scala 850:19]
  assign fpiu_io_in_bits_typeTagOut = ex_reg_ctrl_typeTagOut; // @[FPU.scala 850:19]
  assign fpiu_io_in_bits_wflags = ex_reg_ctrl_wflags; // @[FPU.scala 850:19]
  assign fpiu_io_in_bits_rm = _ex_rm_T_1 ? io_fcsr_rm : ex_reg_inst[14:12]; // @[FPU.scala 850:19]
  assign fpiu_io_in_bits_typ = ex_reg_inst[21:20]; // @[FPU.scala 850:19]
  assign fpiu_io_in_bits_fmt = ex_reg_inst[26:25]; // @[FPU.scala 850:19]
  assign fpiu_io_in_bits_in1 = _fpiu_io_in_bits_req_in1_T_1 ? _fpiu_io_in_bits_req_in1_T_3 : 65'he008000000000000; // @[FPU.scala 850:19]
  assign fpiu_io_in_bits_in2 = _fpiu_io_in_bits_req_in2_T_1 ? _fpiu_io_in_bits_req_in2_T_3 : 65'he008000000000000; // @[FPU.scala 850:19]
  assign ifpu_clock = clock;
  assign ifpu_reset = reset;
  assign ifpu_io_in_valid = ex_reg_valid & ex_reg_ctrl_fromint; // @[FPU.scala 859:20]
  assign ifpu_io_in_bits_typeTagIn = fpiu_io_in_bits_typeTagIn; // @[FPU.scala 860:19]
  assign ifpu_io_in_bits_wflags = fpiu_io_in_bits_wflags; // @[FPU.scala 860:19]
  assign ifpu_io_in_bits_rm = fpiu_io_in_bits_rm; // @[FPU.scala 860:19]
  assign ifpu_io_in_bits_typ = fpiu_io_in_bits_typ; // @[FPU.scala 860:19]
  assign ifpu_io_in_bits_in1 = _ifpu_io_in_bits_in1_T[63:0]; // @[FPU.scala 860:19 FPU.scala 861:23]
  assign fpmu_clock = clock;
  assign fpmu_reset = reset;
  assign fpmu_io_in_valid = ex_reg_valid & ex_reg_ctrl_fastpipe; // @[FPU.scala 864:20]
  assign fpmu_io_in_bits_ren2 = fpiu_io_in_bits_ren2; // @[FPU.scala 865:19]
  assign fpmu_io_in_bits_typeTagOut = fpiu_io_in_bits_typeTagOut; // @[FPU.scala 865:19]
  assign fpmu_io_in_bits_wflags = fpiu_io_in_bits_wflags; // @[FPU.scala 865:19]
  assign fpmu_io_in_bits_rm = fpiu_io_in_bits_rm; // @[FPU.scala 865:19]
  assign fpmu_io_in_bits_in1 = fpiu_io_in_bits_in1; // @[FPU.scala 865:19]
  assign fpmu_io_in_bits_in2 = fpiu_io_in_bits_in2; // @[FPU.scala 865:19]
  assign fpmu_io_lt = fpiu_io_out_bits_lt; // @[FPU.scala 866:14]
  assign dfma_clock = clock;
  assign dfma_reset = reset;
  assign dfma_io_in_valid = _sfma_io_in_valid_T & _dfma_io_in_valid_T_1; // @[FPU.scala 883:28]
  assign dfma_io_in_bits_ren3 = ex_reg_ctrl_ren3; // @[FPU.scala 884:27]
  assign dfma_io_in_bits_swap23 = ex_reg_ctrl_swap23; // @[FPU.scala 884:27]
  assign dfma_io_in_bits_rm = _ex_rm_T_1 ? io_fcsr_rm : ex_reg_inst[14:12]; // @[FPU.scala 884:27]
  assign dfma_io_in_bits_fmaCmd = ex_reg_inst[3:2] | _GEN_179; // @[FPU.scala 884:27]
  assign dfma_io_in_bits_in1 = regfile_ex_rs_0_data; // @[FPU.scala 884:27]
  assign dfma_io_in_bits_in2 = regfile_ex_rs_1_data; // @[FPU.scala 884:27]
  assign dfma_io_in_bits_in3 = regfile_ex_rs_2_data; // @[FPU.scala 884:27]
  assign divSqrt_clock = clock;
  assign divSqrt_reset = divSqrt_killed;
  assign divSqrt_io_inValid = divSqrt_inValid & _memLatencyMask_T_2; // @[FPU.scala 987:26]
  assign divSqrt_io_sqrtOp = mem_ctrl_sqrt; // @[FPU.scala 988:25]
  assign divSqrt_io_a = {divSqrt_io_a_hi,divSqrt_io_a_lo}; // @[FPU.scala 989:20]
  assign divSqrt_io_b = {divSqrt_io_b_hi,divSqrt_io_b_lo}; // @[FPU.scala 990:20]
  assign divSqrt_io_roundingMode = fpiu_io_out_bits_in_rm; // @[FPU.scala 991:31]
  assign divSqrt_1_clock = clock;
  assign divSqrt_1_reset = divSqrt_killed;
  assign divSqrt_1_io_inValid = divSqrt_inValid & _memLatencyMask_T_5; // @[FPU.scala 987:26]
  assign divSqrt_1_io_sqrtOp = mem_ctrl_sqrt; // @[FPU.scala 988:25]
  assign divSqrt_1_io_a = fpiu_io_out_bits_in_in1; // @[FPU.scala 989:20]
  assign divSqrt_1_io_b = fpiu_io_out_bits_in_in2; // @[FPU.scala 990:20]
  assign divSqrt_1_io_roundingMode = fpiu_io_out_bits_in_rm; // @[FPU.scala 991:31]
  assign FPU_cov_read_addr = FPU_state;
  assign FPU_cov_read_data = FPU_cov[FPU_cov_read_addr]; // @[Coverage map for FPU]
  assign FPU_cov_write_data = 1'h1;
  assign FPU_cov_write_addr = FPU_state;
  assign FPU_cov_write_mask = 1'h1;
  assign FPU_cov_write_en = 1'h1;
  assign wbInfo_0_typeTag_shl = {wbInfo_0_typeTag, 16'h0};
  assign wbInfo_0_typeTag_pad = {3'h0,wbInfo_0_typeTag_shl};
  assign wb_reg_valid_shl = {wb_reg_valid, 2'h0};
  assign wb_reg_valid_pad = {17'h0,wb_reg_valid_shl};
  assign mem_ctrl_sqrt_shl = {mem_ctrl_sqrt, 7'h0};
  assign mem_ctrl_sqrt_pad = {12'h0,mem_ctrl_sqrt_shl};
  assign divSqrt_killed_shl = {divSqrt_killed, 19'h0};
  assign divSqrt_killed_pad = divSqrt_killed_shl;
  assign ex_reg_ctrl_typeTagIn_shl = {ex_reg_ctrl_typeTagIn, 7'h0};
  assign ex_reg_ctrl_typeTagIn_pad = {11'h0,ex_reg_ctrl_typeTagIn_shl};
  assign ex_reg_ctrl_fromint_shl = {ex_reg_ctrl_fromint, 2'h0};
  assign ex_reg_ctrl_fromint_pad = {17'h0,ex_reg_ctrl_fromint_shl};
  assign mem_ctrl_typeTagOut_shl = {mem_ctrl_typeTagOut, 7'h0};
  assign mem_ctrl_typeTagOut_pad = {11'h0,mem_ctrl_typeTagOut_shl};
  assign wen_shl = {wen, 5'h0};
  assign wen_pad = {12'h0,wen_shl};
  assign wb_ctrl_toint_shl = {wb_ctrl_toint, 11'h0};
  assign wb_ctrl_toint_pad = {8'h0,wb_ctrl_toint_shl};
  assign ex_reg_ctrl_fastpipe_shl = {ex_reg_ctrl_fastpipe, 18'h0};
  assign ex_reg_ctrl_fastpipe_pad = {1'h0,ex_reg_ctrl_fastpipe_shl};
  assign write_port_busy_shl = {write_port_busy, 14'h0};
  assign write_port_busy_pad = {5'h0,write_port_busy_shl};
  assign mem_ctrl_fastpipe_shl = {mem_ctrl_fastpipe, 5'h0};
  assign mem_ctrl_fastpipe_pad = {14'h0,mem_ctrl_fastpipe_shl};
  assign ex_reg_ctrl_typeTagOut_shl = {ex_reg_ctrl_typeTagOut, 13'h0};
  assign ex_reg_ctrl_typeTagOut_pad = {5'h0,ex_reg_ctrl_typeTagOut_shl};
  assign mem_reg_valid_shl = {mem_reg_valid, 17'h0};
  assign mem_reg_valid_pad = {2'h0,mem_reg_valid_shl};
  assign mem_ctrl_div_shl = {mem_ctrl_div, 13'h0};
  assign mem_ctrl_div_pad = {6'h0,mem_ctrl_div_shl};
  assign wbInfo_0_pipeid_shl = {wbInfo_0_pipeid, 10'h0};
  assign wbInfo_0_pipeid_pad = {8'h0,wbInfo_0_pipeid_shl};
  assign mem_ctrl_toint_shl = {mem_ctrl_toint, 1'h0};
  assign mem_ctrl_toint_pad = {18'h0,mem_ctrl_toint_shl};
  assign ex_reg_ctrl_fma_shl = {ex_reg_ctrl_fma, 4'h0};
  assign ex_reg_ctrl_fma_pad = {15'h0,ex_reg_ctrl_fma_shl};
  assign ex_reg_valid_shl = {ex_reg_valid, 3'h0};
  assign ex_reg_valid_pad = {16'h0,ex_reg_valid_shl};
  assign mem_ctrl_fromint_shl = {mem_ctrl_fromint, 10'h0};
  assign mem_ctrl_fromint_pad = {9'h0,mem_ctrl_fromint_shl};
  assign mem_ctrl_fma_shl = {mem_ctrl_fma, 2'h0};
  assign mem_ctrl_fma_pad = {17'h0,mem_ctrl_fma_shl};
  assign FPU_xor7 = wbInfo_0_typeTag_pad ^ wb_reg_valid_pad;
  assign FPU_xor18 = divSqrt_killed_pad ^ ex_reg_ctrl_typeTagIn_pad;
  assign FPU_xor8 = mem_ctrl_sqrt_pad ^ FPU_xor18;
  assign FPU_xor3 = FPU_xor7 ^ FPU_xor8;
  assign FPU_xor9 = ex_reg_ctrl_fromint_pad ^ mem_ctrl_typeTagOut_pad;
  assign FPU_xor22 = wb_ctrl_toint_pad ^ ex_reg_ctrl_fastpipe_pad;
  assign FPU_xor10 = wen_pad ^ FPU_xor22;
  assign FPU_xor4 = FPU_xor9 ^ FPU_xor10;
  assign FPU_xor1 = FPU_xor3 ^ FPU_xor4;
  assign FPU_xor11 = write_port_busy_pad ^ mem_ctrl_fastpipe_pad;
  assign FPU_xor26 = mem_reg_valid_pad ^ mem_ctrl_div_pad;
  assign FPU_xor12 = ex_reg_ctrl_typeTagOut_pad ^ FPU_xor26;
  assign FPU_xor5 = FPU_xor11 ^ FPU_xor12;
  assign FPU_xor28 = mem_ctrl_toint_pad ^ ex_reg_ctrl_fma_pad;
  assign FPU_xor13 = wbInfo_0_pipeid_pad ^ FPU_xor28;
  assign FPU_xor30 = mem_ctrl_fromint_pad ^ mem_ctrl_fma_pad;
  assign FPU_xor14 = ex_reg_valid_pad ^ FPU_xor30;
  assign FPU_xor6 = FPU_xor13 ^ FPU_xor14;
  assign FPU_xor2 = FPU_xor5 ^ FPU_xor6;
  assign FPU_xor0 = FPU_xor1 ^ FPU_xor2;
  assign fpiu_sum = FPU_covSum + fpiu_io_covSum;
  assign fp_decoder_sum = fpiu_sum + fp_decoder_io_covSum;
  assign ifpu_sum = fp_decoder_sum + ifpu_io_covSum;
  assign sfma_sum = ifpu_sum + sfma_io_covSum;
  assign fpmu_sum = sfma_sum + fpmu_io_covSum;
  assign divSqrt_1_sum = fpmu_sum + divSqrt_1_io_covSum;
  assign dfma_sum = divSqrt_1_sum + dfma_io_covSum;
  assign divSqrt_sum = dfma_sum + divSqrt_io_covSum;
  assign io_covSum = divSqrt_sum;
  assign stopEn0 = load_wb & ~_T_2;
  assign stopEn1 = frfWriteBundle_1_wrenf & ~_T_33;
  assign fpiu_metaAssert_wire = fpiu_metaAssert;
  assign divSqrt_metaAssert_wire = divSqrt_metaAssert;
  assign fp_decoder_metaAssert_wire = fp_decoder_metaAssert;
  assign dfma_metaAssert_wire = dfma_metaAssert;
  assign ifpu_metaAssert_wire = ifpu_metaAssert;
  assign divSqrt_1_metaAssert_wire = divSqrt_1_metaAssert;
  assign sfma_metaAssert_wire = sfma_metaAssert;
  assign fpmu_metaAssert_wire = fpmu_metaAssert;
  assign FPU_or3 = stopEn0 | stopEn1;
  assign FPU_or10 = divSqrt_metaAssert_wire | divSqrt_1_metaAssert_wire;
  assign FPU_or4 = fp_decoder_metaAssert_wire | FPU_or10;
  assign FPU_or1 = FPU_or3 | FPU_or4;
  assign FPU_or5 = fpiu_metaAssert_wire | dfma_metaAssert_wire;
  assign FPU_or14 = ifpu_metaAssert_wire | sfma_metaAssert_wire;
  assign FPU_or6 = fpmu_metaAssert_wire | FPU_or14;
  assign FPU_or2 = FPU_or5 | FPU_or6;
  assign FPU_or0 = FPU_or1 | FPU_or2;
  assign metaAssert = FPU_metaAssert;
  assign fpiu_metaReset = metaReset | fpiu_halt;
  assign ifpu_metaReset = metaReset | ifpu_halt;
  assign sfma_metaReset = metaReset | sfma_halt;
  assign fpmu_metaReset = metaReset | fpmu_halt;
  assign divSqrt_1_metaReset = metaReset | divSqrt_1_halt;
  assign dfma_metaReset = metaReset | dfma_halt;
  assign divSqrt_metaReset = metaReset | divSqrt_halt;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {3{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    regfile[initvar] = _RAND_0[64:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ex_reg_valid = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ex_reg_inst = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  ex_reg_ctrl_ren2 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  ex_reg_ctrl_ren3 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  ex_reg_ctrl_swap23 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  ex_reg_ctrl_typeTagIn = _RAND_6[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  ex_reg_ctrl_typeTagOut = _RAND_7[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  ex_reg_ctrl_fromint = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  ex_reg_ctrl_toint = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  ex_reg_ctrl_fastpipe = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  ex_reg_ctrl_fma = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  ex_reg_ctrl_div = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  ex_reg_ctrl_sqrt = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  ex_reg_ctrl_wflags = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  ex_ra_0 = _RAND_15[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  ex_ra_1 = _RAND_16[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  ex_ra_2 = _RAND_17[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  load_wb = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  load_wb_typeTag = _RAND_19[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {2{`RANDOM}};
  load_wb_data = _RAND_20[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  load_wb_tag = _RAND_21[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  mem_reg_valid = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  mem_reg_inst = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  wb_reg_valid = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  mem_ctrl_typeTagOut = _RAND_25[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  mem_ctrl_fromint = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  mem_ctrl_toint = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  mem_ctrl_fastpipe = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  mem_ctrl_fma = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  mem_ctrl_div = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  mem_ctrl_sqrt = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  mem_ctrl_wflags = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  wb_ctrl_toint = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  divSqrt_waddr = _RAND_34[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  wen = _RAND_35[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  wbInfo_0_rd = _RAND_36[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  wbInfo_0_typeTag = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  wbInfo_0_pipeid = _RAND_38[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  wbInfo_1_rd = _RAND_39[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  wbInfo_1_typeTag = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  wbInfo_1_pipeid = _RAND_41[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  wbInfo_2_rd = _RAND_42[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  wbInfo_2_typeTag = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  wbInfo_2_pipeid = _RAND_44[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  write_port_busy = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  divSqrt_killed = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  wb_toint_exc = _RAND_47[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  io_sboard_set_REG = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  FPU_state = _RAND_49[19:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1048576; initvar = initvar+1)
    FPU_cov[initvar] = _RAND_50[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  FPU_covSum = _RAND_51[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  FPU_metaAssert = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(regfile_MPORT_en & regfile_MPORT_mask) begin
      regfile[regfile_MPORT_addr] <= regfile_MPORT_data; // @[FPU.scala 796:20]
    end
    if(regfile_MPORT_1_en & regfile_MPORT_1_mask) begin
      regfile[regfile_MPORT_1_addr] <= regfile_MPORT_1_data; // @[FPU.scala 796:20]
    end
    if (metaReset) begin
      ex_reg_valid <= 1'h0;
    end else if (reset) begin
      ex_reg_valid <= 1'h0;
    end else begin
      ex_reg_valid <= io_valid;
    end
    if (metaReset) begin
      ex_reg_inst <= 32'h0;
    end else if (io_valid) begin
      ex_reg_inst <= io_inst;
    end
    if (metaReset) begin
      ex_reg_ctrl_ren2 <= 1'h0;
    end else if (io_valid) begin
      ex_reg_ctrl_ren2 <= fp_decoder_io_sigs_ren2;
    end
    if (metaReset) begin
      ex_reg_ctrl_ren3 <= 1'h0;
    end else if (io_valid) begin
      ex_reg_ctrl_ren3 <= fp_decoder_io_sigs_ren3;
    end
    if (metaReset) begin
      ex_reg_ctrl_swap23 <= 1'h0;
    end else if (io_valid) begin
      ex_reg_ctrl_swap23 <= fp_decoder_io_sigs_swap23;
    end
    if (metaReset) begin
      ex_reg_ctrl_typeTagIn <= 2'h0;
    end else if (io_valid) begin
      ex_reg_ctrl_typeTagIn <= fp_decoder_io_sigs_typeTagIn;
    end
    if (metaReset) begin
      ex_reg_ctrl_typeTagOut <= 2'h0;
    end else if (io_valid) begin
      ex_reg_ctrl_typeTagOut <= fp_decoder_io_sigs_typeTagOut;
    end
    if (metaReset) begin
      ex_reg_ctrl_fromint <= 1'h0;
    end else if (io_valid) begin
      ex_reg_ctrl_fromint <= fp_decoder_io_sigs_fromint;
    end
    if (metaReset) begin
      ex_reg_ctrl_toint <= 1'h0;
    end else if (io_valid) begin
      ex_reg_ctrl_toint <= fp_decoder_io_sigs_toint;
    end
    if (metaReset) begin
      ex_reg_ctrl_fastpipe <= 1'h0;
    end else if (io_valid) begin
      ex_reg_ctrl_fastpipe <= fp_decoder_io_sigs_fastpipe;
    end
    if (metaReset) begin
      ex_reg_ctrl_fma <= 1'h0;
    end else if (io_valid) begin
      ex_reg_ctrl_fma <= fp_decoder_io_sigs_fma;
    end
    if (metaReset) begin
      ex_reg_ctrl_div <= 1'h0;
    end else if (io_valid) begin
      ex_reg_ctrl_div <= fp_decoder_io_sigs_div;
    end
    if (metaReset) begin
      ex_reg_ctrl_sqrt <= 1'h0;
    end else if (io_valid) begin
      ex_reg_ctrl_sqrt <= fp_decoder_io_sigs_sqrt;
    end
    if (metaReset) begin
      ex_reg_ctrl_wflags <= 1'h0;
    end else if (io_valid) begin
      ex_reg_ctrl_wflags <= fp_decoder_io_sigs_wflags;
    end
    if (metaReset) begin
      ex_ra_0 <= 5'h0;
    end else if (io_valid) begin
      if (fp_decoder_io_sigs_ren2) begin
        if (fp_decoder_io_sigs_swap12) begin
          ex_ra_0 <= io_inst[24:20];
        end else if (fp_decoder_io_sigs_ren1) begin
          if (~fp_decoder_io_sigs_swap12) begin
            ex_ra_0 <= io_inst[19:15];
          end
        end
      end else if (fp_decoder_io_sigs_ren1) begin
        if (~fp_decoder_io_sigs_swap12) begin
          ex_ra_0 <= io_inst[19:15];
        end
      end
    end
    if (metaReset) begin
      ex_ra_1 <= 5'h0;
    end else if (io_valid) begin
      if (fp_decoder_io_sigs_ren2) begin
        if (_T_11) begin
          ex_ra_1 <= io_inst[24:20];
        end else if (fp_decoder_io_sigs_ren1) begin
          if (fp_decoder_io_sigs_swap12) begin
            ex_ra_1 <= io_inst[19:15];
          end
        end
      end else if (fp_decoder_io_sigs_ren1) begin
        if (fp_decoder_io_sigs_swap12) begin
          ex_ra_1 <= io_inst[19:15];
        end
      end
    end
    if (metaReset) begin
      ex_ra_2 <= 5'h0;
    end else if (io_valid) begin
      if (fp_decoder_io_sigs_ren3) begin
        ex_ra_2 <= io_inst[31:27];
      end else if (fp_decoder_io_sigs_ren2) begin
        if (fp_decoder_io_sigs_swap23) begin
          ex_ra_2 <= io_inst[24:20];
        end
      end
    end
    if (metaReset) begin
      load_wb <= 1'h0;
    end else begin
      load_wb <= io_dmem_resp_val;
    end
    if (metaReset) begin
      load_wb_typeTag <= 2'h0;
    end else if (io_dmem_resp_val) begin
      load_wb_typeTag <= _load_wb_typeTag_T_2;
    end
    if (metaReset) begin
      load_wb_data <= 64'h0;
    end else if (io_dmem_resp_val) begin
      load_wb_data <= io_dmem_resp_data;
    end
    if (metaReset) begin
      load_wb_tag <= 5'h0;
    end else if (io_dmem_resp_val) begin
      load_wb_tag <= io_dmem_resp_tag;
    end
    if (metaReset) begin
      mem_reg_valid <= 1'h0;
    end else if (reset) begin
      mem_reg_valid <= 1'h0;
    end else begin
      mem_reg_valid <= _mem_reg_valid_T_1;
    end
    if (metaReset) begin
      mem_reg_inst <= 32'h0;
    end else if (ex_reg_valid) begin
      mem_reg_inst <= ex_reg_inst;
    end
    if (metaReset) begin
      wb_reg_valid <= 1'h0;
    end else if (reset) begin
      wb_reg_valid <= 1'h0;
    end else begin
      wb_reg_valid <= wb_reg_valid_x7;
    end
    if (metaReset) begin
      mem_ctrl_typeTagOut <= 2'h0;
    end else if (ex_reg_valid) begin
      mem_ctrl_typeTagOut <= ex_reg_ctrl_typeTagOut;
    end
    if (metaReset) begin
      mem_ctrl_fromint <= 1'h0;
    end else if (ex_reg_valid) begin
      mem_ctrl_fromint <= ex_reg_ctrl_fromint;
    end
    if (metaReset) begin
      mem_ctrl_toint <= 1'h0;
    end else if (ex_reg_valid) begin
      mem_ctrl_toint <= ex_reg_ctrl_toint;
    end
    if (metaReset) begin
      mem_ctrl_fastpipe <= 1'h0;
    end else if (ex_reg_valid) begin
      mem_ctrl_fastpipe <= ex_reg_ctrl_fastpipe;
    end
    if (metaReset) begin
      mem_ctrl_fma <= 1'h0;
    end else if (ex_reg_valid) begin
      mem_ctrl_fma <= ex_reg_ctrl_fma;
    end
    if (metaReset) begin
      mem_ctrl_div <= 1'h0;
    end else if (ex_reg_valid) begin
      mem_ctrl_div <= ex_reg_ctrl_div;
    end
    if (metaReset) begin
      mem_ctrl_sqrt <= 1'h0;
    end else if (ex_reg_valid) begin
      mem_ctrl_sqrt <= ex_reg_ctrl_sqrt;
    end
    if (metaReset) begin
      mem_ctrl_wflags <= 1'h0;
    end else if (ex_reg_valid) begin
      mem_ctrl_wflags <= ex_reg_ctrl_wflags;
    end
    if (metaReset) begin
      wb_ctrl_toint <= 1'h0;
    end else if (mem_reg_valid) begin
      wb_ctrl_toint <= mem_ctrl_toint;
    end
    if (metaReset) begin
      divSqrt_waddr <= 5'h0;
    end else if (divSqrt_inValid) begin
      divSqrt_waddr <= mem_reg_inst[11:7];
    end
    if (metaReset) begin
      wen <= 3'h0;
    end else if (reset) begin
      wen <= 3'h0;
    end else if (mem_wen) begin
      if (~killm) begin
        wen <= _wen_T_2;
      end else begin
        wen <= {{1'd0}, wen[2:1]};
      end
    end else begin
      wen <= {{1'd0}, wen[2:1]};
    end
    if (metaReset) begin
      wbInfo_0_rd <= 5'h0;
    end else if (mem_wen) begin
      if (_T_20) begin
        wbInfo_0_rd <= mem_reg_inst[11:7];
      end else if (wen[1]) begin
        wbInfo_0_rd <= wbInfo_1_rd;
      end
    end else if (wen[1]) begin
      wbInfo_0_rd <= wbInfo_1_rd;
    end
    if (metaReset) begin
      wbInfo_0_typeTag <= 1'h0;
    end else begin
      wbInfo_0_typeTag <= _GEN_136[0];
    end
    if (metaReset) begin
      wbInfo_0_pipeid <= 2'h0;
    end else if (mem_wen) begin
      if (_T_20) begin
        wbInfo_0_pipeid <= _wbInfo_0_pipeid_T_10;
      end else if (wen[1]) begin
        wbInfo_0_pipeid <= wbInfo_1_pipeid;
      end
    end else if (wen[1]) begin
      wbInfo_0_pipeid <= wbInfo_1_pipeid;
    end
    if (metaReset) begin
      wbInfo_1_rd <= 5'h0;
    end else if (mem_wen) begin
      if (_T_23) begin
        wbInfo_1_rd <= mem_reg_inst[11:7];
      end else if (wen[2]) begin
        wbInfo_1_rd <= wbInfo_2_rd;
      end
    end else if (wen[2]) begin
      wbInfo_1_rd <= wbInfo_2_rd;
    end
    if (metaReset) begin
      wbInfo_1_typeTag <= 1'h0;
    end else begin
      wbInfo_1_typeTag <= _GEN_140[0];
    end
    if (metaReset) begin
      wbInfo_1_pipeid <= 2'h0;
    end else if (mem_wen) begin
      if (_T_23) begin
        wbInfo_1_pipeid <= _wbInfo_0_pipeid_T_10;
      end else if (wen[2]) begin
        wbInfo_1_pipeid <= wbInfo_2_pipeid;
      end
    end else if (wen[2]) begin
      wbInfo_1_pipeid <= wbInfo_2_pipeid;
    end
    if (metaReset) begin
      wbInfo_2_rd <= 5'h0;
    end else if (mem_wen) begin
      if (_T_26) begin
        wbInfo_2_rd <= mem_reg_inst[11:7];
      end
    end
    if (metaReset) begin
      wbInfo_2_typeTag <= 1'h0;
    end else begin
      wbInfo_2_typeTag <= _GEN_144[0];
    end
    if (metaReset) begin
      wbInfo_2_pipeid <= 2'h0;
    end else if (mem_wen) begin
      if (_T_26) begin
        wbInfo_2_pipeid <= _wbInfo_0_pipeid_T_10;
      end
    end
    if (metaReset) begin
      write_port_busy <= 1'h0;
    end else if (ex_reg_valid) begin
      write_port_busy <= _write_port_busy_T_27;
    end
    if (metaReset) begin
      divSqrt_killed <= 1'h0;
    end else begin
      divSqrt_killed <= reset | _divSqrt_killed_T;
    end
    if (metaReset) begin
      wb_toint_exc <= 5'h0;
    end else if (mem_ctrl_toint) begin
      wb_toint_exc <= fpiu_io_out_bits_exc;
    end
    if (metaReset) begin
      io_sboard_set_REG <= 1'h0;
    end else begin
      io_sboard_set_REG <= _io_sboard_set_x27_T_3 | mem_ctrl_sqrt;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (load_wb & ~_T_2) begin
          $fwrite(32'h80000002,"Assertion failed\n    at FPU.scala:800 assert(consistent(wdata))\n"); // @[FPU.scala 800:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (load_wb & ~_T_2) begin
          $fatal; // @[FPU.scala 800:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (load_wb & ~reset) begin
          //$fwrite(32'h80000002,"12487: %d %x",load_wb_tag,load_wb_data);
          $fwrite(32'h80000002,"f%d p%d 0x%x\n",load_wb_tag,_T_5,load_wb_data); // @[FPU.scala 802:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (frfWriteBundle_1_wrenf & ~_T_33) begin
          $fwrite(32'h80000002,"Assertion failed\n    at FPU.scala:938 assert(consistent(wdata))\n"); // @[FPU.scala 938:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (frfWriteBundle_1_wrenf & ~_T_33) begin
          $fatal; // @[FPU.scala 938:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (frfWriteBundle_1_wrenf & ~reset) begin
          //$fwrite(32'h80000002,"12521: %d %x",waddr,_T_40);
          $fwrite(32'h80000002,"f%d p%d 0x%x\n",waddr,_T_36,_T_40); // @[FPU.scala 941:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    FPU_state <= FPU_xor0;
    if (!(FPU_cov_read_data)) begin
      FPU_covSum <= FPU_covSum + 1'h1;
    end
    if (metaReset) begin
      FPU_metaAssert <= 1'h0;
    end else begin
      FPU_metaAssert <= FPU_metaAssert | FPU_or0;
    end
  end
  always @(posedge clock) begin
    if(FPU_cov_write_en & FPU_cov_write_mask) begin
      FPU_cov[FPU_cov_write_addr] <= FPU_cov_write_data; // @[Coverage map for FPU]
    end
  end
endmodule
module HellaCacheArbiter(
  input         clock,
  output        io_requestor_0_req_ready,
  input         io_requestor_0_req_valid,
  input  [39:0] io_requestor_0_req_bits_addr,
  input         io_requestor_0_s1_kill,
  output        io_requestor_0_s2_nack,
  output        io_requestor_0_resp_valid,
  output [63:0] io_requestor_0_resp_bits_data,
  output        io_requestor_0_s2_xcpt_ae_ld,
  output        io_requestor_1_req_ready,
  input         io_requestor_1_req_valid,
  input  [39:0] io_requestor_1_req_bits_addr,
  input  [6:0]  io_requestor_1_req_bits_tag,
  input  [4:0]  io_requestor_1_req_bits_cmd,
  input  [1:0]  io_requestor_1_req_bits_size,
  input         io_requestor_1_req_bits_signed,
  input         io_requestor_1_s1_kill,
  input  [63:0] io_requestor_1_s1_data_data,
  output        io_requestor_1_s2_nack,
  output        io_requestor_1_resp_valid,
  output [6:0]  io_requestor_1_resp_bits_tag,
  output [1:0]  io_requestor_1_resp_bits_size,
  output [63:0] io_requestor_1_resp_bits_data,
  output        io_requestor_1_resp_bits_replay,
  output        io_requestor_1_resp_bits_has_data,
  output [63:0] io_requestor_1_resp_bits_data_word_bypass,
  output        io_requestor_1_replay_next,
  output        io_requestor_1_s2_xcpt_ma_ld,
  output        io_requestor_1_s2_xcpt_ma_st,
  output        io_requestor_1_s2_xcpt_pf_ld,
  output        io_requestor_1_s2_xcpt_pf_st,
  output        io_requestor_1_s2_xcpt_ae_ld,
  output        io_requestor_1_s2_xcpt_ae_st,
  output        io_requestor_1_ordered,
  output        io_requestor_1_perf_release,
  output        io_requestor_1_perf_grant,
  input         io_mem_req_ready,
  output        io_mem_req_valid,
  output [39:0] io_mem_req_bits_addr,
  output [6:0]  io_mem_req_bits_tag,
  output [4:0]  io_mem_req_bits_cmd,
  output [1:0]  io_mem_req_bits_size,
  output        io_mem_req_bits_signed,
  output        io_mem_req_bits_phys,
  output        io_mem_s1_kill,
  output [63:0] io_mem_s1_data_data,
  input         io_mem_s2_nack,
  input         io_mem_resp_valid,
  input  [6:0]  io_mem_resp_bits_tag,
  input  [1:0]  io_mem_resp_bits_size,
  input  [63:0] io_mem_resp_bits_data,
  input         io_mem_resp_bits_replay,
  input         io_mem_resp_bits_has_data,
  input  [63:0] io_mem_resp_bits_data_word_bypass,
  input         io_mem_replay_next,
  input         io_mem_s2_xcpt_ma_ld,
  input         io_mem_s2_xcpt_ma_st,
  input         io_mem_s2_xcpt_pf_ld,
  input         io_mem_s2_xcpt_pf_st,
  input         io_mem_s2_xcpt_ae_ld,
  input         io_mem_s2_xcpt_ae_st,
  input         io_mem_ordered,
  input         io_mem_perf_release,
  input         io_mem_perf_grant,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  reg  s1_id; // @[HellaCacheArbiter.scala 19:20]
  reg [31:0] _RAND_0;
  reg  s2_id; // @[HellaCacheArbiter.scala 20:20]
  reg [31:0] _RAND_1;
  wire [7:0] _io_mem_req_bits_tag_T; // @[Cat.scala 30:58]
  wire [7:0] _GEN_1; // @[HellaCacheArbiter.scala 49:26]
  wire  tag_hit; // @[HellaCacheArbiter.scala 59:57]
  reg  HellaCacheArbiter_state; // @[Register tracking HellaCacheArbiter state]
  reg [31:0] _RAND_2;
  reg  HellaCacheArbiter_cov [0:1]; // @[Coverage map for HellaCacheArbiter]
  reg [31:0] _RAND_3;
  wire  HellaCacheArbiter_cov_read_data; // @[Coverage map for HellaCacheArbiter]
  wire  HellaCacheArbiter_cov_read_addr; // @[Coverage map for HellaCacheArbiter]
  wire  HellaCacheArbiter_cov_write_data; // @[Coverage map for HellaCacheArbiter]
  wire  HellaCacheArbiter_cov_write_addr; // @[Coverage map for HellaCacheArbiter]
  wire  HellaCacheArbiter_cov_write_mask; // @[Coverage map for HellaCacheArbiter]
  wire  HellaCacheArbiter_cov_write_en; // @[Coverage map for HellaCacheArbiter]
  reg [29:0] HellaCacheArbiter_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_4;
  wire  s1_id_shl;
  wire  s1_id_pad;
  assign _io_mem_req_bits_tag_T = {io_requestor_1_req_bits_tag,1'h1}; // @[Cat.scala 30:58]
  assign _GEN_1 = io_requestor_0_req_valid ? 8'h0 : _io_mem_req_bits_tag_T; // @[HellaCacheArbiter.scala 49:26]
  assign tag_hit = ~io_mem_resp_bits_tag[0]; // @[HellaCacheArbiter.scala 59:57]
  assign io_requestor_0_req_ready = io_mem_req_ready; // @[HellaCacheArbiter.scala 25:31]
  assign io_requestor_0_s2_nack = io_mem_s2_nack & ~s2_id; // @[HellaCacheArbiter.scala 64:31]
  assign io_requestor_0_resp_valid = io_mem_resp_valid & tag_hit; // @[HellaCacheArbiter.scala 60:18]
  assign io_requestor_0_resp_bits_data = io_mem_resp_bits_data; // @[HellaCacheArbiter.scala 69:17]
  assign io_requestor_0_s2_xcpt_ae_ld = io_mem_s2_xcpt_ae_ld; // @[HellaCacheArbiter.scala 61:31]
  assign io_requestor_1_req_ready = io_requestor_0_req_ready & ~io_requestor_0_req_valid; // @[HellaCacheArbiter.scala 27:33]
  assign io_requestor_1_s2_nack = io_mem_s2_nack & s2_id; // @[HellaCacheArbiter.scala 64:31]
  assign io_requestor_1_resp_valid = io_mem_resp_valid & io_mem_resp_bits_tag[0]; // @[HellaCacheArbiter.scala 60:18]
  assign io_requestor_1_resp_bits_tag = {{1'd0}, io_mem_resp_bits_tag[6:1]}; // @[HellaCacheArbiter.scala 69:17 HellaCacheArbiter.scala 70:21]
  assign io_requestor_1_resp_bits_size = io_mem_resp_bits_size; // @[HellaCacheArbiter.scala 69:17]
  assign io_requestor_1_resp_bits_data = io_mem_resp_bits_data; // @[HellaCacheArbiter.scala 69:17]
  assign io_requestor_1_resp_bits_replay = io_mem_resp_bits_replay; // @[HellaCacheArbiter.scala 69:17]
  assign io_requestor_1_resp_bits_has_data = io_mem_resp_bits_has_data; // @[HellaCacheArbiter.scala 69:17]
  assign io_requestor_1_resp_bits_data_word_bypass = io_mem_resp_bits_data_word_bypass; // @[HellaCacheArbiter.scala 69:17]
  assign io_requestor_1_replay_next = io_mem_replay_next; // @[HellaCacheArbiter.scala 72:35]
  assign io_requestor_1_s2_xcpt_ma_ld = io_mem_s2_xcpt_ma_ld; // @[HellaCacheArbiter.scala 61:31]
  assign io_requestor_1_s2_xcpt_ma_st = io_mem_s2_xcpt_ma_st; // @[HellaCacheArbiter.scala 61:31]
  assign io_requestor_1_s2_xcpt_pf_ld = io_mem_s2_xcpt_pf_ld; // @[HellaCacheArbiter.scala 61:31]
  assign io_requestor_1_s2_xcpt_pf_st = io_mem_s2_xcpt_pf_st; // @[HellaCacheArbiter.scala 61:31]
  assign io_requestor_1_s2_xcpt_ae_ld = io_mem_s2_xcpt_ae_ld; // @[HellaCacheArbiter.scala 61:31]
  assign io_requestor_1_s2_xcpt_ae_st = io_mem_s2_xcpt_ae_st; // @[HellaCacheArbiter.scala 61:31]
  assign io_requestor_1_ordered = io_mem_ordered; // @[HellaCacheArbiter.scala 62:31]
  assign io_requestor_1_perf_release = io_mem_perf_release; // @[HellaCacheArbiter.scala 63:28]
  assign io_requestor_1_perf_grant = io_mem_perf_grant; // @[HellaCacheArbiter.scala 63:28]
  assign io_mem_req_valid = io_requestor_0_req_valid | io_requestor_1_req_valid; // @[HellaCacheArbiter.scala 24:22]
  assign io_mem_req_bits_addr = io_requestor_0_req_valid ? io_requestor_0_req_bits_addr : io_requestor_1_req_bits_addr; // @[HellaCacheArbiter.scala 32:25 HellaCacheArbiter.scala 32:25]
  assign io_mem_req_bits_tag = _GEN_1[6:0]; // @[HellaCacheArbiter.scala 32:25 HellaCacheArbiter.scala 33:29 HellaCacheArbiter.scala 32:25 HellaCacheArbiter.scala 33:29]
  assign io_mem_req_bits_cmd = io_requestor_0_req_valid ? 5'h0 : io_requestor_1_req_bits_cmd; // @[HellaCacheArbiter.scala 32:25 HellaCacheArbiter.scala 32:25]
  assign io_mem_req_bits_size = io_requestor_0_req_valid ? 2'h3 : io_requestor_1_req_bits_size; // @[HellaCacheArbiter.scala 32:25 HellaCacheArbiter.scala 32:25]
  assign io_mem_req_bits_signed = io_requestor_0_req_valid ? 1'h0 : io_requestor_1_req_bits_signed; // @[HellaCacheArbiter.scala 32:25 HellaCacheArbiter.scala 32:25]
  assign io_mem_req_bits_phys = io_requestor_0_req_valid; // @[HellaCacheArbiter.scala 32:25 HellaCacheArbiter.scala 32:25]
  assign io_mem_s1_kill = s1_id ? io_requestor_1_s1_kill : io_requestor_0_s1_kill; // @[HellaCacheArbiter.scala 37:24 HellaCacheArbiter.scala 37:24]
  assign io_mem_s1_data_data = s1_id ? io_requestor_1_s1_data_data : 64'h0; // @[HellaCacheArbiter.scala 38:24 HellaCacheArbiter.scala 38:24]
  assign HellaCacheArbiter_cov_read_addr = HellaCacheArbiter_state;
  assign HellaCacheArbiter_cov_read_data = HellaCacheArbiter_cov[HellaCacheArbiter_cov_read_addr]; // @[Coverage map for HellaCacheArbiter]
  assign HellaCacheArbiter_cov_write_data = 1'h1;
  assign HellaCacheArbiter_cov_write_addr = HellaCacheArbiter_state;
  assign HellaCacheArbiter_cov_write_mask = 1'h1;
  assign HellaCacheArbiter_cov_write_en = 1'h1;
  assign s1_id_shl = s1_id;
  assign s1_id_pad = s1_id_shl;
  assign io_covSum = HellaCacheArbiter_covSum;
  assign metaAssert = 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s1_id = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  s2_id = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  HellaCacheArbiter_state = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    HellaCacheArbiter_cov[initvar] = _RAND_3[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  HellaCacheArbiter_covSum = _RAND_4[29:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      s1_id <= 1'h0;
    end else if (io_requestor_0_req_valid) begin
      s1_id <= 1'h0;
    end else begin
      s1_id <= 1'h1;
    end
    if (metaReset) begin
      s2_id <= 1'h0;
    end else begin
      s2_id <= s1_id;
    end
    HellaCacheArbiter_state <= s1_id_pad;
    if (!(HellaCacheArbiter_cov_read_data)) begin
      HellaCacheArbiter_covSum <= HellaCacheArbiter_covSum + 1'h1;
    end
  end
  always @(posedge clock) begin
    if(HellaCacheArbiter_cov_write_en & HellaCacheArbiter_cov_write_mask) begin
      HellaCacheArbiter_cov[HellaCacheArbiter_cov_write_addr] <= HellaCacheArbiter_cov_write_data; // @[Coverage map for HellaCacheArbiter]
    end
  end
endmodule
module PTW(
  input         clock,
  input         reset,
  output        io_requestor_0_req_ready,
  input         io_requestor_0_req_valid,
  input  [26:0] io_requestor_0_req_bits_bits_addr,
  output        io_requestor_0_resp_valid,
  output        io_requestor_0_resp_bits_ae,
  output [53:0] io_requestor_0_resp_bits_pte_ppn,
  output        io_requestor_0_resp_bits_pte_d,
  output        io_requestor_0_resp_bits_pte_a,
  output        io_requestor_0_resp_bits_pte_g,
  output        io_requestor_0_resp_bits_pte_u,
  output        io_requestor_0_resp_bits_pte_x,
  output        io_requestor_0_resp_bits_pte_w,
  output        io_requestor_0_resp_bits_pte_r,
  output        io_requestor_0_resp_bits_pte_v,
  output [1:0]  io_requestor_0_resp_bits_level,
  output        io_requestor_0_resp_bits_homogeneous,
  output [3:0]  io_requestor_0_ptbr_mode,
  output        io_requestor_0_status_debug,
  output [1:0]  io_requestor_0_status_dprv,
  output        io_requestor_0_status_mxr,
  output        io_requestor_0_status_sum,
  output        io_requestor_0_pmp_0_cfg_l,
  output [1:0]  io_requestor_0_pmp_0_cfg_a,
  output        io_requestor_0_pmp_0_cfg_x,
  output        io_requestor_0_pmp_0_cfg_w,
  output        io_requestor_0_pmp_0_cfg_r,
  output [29:0] io_requestor_0_pmp_0_addr,
  output [31:0] io_requestor_0_pmp_0_mask,
  output        io_requestor_0_pmp_1_cfg_l,
  output [1:0]  io_requestor_0_pmp_1_cfg_a,
  output        io_requestor_0_pmp_1_cfg_x,
  output        io_requestor_0_pmp_1_cfg_w,
  output        io_requestor_0_pmp_1_cfg_r,
  output [29:0] io_requestor_0_pmp_1_addr,
  output [31:0] io_requestor_0_pmp_1_mask,
  output        io_requestor_0_pmp_2_cfg_l,
  output [1:0]  io_requestor_0_pmp_2_cfg_a,
  output        io_requestor_0_pmp_2_cfg_x,
  output        io_requestor_0_pmp_2_cfg_w,
  output        io_requestor_0_pmp_2_cfg_r,
  output [29:0] io_requestor_0_pmp_2_addr,
  output [31:0] io_requestor_0_pmp_2_mask,
  output        io_requestor_0_pmp_3_cfg_l,
  output [1:0]  io_requestor_0_pmp_3_cfg_a,
  output        io_requestor_0_pmp_3_cfg_x,
  output        io_requestor_0_pmp_3_cfg_w,
  output        io_requestor_0_pmp_3_cfg_r,
  output [29:0] io_requestor_0_pmp_3_addr,
  output [31:0] io_requestor_0_pmp_3_mask,
  output        io_requestor_0_pmp_4_cfg_l,
  output [1:0]  io_requestor_0_pmp_4_cfg_a,
  output        io_requestor_0_pmp_4_cfg_x,
  output        io_requestor_0_pmp_4_cfg_w,
  output        io_requestor_0_pmp_4_cfg_r,
  output [29:0] io_requestor_0_pmp_4_addr,
  output [31:0] io_requestor_0_pmp_4_mask,
  output        io_requestor_0_pmp_5_cfg_l,
  output [1:0]  io_requestor_0_pmp_5_cfg_a,
  output        io_requestor_0_pmp_5_cfg_x,
  output        io_requestor_0_pmp_5_cfg_w,
  output        io_requestor_0_pmp_5_cfg_r,
  output [29:0] io_requestor_0_pmp_5_addr,
  output [31:0] io_requestor_0_pmp_5_mask,
  output        io_requestor_0_pmp_6_cfg_l,
  output [1:0]  io_requestor_0_pmp_6_cfg_a,
  output        io_requestor_0_pmp_6_cfg_x,
  output        io_requestor_0_pmp_6_cfg_w,
  output        io_requestor_0_pmp_6_cfg_r,
  output [29:0] io_requestor_0_pmp_6_addr,
  output [31:0] io_requestor_0_pmp_6_mask,
  output        io_requestor_0_pmp_7_cfg_l,
  output [1:0]  io_requestor_0_pmp_7_cfg_a,
  output        io_requestor_0_pmp_7_cfg_x,
  output        io_requestor_0_pmp_7_cfg_w,
  output        io_requestor_0_pmp_7_cfg_r,
  output [29:0] io_requestor_0_pmp_7_addr,
  output [31:0] io_requestor_0_pmp_7_mask,
  output        io_requestor_1_req_ready,
  input         io_requestor_1_req_valid,
  input         io_requestor_1_req_bits_valid,
  input  [26:0] io_requestor_1_req_bits_bits_addr,
  output        io_requestor_1_resp_valid,
  output        io_requestor_1_resp_bits_ae,
  output [53:0] io_requestor_1_resp_bits_pte_ppn,
  output        io_requestor_1_resp_bits_pte_d,
  output        io_requestor_1_resp_bits_pte_a,
  output        io_requestor_1_resp_bits_pte_g,
  output        io_requestor_1_resp_bits_pte_u,
  output        io_requestor_1_resp_bits_pte_x,
  output        io_requestor_1_resp_bits_pte_w,
  output        io_requestor_1_resp_bits_pte_r,
  output        io_requestor_1_resp_bits_pte_v,
  output [1:0]  io_requestor_1_resp_bits_level,
  output        io_requestor_1_resp_bits_homogeneous,
  output [3:0]  io_requestor_1_ptbr_mode,
  output        io_requestor_1_status_debug,
  output [1:0]  io_requestor_1_status_prv,
  output        io_requestor_1_pmp_0_cfg_l,
  output [1:0]  io_requestor_1_pmp_0_cfg_a,
  output        io_requestor_1_pmp_0_cfg_x,
  output        io_requestor_1_pmp_0_cfg_w,
  output        io_requestor_1_pmp_0_cfg_r,
  output [29:0] io_requestor_1_pmp_0_addr,
  output [31:0] io_requestor_1_pmp_0_mask,
  output        io_requestor_1_pmp_1_cfg_l,
  output [1:0]  io_requestor_1_pmp_1_cfg_a,
  output        io_requestor_1_pmp_1_cfg_x,
  output        io_requestor_1_pmp_1_cfg_w,
  output        io_requestor_1_pmp_1_cfg_r,
  output [29:0] io_requestor_1_pmp_1_addr,
  output [31:0] io_requestor_1_pmp_1_mask,
  output        io_requestor_1_pmp_2_cfg_l,
  output [1:0]  io_requestor_1_pmp_2_cfg_a,
  output        io_requestor_1_pmp_2_cfg_x,
  output        io_requestor_1_pmp_2_cfg_w,
  output        io_requestor_1_pmp_2_cfg_r,
  output [29:0] io_requestor_1_pmp_2_addr,
  output [31:0] io_requestor_1_pmp_2_mask,
  output        io_requestor_1_pmp_3_cfg_l,
  output [1:0]  io_requestor_1_pmp_3_cfg_a,
  output        io_requestor_1_pmp_3_cfg_x,
  output        io_requestor_1_pmp_3_cfg_w,
  output        io_requestor_1_pmp_3_cfg_r,
  output [29:0] io_requestor_1_pmp_3_addr,
  output [31:0] io_requestor_1_pmp_3_mask,
  output        io_requestor_1_pmp_4_cfg_l,
  output [1:0]  io_requestor_1_pmp_4_cfg_a,
  output        io_requestor_1_pmp_4_cfg_x,
  output        io_requestor_1_pmp_4_cfg_w,
  output        io_requestor_1_pmp_4_cfg_r,
  output [29:0] io_requestor_1_pmp_4_addr,
  output [31:0] io_requestor_1_pmp_4_mask,
  output        io_requestor_1_pmp_5_cfg_l,
  output [1:0]  io_requestor_1_pmp_5_cfg_a,
  output        io_requestor_1_pmp_5_cfg_x,
  output        io_requestor_1_pmp_5_cfg_w,
  output        io_requestor_1_pmp_5_cfg_r,
  output [29:0] io_requestor_1_pmp_5_addr,
  output [31:0] io_requestor_1_pmp_5_mask,
  output        io_requestor_1_pmp_6_cfg_l,
  output [1:0]  io_requestor_1_pmp_6_cfg_a,
  output        io_requestor_1_pmp_6_cfg_x,
  output        io_requestor_1_pmp_6_cfg_w,
  output        io_requestor_1_pmp_6_cfg_r,
  output [29:0] io_requestor_1_pmp_6_addr,
  output [31:0] io_requestor_1_pmp_6_mask,
  output        io_requestor_1_pmp_7_cfg_l,
  output [1:0]  io_requestor_1_pmp_7_cfg_a,
  output        io_requestor_1_pmp_7_cfg_x,
  output        io_requestor_1_pmp_7_cfg_w,
  output        io_requestor_1_pmp_7_cfg_r,
  output [29:0] io_requestor_1_pmp_7_addr,
  output [31:0] io_requestor_1_pmp_7_mask,
  output [63:0] io_requestor_1_customCSRs_csrs_0_value,
  input         io_mem_req_ready,
  output        io_mem_req_valid,
  output [39:0] io_mem_req_bits_addr,
  output        io_mem_s1_kill,
  input         io_mem_s2_nack,
  input         io_mem_resp_valid,
  input  [63:0] io_mem_resp_bits_data,
  input         io_mem_s2_xcpt_ae_ld,
  input  [3:0]  io_dpath_ptbr_mode,
  input  [43:0] io_dpath_ptbr_ppn,
  input         io_dpath_sfence_valid,
  input         io_dpath_sfence_bits_rs1,
  input         io_dpath_status_debug,
  input  [1:0]  io_dpath_status_dprv,
  input  [1:0]  io_dpath_status_prv,
  input         io_dpath_status_mxr,
  input         io_dpath_status_sum,
  input         io_dpath_pmp_0_cfg_l,
  input  [1:0]  io_dpath_pmp_0_cfg_a,
  input         io_dpath_pmp_0_cfg_x,
  input         io_dpath_pmp_0_cfg_w,
  input         io_dpath_pmp_0_cfg_r,
  input  [29:0] io_dpath_pmp_0_addr,
  input  [31:0] io_dpath_pmp_0_mask,
  input         io_dpath_pmp_1_cfg_l,
  input  [1:0]  io_dpath_pmp_1_cfg_a,
  input         io_dpath_pmp_1_cfg_x,
  input         io_dpath_pmp_1_cfg_w,
  input         io_dpath_pmp_1_cfg_r,
  input  [29:0] io_dpath_pmp_1_addr,
  input  [31:0] io_dpath_pmp_1_mask,
  input         io_dpath_pmp_2_cfg_l,
  input  [1:0]  io_dpath_pmp_2_cfg_a,
  input         io_dpath_pmp_2_cfg_x,
  input         io_dpath_pmp_2_cfg_w,
  input         io_dpath_pmp_2_cfg_r,
  input  [29:0] io_dpath_pmp_2_addr,
  input  [31:0] io_dpath_pmp_2_mask,
  input         io_dpath_pmp_3_cfg_l,
  input  [1:0]  io_dpath_pmp_3_cfg_a,
  input         io_dpath_pmp_3_cfg_x,
  input         io_dpath_pmp_3_cfg_w,
  input         io_dpath_pmp_3_cfg_r,
  input  [29:0] io_dpath_pmp_3_addr,
  input  [31:0] io_dpath_pmp_3_mask,
  input         io_dpath_pmp_4_cfg_l,
  input  [1:0]  io_dpath_pmp_4_cfg_a,
  input         io_dpath_pmp_4_cfg_x,
  input         io_dpath_pmp_4_cfg_w,
  input         io_dpath_pmp_4_cfg_r,
  input  [29:0] io_dpath_pmp_4_addr,
  input  [31:0] io_dpath_pmp_4_mask,
  input         io_dpath_pmp_5_cfg_l,
  input  [1:0]  io_dpath_pmp_5_cfg_a,
  input         io_dpath_pmp_5_cfg_x,
  input         io_dpath_pmp_5_cfg_w,
  input         io_dpath_pmp_5_cfg_r,
  input  [29:0] io_dpath_pmp_5_addr,
  input  [31:0] io_dpath_pmp_5_mask,
  input         io_dpath_pmp_6_cfg_l,
  input  [1:0]  io_dpath_pmp_6_cfg_a,
  input         io_dpath_pmp_6_cfg_x,
  input         io_dpath_pmp_6_cfg_w,
  input         io_dpath_pmp_6_cfg_r,
  input  [29:0] io_dpath_pmp_6_addr,
  input  [31:0] io_dpath_pmp_6_mask,
  input         io_dpath_pmp_7_cfg_l,
  input  [1:0]  io_dpath_pmp_7_cfg_a,
  input         io_dpath_pmp_7_cfg_x,
  input         io_dpath_pmp_7_cfg_w,
  input         io_dpath_pmp_7_cfg_r,
  input  [29:0] io_dpath_pmp_7_addr,
  input  [31:0] io_dpath_pmp_7_mask,
  output        io_dpath_perf_l2hit,
  output        io_dpath_perf_pte_miss,
  output        io_dpath_perf_pte_hit,
  input  [63:0] io_dpath_customCSRs_csrs_0_value,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  wire  arb_io_in_0_ready; // @[PTW.scala 112:19]
  wire  arb_io_in_0_valid; // @[PTW.scala 112:19]
  wire [26:0] arb_io_in_0_bits_bits_addr; // @[PTW.scala 112:19]
  wire  arb_io_in_1_ready; // @[PTW.scala 112:19]
  wire  arb_io_in_1_valid; // @[PTW.scala 112:19]
  wire  arb_io_in_1_bits_valid; // @[PTW.scala 112:19]
  wire [26:0] arb_io_in_1_bits_bits_addr; // @[PTW.scala 112:19]
  wire  arb_io_out_ready; // @[PTW.scala 112:19]
  wire  arb_io_out_valid; // @[PTW.scala 112:19]
  wire  arb_io_out_bits_valid; // @[PTW.scala 112:19]
  wire [26:0] arb_io_out_bits_bits_addr; // @[PTW.scala 112:19]
  wire  arb_io_chosen; // @[PTW.scala 112:19]
  wire [29:0] arb_io_covSum; // @[PTW.scala 112:19]
  wire  arb_metaAssert; // @[PTW.scala 112:19]
  wire [2:0] state_barrier_io_x; // @[package.scala 258:25]
  wire [2:0] state_barrier_io_y; // @[package.scala 258:25]
  wire [29:0] state_barrier_io_covSum; // @[package.scala 258:25]
  wire  state_barrier_metaAssert; // @[package.scala 258:25]
  wire [53:0] r_pte_barrier_io_x_ppn; // @[package.scala 258:25]
  wire  r_pte_barrier_io_x_d; // @[package.scala 258:25]
  wire  r_pte_barrier_io_x_a; // @[package.scala 258:25]
  wire  r_pte_barrier_io_x_g; // @[package.scala 258:25]
  wire  r_pte_barrier_io_x_u; // @[package.scala 258:25]
  wire  r_pte_barrier_io_x_x; // @[package.scala 258:25]
  wire  r_pte_barrier_io_x_w; // @[package.scala 258:25]
  wire  r_pte_barrier_io_x_r; // @[package.scala 258:25]
  wire  r_pte_barrier_io_x_v; // @[package.scala 258:25]
  wire [53:0] r_pte_barrier_io_y_ppn; // @[package.scala 258:25]
  wire  r_pte_barrier_io_y_d; // @[package.scala 258:25]
  wire  r_pte_barrier_io_y_a; // @[package.scala 258:25]
  wire  r_pte_barrier_io_y_g; // @[package.scala 258:25]
  wire  r_pte_barrier_io_y_u; // @[package.scala 258:25]
  wire  r_pte_barrier_io_y_x; // @[package.scala 258:25]
  wire  r_pte_barrier_io_y_w; // @[package.scala 258:25]
  wire  r_pte_barrier_io_y_r; // @[package.scala 258:25]
  wire  r_pte_barrier_io_y_v; // @[package.scala 258:25]
  wire [29:0] r_pte_barrier_io_covSum; // @[package.scala 258:25]
  wire  r_pte_barrier_metaAssert; // @[package.scala 258:25]
  reg [2:0] state; // @[PTW.scala 109:18]
  reg [31:0] _RAND_0;
  wire  _arb_io_out_ready_T; // @[PTW.scala 114:30]
  reg  l2_refill; // @[PTW.scala 201:26]
  reg [31:0] _RAND_1;
  reg  resp_valid_0; // @[PTW.scala 116:23]
  reg [31:0] _RAND_2;
  reg  resp_valid_1; // @[PTW.scala 116:23]
  reg [31:0] _RAND_3;
  wire  _clock_en_T; // @[PTW.scala 118:24]
  reg  invalidated; // @[PTW.scala 125:24]
  reg [31:0] _RAND_4;
  reg [1:0] count; // @[PTW.scala 126:18]
  reg [31:0] _RAND_5;
  reg  resp_ae; // @[PTW.scala 127:24]
  reg [31:0] _RAND_6;
  reg [26:0] r_req_addr; // @[PTW.scala 130:18]
  reg [31:0] _RAND_7;
  reg  r_req_dest; // @[PTW.scala 131:23]
  reg [31:0] _RAND_8;
  reg [53:0] r_pte_ppn; // @[PTW.scala 132:18]
  reg [63:0] _RAND_9;
  reg  r_pte_d; // @[PTW.scala 132:18]
  reg [31:0] _RAND_10;
  reg  r_pte_a; // @[PTW.scala 132:18]
  reg [31:0] _RAND_11;
  reg  r_pte_g; // @[PTW.scala 132:18]
  reg [31:0] _RAND_12;
  reg  r_pte_u; // @[PTW.scala 132:18]
  reg [31:0] _RAND_13;
  reg  r_pte_x; // @[PTW.scala 132:18]
  reg [31:0] _RAND_14;
  reg  r_pte_w; // @[PTW.scala 132:18]
  reg [31:0] _RAND_15;
  reg  r_pte_r; // @[PTW.scala 132:18]
  reg [31:0] _RAND_16;
  reg  r_pte_v; // @[PTW.scala 132:18]
  reg [31:0] _RAND_17;
  reg  mem_resp_valid; // @[PTW.scala 134:31]
  reg [31:0] _RAND_18;
  reg [63:0] mem_resp_data; // @[PTW.scala 135:30]
  reg [63:0] _RAND_19;
  wire  tmp_v; // @[PTW.scala 146:33]
  wire  tmp_r; // @[PTW.scala 146:33]
  wire  tmp_w; // @[PTW.scala 146:33]
  wire  tmp_x; // @[PTW.scala 146:33]
  wire  tmp_u; // @[PTW.scala 146:33]
  wire  tmp_g; // @[PTW.scala 146:33]
  wire  tmp_a; // @[PTW.scala 146:33]
  wire  tmp_d; // @[PTW.scala 146:33]
  wire [53:0] tmp_ppn; // @[PTW.scala 146:33]
  wire  _T_11; // @[PTW.scala 149:17]
  wire  _T_12; // @[PTW.scala 149:26]
  wire  _T_13; // @[PTW.scala 152:21]
  wire  _T_15; // @[PTW.scala 152:95]
  wire  _T_16; // @[PTW.scala 152:26]
  wire  _GEN_0; // @[PTW.scala 152:102]
  wire  _T_17; // @[PTW.scala 152:21]
  wire  _T_19; // @[PTW.scala 152:95]
  wire  _T_20; // @[PTW.scala 152:26]
  wire  _GEN_1; // @[PTW.scala 152:102]
  wire  res_v; // @[PTW.scala 149:36]
  wire  invalid_paddr; // @[PTW.scala 154:32]
  wire  _traverse_T_1; // @[PTW.scala 72:33]
  wire  _traverse_T_3; // @[PTW.scala 72:39]
  wire  _traverse_T_5; // @[PTW.scala 72:45]
  wire  _traverse_T_7; // @[PTW.scala 156:30]
  wire  _traverse_T_8; // @[PTW.scala 156:57]
  wire  traverse; // @[PTW.scala 156:48]
  wire [8:0] vpn_idxs_0; // @[PTW.scala 158:60]
  wire [8:0] vpn_idxs_1; // @[PTW.scala 158:90]
  wire [8:0] vpn_idxs_2; // @[PTW.scala 158:90]
  wire  _pte_addr_vpn_idx_T; // @[package.scala 32:86]
  wire [8:0] _pte_addr_vpn_idx_T_1; // @[package.scala 32:76]
  wire  _pte_addr_vpn_idx_T_2; // @[package.scala 32:86]
  wire [8:0] _pte_addr_vpn_idx_T_3; // @[package.scala 32:76]
  wire  _pte_addr_vpn_idx_T_4; // @[package.scala 32:86]
  wire [8:0] vpn_idx; // @[package.scala 32:76]
  wire [62:0] _pte_addr_T; // @[Cat.scala 30:58]
  wire [65:0] pte_addr; // @[PTW.scala 160:29]
  wire [35:0] fragmented_superpage_ppn_choices_hi; // @[PTW.scala 163:69]
  wire [17:0] fragmented_superpage_ppn_choices_lo; // @[PTW.scala 163:99]
  wire [53:0] choices_0; // @[Cat.scala 30:58]
  wire [44:0] fragmented_superpage_ppn_choices_hi_1; // @[PTW.scala 163:69]
  wire [53:0] choices_1; // @[Cat.scala 30:58]
  wire  fragmented_superpage_ppn_truncIdx; // @[package.scala 31:49]
  wire [53:0] fragmented_superpage_ppn; // @[package.scala 32:76]
  wire  _T_22; // @[Decoupled.scala 40:37]
  reg [6:0] state_reg; // @[Replacement.scala 168:70]
  reg [31:0] _RAND_20;
  reg [7:0] valid; // @[PTW.scala 175:24]
  reg [31:0] _RAND_21;
  reg [31:0] tags_0; // @[PTW.scala 176:19]
  reg [31:0] _RAND_22;
  reg [31:0] tags_1; // @[PTW.scala 176:19]
  reg [31:0] _RAND_23;
  reg [31:0] tags_2; // @[PTW.scala 176:19]
  reg [31:0] _RAND_24;
  reg [31:0] tags_3; // @[PTW.scala 176:19]
  reg [31:0] _RAND_25;
  reg [31:0] tags_4; // @[PTW.scala 176:19]
  reg [31:0] _RAND_26;
  reg [31:0] tags_5; // @[PTW.scala 176:19]
  reg [31:0] _RAND_27;
  reg [31:0] tags_6; // @[PTW.scala 176:19]
  reg [31:0] _RAND_28;
  reg [31:0] tags_7; // @[PTW.scala 176:19]
  reg [31:0] _RAND_29;
  reg [19:0] data_0; // @[PTW.scala 177:19]
  reg [31:0] _RAND_30;
  reg [19:0] data_1; // @[PTW.scala 177:19]
  reg [31:0] _RAND_31;
  reg [19:0] data_2; // @[PTW.scala 177:19]
  reg [31:0] _RAND_32;
  reg [19:0] data_3; // @[PTW.scala 177:19]
  reg [31:0] _RAND_33;
  reg [19:0] data_4; // @[PTW.scala 177:19]
  reg [31:0] _RAND_34;
  reg [19:0] data_5; // @[PTW.scala 177:19]
  reg [31:0] _RAND_35;
  reg [19:0] data_6; // @[PTW.scala 177:19]
  reg [31:0] _RAND_36;
  reg [19:0] data_7; // @[PTW.scala 177:19]
  reg [31:0] _RAND_37;
  wire [65:0] _GEN_115; // @[PTW.scala 179:27]
  wire  lo_lo_lo; // @[PTW.scala 179:27]
  wire [65:0] _GEN_116; // @[PTW.scala 179:27]
  wire  lo_lo_hi; // @[PTW.scala 179:27]
  wire [65:0] _GEN_117; // @[PTW.scala 179:27]
  wire  lo_hi_lo; // @[PTW.scala 179:27]
  wire [65:0] _GEN_118; // @[PTW.scala 179:27]
  wire  lo_hi_hi; // @[PTW.scala 179:27]
  wire [65:0] _GEN_119; // @[PTW.scala 179:27]
  wire  hi_lo_lo; // @[PTW.scala 179:27]
  wire [65:0] _GEN_120; // @[PTW.scala 179:27]
  wire  hi_lo_hi; // @[PTW.scala 179:27]
  wire [65:0] _GEN_121; // @[PTW.scala 179:27]
  wire  hi_hi_lo; // @[PTW.scala 179:27]
  wire [65:0] _GEN_122; // @[PTW.scala 179:27]
  wire  hi_hi_hi; // @[PTW.scala 179:27]
  wire [7:0] _T_23; // @[Cat.scala 30:58]
  wire [7:0] hits; // @[PTW.scala 179:48]
  wire  hit; // @[PTW.scala 180:20]
  wire  _T_24; // @[PTW.scala 181:26]
  wire  _T_26; // @[PTW.scala 181:38]
  wire  _T_28; // @[PTW.scala 181:46]
  wire  _T_29; // @[PTW.scala 182:25]
  wire  hi_1; // @[Replacement.scala 243:38]
  wire [2:0] left_subtree_state; // @[package.scala 154:13]
  wire [2:0] right_subtree_state; // @[Replacement.scala 245:38]
  wire  hi_2; // @[Replacement.scala 243:38]
  wire  left_subtree_state_1; // @[package.scala 154:13]
  wire  right_subtree_state_1; // @[Replacement.scala 245:38]
  wire  lo_1; // @[Replacement.scala 250:16]
  wire [1:0] _T_32; // @[Cat.scala 30:58]
  wire  hi_3; // @[Replacement.scala 243:38]
  wire  left_subtree_state_2; // @[package.scala 154:13]
  wire  right_subtree_state_2; // @[Replacement.scala 245:38]
  wire  lo_2; // @[Replacement.scala 250:16]
  wire [1:0] _T_35; // @[Cat.scala 30:58]
  wire [1:0] lo_3; // @[Replacement.scala 250:16]
  wire [2:0] _T_36; // @[Cat.scala 30:58]
  wire  _T_38; // @[OneHot.scala 47:40]
  wire  _T_39; // @[OneHot.scala 47:40]
  wire  _T_40; // @[OneHot.scala 47:40]
  wire  _T_41; // @[OneHot.scala 47:40]
  wire  _T_42; // @[OneHot.scala 47:40]
  wire  _T_43; // @[OneHot.scala 47:40]
  wire  _T_44; // @[OneHot.scala 47:40]
  wire [2:0] _T_46; // @[Mux.scala 47:69]
  wire [2:0] _T_47; // @[Mux.scala 47:69]
  wire [2:0] _T_48; // @[Mux.scala 47:69]
  wire [2:0] _T_49; // @[Mux.scala 47:69]
  wire [2:0] _T_50; // @[Mux.scala 47:69]
  wire [2:0] _T_51; // @[Mux.scala 47:69]
  wire [2:0] _T_52; // @[Mux.scala 47:69]
  wire [2:0] r; // @[PTW.scala 182:18]
  wire [7:0] _T_53; // @[OneHot.scala 58:35]
  wire [7:0] _T_54; // @[PTW.scala 183:22]
  wire [53:0] res_ppn; // @[PTW.scala 148:13]
  wire  _T_55; // @[PTW.scala 187:24]
  wire  _T_56; // @[PTW.scala 187:15]
  wire [3:0] hi_4; // @[OneHot.scala 30:18]
  wire [3:0] lo_4; // @[OneHot.scala 31:18]
  wire  hi_5; // @[OneHot.scala 32:14]
  wire [3:0] _T_57; // @[OneHot.scala 32:28]
  wire [1:0] hi_6; // @[OneHot.scala 30:18]
  wire [1:0] lo_5; // @[OneHot.scala 31:18]
  wire  hi_7; // @[OneHot.scala 32:14]
  wire [1:0] _T_58; // @[OneHot.scala 32:28]
  wire  lo_6; // @[CircuitMath.scala 30:8]
  wire [2:0] state_reg_touch_way_sized; // @[Cat.scala 30:58]
  wire  state_reg_hi_hi; // @[Replacement.scala 196:33]
  wire  state_reg_hi_hi_1; // @[Replacement.scala 196:33]
  wire  state_reg_hi_lo; // @[Replacement.scala 203:16]
  wire  state_reg_lo; // @[Replacement.scala 206:16]
  wire [2:0] _state_reg_T_7; // @[Cat.scala 30:58]
  wire [2:0] state_reg_hi_lo_1; // @[Replacement.scala 203:16]
  wire  state_reg_hi_lo_2; // @[Replacement.scala 203:16]
  wire  state_reg_lo_1; // @[Replacement.scala 206:16]
  wire [2:0] _state_reg_T_15; // @[Cat.scala 30:58]
  wire [2:0] state_reg_lo_2; // @[Replacement.scala 206:16]
  wire [6:0] _state_reg_T_16; // @[Cat.scala 30:58]
  wire  _T_61; // @[PTW.scala 188:33]
  wire  pte_cache_hit; // @[PTW.scala 193:10]
  wire [19:0] _T_79; // @[Mux.scala 27:72]
  wire [19:0] _T_80; // @[Mux.scala 27:72]
  wire [19:0] _T_81; // @[Mux.scala 27:72]
  wire [19:0] _T_82; // @[Mux.scala 27:72]
  wire [19:0] _T_83; // @[Mux.scala 27:72]
  wire [19:0] _T_84; // @[Mux.scala 27:72]
  wire [19:0] _T_85; // @[Mux.scala 27:72]
  wire [19:0] _T_86; // @[Mux.scala 27:72]
  wire [19:0] _T_87; // @[Mux.scala 27:72]
  wire [19:0] _T_88; // @[Mux.scala 27:72]
  wire [19:0] _T_89; // @[Mux.scala 27:72]
  wire [19:0] _T_90; // @[Mux.scala 27:72]
  wire [19:0] _T_91; // @[Mux.scala 27:72]
  wire [19:0] _T_92; // @[Mux.scala 27:72]
  wire [19:0] pte_cache_data; // @[Mux.scala 27:72]
  reg  pte_hit; // @[PTW.scala 195:24]
  reg [31:0] _RAND_38;
  wire  _io_dpath_perf_pte_hit_T_1; // @[PTW.scala 197:36]
  wire  _T_94; // @[PTW.scala 198:59]
  wire  _T_95; // @[PTW.scala 198:32]
  wire  _T_98; // @[PTW.scala 198:9]
  wire  _invalidated_T_1; // @[PTW.scala 285:56]
  wire  _io_mem_req_valid_T_1; // @[PTW.scala 287:48]
  wire [65:0] _pmaPgLevelHomogeneous_T_6; // @[Parameters.scala 137:31]
  wire [66:0] _pmaPgLevelHomogeneous_T_7; // @[Parameters.scala 137:49]
  wire [66:0] _pmaPgLevelHomogeneous_T_9; // @[Parameters.scala 137:52]
  wire  _pmaPgLevelHomogeneous_T_10; // @[Parameters.scala 137:67]
  wire [65:0] _pmaPgLevelHomogeneous_T_11; // @[Parameters.scala 137:31]
  wire [66:0] _pmaPgLevelHomogeneous_T_12; // @[Parameters.scala 137:49]
  wire [66:0] _pmaPgLevelHomogeneous_T_14; // @[Parameters.scala 137:52]
  wire  _pmaPgLevelHomogeneous_T_15; // @[Parameters.scala 137:67]
  wire [65:0] _pmaPgLevelHomogeneous_T_16; // @[Parameters.scala 137:31]
  wire [66:0] _pmaPgLevelHomogeneous_T_17; // @[Parameters.scala 137:49]
  wire [66:0] _pmaPgLevelHomogeneous_T_19; // @[Parameters.scala 137:52]
  wire  _pmaPgLevelHomogeneous_T_20; // @[Parameters.scala 137:67]
  wire  _pmaPgLevelHomogeneous_T_22; // @[TLBPermissions.scala 99:65]
  wire  pmaPgLevelHomogeneous_1; // @[TLBPermissions.scala 99:65]
  wire [66:0] _pmaPgLevelHomogeneous_T_26; // @[Parameters.scala 137:49]
  wire [66:0] _pmaPgLevelHomogeneous_T_53; // @[Parameters.scala 137:52]
  wire  _pmaPgLevelHomogeneous_T_54; // @[Parameters.scala 137:67]
  wire [65:0] _pmaPgLevelHomogeneous_T_55; // @[Parameters.scala 137:31]
  wire [66:0] _pmaPgLevelHomogeneous_T_56; // @[Parameters.scala 137:49]
  wire [66:0] _pmaPgLevelHomogeneous_T_58; // @[Parameters.scala 137:52]
  wire  _pmaPgLevelHomogeneous_T_59; // @[Parameters.scala 137:67]
  wire [65:0] _pmaPgLevelHomogeneous_T_60; // @[Parameters.scala 137:31]
  wire [66:0] _pmaPgLevelHomogeneous_T_61; // @[Parameters.scala 137:49]
  wire [66:0] _pmaPgLevelHomogeneous_T_63; // @[Parameters.scala 137:52]
  wire  _pmaPgLevelHomogeneous_T_64; // @[Parameters.scala 137:67]
  wire [65:0] _pmaPgLevelHomogeneous_T_65; // @[Parameters.scala 137:31]
  wire [66:0] _pmaPgLevelHomogeneous_T_66; // @[Parameters.scala 137:49]
  wire [66:0] _pmaPgLevelHomogeneous_T_68; // @[Parameters.scala 137:52]
  wire  _pmaPgLevelHomogeneous_T_69; // @[Parameters.scala 137:67]
  wire  _pmaPgLevelHomogeneous_T_86; // @[TLBPermissions.scala 99:65]
  wire  _pmaPgLevelHomogeneous_T_87; // @[TLBPermissions.scala 99:65]
  wire  _pmaPgLevelHomogeneous_T_88; // @[TLBPermissions.scala 99:65]
  wire  _pmaPgLevelHomogeneous_T_89; // @[TLBPermissions.scala 99:65]
  wire  _pmaPgLevelHomogeneous_T_90; // @[TLBPermissions.scala 99:65]
  wire  pmaPgLevelHomogeneous_2; // @[TLBPermissions.scala 99:65]
  wire  _pmaHomogeneous_T_1; // @[package.scala 32:76]
  wire  _pmaHomogeneous_T_3; // @[package.scala 32:76]
  wire  pmaHomogeneous; // @[package.scala 32:76]
  wire [65:0] _pmpHomogeneous_T_1; // @[PTW.scala 309:92]
  wire  _pmpHomogeneous_maskHomogeneous_T_4; // @[package.scala 32:76]
  wire  _pmpHomogeneous_maskHomogeneous_T_6; // @[package.scala 32:76]
  wire  pmpHomogeneous_maskHomogeneous; // @[package.scala 32:76]
  wire [31:0] _pmpHomogeneous_T_3; // @[PMP.scala 62:36]
  wire [31:0] _pmpHomogeneous_T_5; // @[PMP.scala 62:48]
  wire [65:0] _GEN_123; // @[PMP.scala 100:53]
  wire [65:0] _pmpHomogeneous_T_7; // @[PMP.scala 100:53]
  wire  _pmpHomogeneous_T_9; // @[PMP.scala 100:78]
  wire  _pmpHomogeneous_T_16; // @[PMP.scala 100:78]
  wire  _pmpHomogeneous_T_23; // @[PMP.scala 100:78]
  wire  _pmpHomogeneous_T_25; // @[package.scala 32:76]
  wire  _pmpHomogeneous_T_27; // @[package.scala 32:76]
  wire  _pmpHomogeneous_T_29; // @[package.scala 32:76]
  wire  _pmpHomogeneous_T_30; // @[PMP.scala 100:21]
  wire  _pmpHomogeneous_beginsAfterUpper_T_4; // @[PMP.scala 109:32]
  wire  pmpHomogeneous_beginsAfterUpper; // @[PMP.scala 109:28]
  wire [31:0] _pmpHomogeneous_pgMask_T_1; // @[package.scala 32:76]
  wire [31:0] _pmpHomogeneous_pgMask_T_3; // @[package.scala 32:76]
  wire [31:0] pmpHomogeneous_pgMask; // @[package.scala 32:76]
  wire [65:0] _GEN_127; // @[PMP.scala 112:30]
  wire [65:0] _pmpHomogeneous_endsBeforeLower_T; // @[PMP.scala 112:30]
  wire [31:0] _pmpHomogeneous_endsBeforeUpper_T_5; // @[PMP.scala 113:53]
  wire [65:0] _GEN_129; // @[PMP.scala 113:40]
  wire  pmpHomogeneous_endsBeforeUpper; // @[PMP.scala 113:40]
  wire  _pmpHomogeneous_T_35; // @[PMP.scala 115:41]
  wire  _pmpHomogeneous_T_36; // @[PMP.scala 120:58]
  wire  _pmpHomogeneous_T_37; // @[PMP.scala 120:8]
  wire  _pmpHomogeneous_maskHomogeneous_T_12; // @[package.scala 32:76]
  wire  _pmpHomogeneous_maskHomogeneous_T_14; // @[package.scala 32:76]
  wire  pmpHomogeneous_maskHomogeneous_1; // @[package.scala 32:76]
  wire [31:0] _pmpHomogeneous_T_40; // @[PMP.scala 62:36]
  wire [31:0] _pmpHomogeneous_T_42; // @[PMP.scala 62:48]
  wire [65:0] _GEN_130; // @[PMP.scala 100:53]
  wire [65:0] _pmpHomogeneous_T_44; // @[PMP.scala 100:53]
  wire  _pmpHomogeneous_T_46; // @[PMP.scala 100:78]
  wire  _pmpHomogeneous_T_53; // @[PMP.scala 100:78]
  wire  _pmpHomogeneous_T_60; // @[PMP.scala 100:78]
  wire  _pmpHomogeneous_T_62; // @[package.scala 32:76]
  wire  _pmpHomogeneous_T_64; // @[package.scala 32:76]
  wire  _pmpHomogeneous_T_66; // @[package.scala 32:76]
  wire  _pmpHomogeneous_T_67; // @[PMP.scala 100:21]
  wire  _pmpHomogeneous_beginsAfterUpper_T_9; // @[PMP.scala 109:32]
  wire  pmpHomogeneous_beginsAfterUpper_1; // @[PMP.scala 109:28]
  wire [31:0] _pmpHomogeneous_endsBeforeUpper_T_11; // @[PMP.scala 113:53]
  wire [65:0] _GEN_138; // @[PMP.scala 113:40]
  wire  pmpHomogeneous_endsBeforeUpper_1; // @[PMP.scala 113:40]
  wire  _pmpHomogeneous_T_70; // @[PMP.scala 115:21]
  wire  _pmpHomogeneous_T_71; // @[PMP.scala 115:62]
  wire  _pmpHomogeneous_T_72; // @[PMP.scala 115:41]
  wire  _pmpHomogeneous_T_73; // @[PMP.scala 120:58]
  wire  _pmpHomogeneous_T_74; // @[PMP.scala 120:8]
  wire  _pmpHomogeneous_T_75; // @[PMP.scala 140:10]
  wire  _pmpHomogeneous_maskHomogeneous_T_20; // @[package.scala 32:76]
  wire  _pmpHomogeneous_maskHomogeneous_T_22; // @[package.scala 32:76]
  wire  pmpHomogeneous_maskHomogeneous_2; // @[package.scala 32:76]
  wire [31:0] _pmpHomogeneous_T_77; // @[PMP.scala 62:36]
  wire [31:0] _pmpHomogeneous_T_79; // @[PMP.scala 62:48]
  wire [65:0] _GEN_139; // @[PMP.scala 100:53]
  wire [65:0] _pmpHomogeneous_T_81; // @[PMP.scala 100:53]
  wire  _pmpHomogeneous_T_83; // @[PMP.scala 100:78]
  wire  _pmpHomogeneous_T_90; // @[PMP.scala 100:78]
  wire  _pmpHomogeneous_T_97; // @[PMP.scala 100:78]
  wire  _pmpHomogeneous_T_99; // @[package.scala 32:76]
  wire  _pmpHomogeneous_T_101; // @[package.scala 32:76]
  wire  _pmpHomogeneous_T_103; // @[package.scala 32:76]
  wire  _pmpHomogeneous_T_104; // @[PMP.scala 100:21]
  wire  _pmpHomogeneous_beginsAfterUpper_T_14; // @[PMP.scala 109:32]
  wire  pmpHomogeneous_beginsAfterUpper_2; // @[PMP.scala 109:28]
  wire [31:0] _pmpHomogeneous_endsBeforeUpper_T_17; // @[PMP.scala 113:53]
  wire [65:0] _GEN_147; // @[PMP.scala 113:40]
  wire  pmpHomogeneous_endsBeforeUpper_2; // @[PMP.scala 113:40]
  wire  _pmpHomogeneous_T_107; // @[PMP.scala 115:21]
  wire  _pmpHomogeneous_T_108; // @[PMP.scala 115:62]
  wire  _pmpHomogeneous_T_109; // @[PMP.scala 115:41]
  wire  _pmpHomogeneous_T_110; // @[PMP.scala 120:58]
  wire  _pmpHomogeneous_T_111; // @[PMP.scala 120:8]
  wire  _pmpHomogeneous_T_112; // @[PMP.scala 140:10]
  wire  _pmpHomogeneous_maskHomogeneous_T_28; // @[package.scala 32:76]
  wire  _pmpHomogeneous_maskHomogeneous_T_30; // @[package.scala 32:76]
  wire  pmpHomogeneous_maskHomogeneous_3; // @[package.scala 32:76]
  wire [31:0] _pmpHomogeneous_T_114; // @[PMP.scala 62:36]
  wire [31:0] _pmpHomogeneous_T_116; // @[PMP.scala 62:48]
  wire [65:0] _GEN_148; // @[PMP.scala 100:53]
  wire [65:0] _pmpHomogeneous_T_118; // @[PMP.scala 100:53]
  wire  _pmpHomogeneous_T_120; // @[PMP.scala 100:78]
  wire  _pmpHomogeneous_T_127; // @[PMP.scala 100:78]
  wire  _pmpHomogeneous_T_134; // @[PMP.scala 100:78]
  wire  _pmpHomogeneous_T_136; // @[package.scala 32:76]
  wire  _pmpHomogeneous_T_138; // @[package.scala 32:76]
  wire  _pmpHomogeneous_T_140; // @[package.scala 32:76]
  wire  _pmpHomogeneous_T_141; // @[PMP.scala 100:21]
  wire  _pmpHomogeneous_beginsAfterUpper_T_19; // @[PMP.scala 109:32]
  wire  pmpHomogeneous_beginsAfterUpper_3; // @[PMP.scala 109:28]
  wire [31:0] _pmpHomogeneous_endsBeforeUpper_T_23; // @[PMP.scala 113:53]
  wire [65:0] _GEN_156; // @[PMP.scala 113:40]
  wire  pmpHomogeneous_endsBeforeUpper_3; // @[PMP.scala 113:40]
  wire  _pmpHomogeneous_T_144; // @[PMP.scala 115:21]
  wire  _pmpHomogeneous_T_145; // @[PMP.scala 115:62]
  wire  _pmpHomogeneous_T_146; // @[PMP.scala 115:41]
  wire  _pmpHomogeneous_T_147; // @[PMP.scala 120:58]
  wire  _pmpHomogeneous_T_148; // @[PMP.scala 120:8]
  wire  _pmpHomogeneous_T_149; // @[PMP.scala 140:10]
  wire  _pmpHomogeneous_maskHomogeneous_T_36; // @[package.scala 32:76]
  wire  _pmpHomogeneous_maskHomogeneous_T_38; // @[package.scala 32:76]
  wire  pmpHomogeneous_maskHomogeneous_4; // @[package.scala 32:76]
  wire [31:0] _pmpHomogeneous_T_151; // @[PMP.scala 62:36]
  wire [31:0] _pmpHomogeneous_T_153; // @[PMP.scala 62:48]
  wire [65:0] _GEN_157; // @[PMP.scala 100:53]
  wire [65:0] _pmpHomogeneous_T_155; // @[PMP.scala 100:53]
  wire  _pmpHomogeneous_T_157; // @[PMP.scala 100:78]
  wire  _pmpHomogeneous_T_164; // @[PMP.scala 100:78]
  wire  _pmpHomogeneous_T_171; // @[PMP.scala 100:78]
  wire  _pmpHomogeneous_T_173; // @[package.scala 32:76]
  wire  _pmpHomogeneous_T_175; // @[package.scala 32:76]
  wire  _pmpHomogeneous_T_177; // @[package.scala 32:76]
  wire  _pmpHomogeneous_T_178; // @[PMP.scala 100:21]
  wire  _pmpHomogeneous_beginsAfterUpper_T_24; // @[PMP.scala 109:32]
  wire  pmpHomogeneous_beginsAfterUpper_4; // @[PMP.scala 109:28]
  wire [31:0] _pmpHomogeneous_endsBeforeUpper_T_29; // @[PMP.scala 113:53]
  wire [65:0] _GEN_165; // @[PMP.scala 113:40]
  wire  pmpHomogeneous_endsBeforeUpper_4; // @[PMP.scala 113:40]
  wire  _pmpHomogeneous_T_181; // @[PMP.scala 115:21]
  wire  _pmpHomogeneous_T_182; // @[PMP.scala 115:62]
  wire  _pmpHomogeneous_T_183; // @[PMP.scala 115:41]
  wire  _pmpHomogeneous_T_184; // @[PMP.scala 120:58]
  wire  _pmpHomogeneous_T_185; // @[PMP.scala 120:8]
  wire  _pmpHomogeneous_T_186; // @[PMP.scala 140:10]
  wire  _pmpHomogeneous_maskHomogeneous_T_44; // @[package.scala 32:76]
  wire  _pmpHomogeneous_maskHomogeneous_T_46; // @[package.scala 32:76]
  wire  pmpHomogeneous_maskHomogeneous_5; // @[package.scala 32:76]
  wire [31:0] _pmpHomogeneous_T_188; // @[PMP.scala 62:36]
  wire [31:0] _pmpHomogeneous_T_190; // @[PMP.scala 62:48]
  wire [65:0] _GEN_166; // @[PMP.scala 100:53]
  wire [65:0] _pmpHomogeneous_T_192; // @[PMP.scala 100:53]
  wire  _pmpHomogeneous_T_194; // @[PMP.scala 100:78]
  wire  _pmpHomogeneous_T_201; // @[PMP.scala 100:78]
  wire  _pmpHomogeneous_T_208; // @[PMP.scala 100:78]
  wire  _pmpHomogeneous_T_210; // @[package.scala 32:76]
  wire  _pmpHomogeneous_T_212; // @[package.scala 32:76]
  wire  _pmpHomogeneous_T_214; // @[package.scala 32:76]
  wire  _pmpHomogeneous_T_215; // @[PMP.scala 100:21]
  wire  _pmpHomogeneous_beginsAfterUpper_T_29; // @[PMP.scala 109:32]
  wire  pmpHomogeneous_beginsAfterUpper_5; // @[PMP.scala 109:28]
  wire [31:0] _pmpHomogeneous_endsBeforeUpper_T_35; // @[PMP.scala 113:53]
  wire [65:0] _GEN_174; // @[PMP.scala 113:40]
  wire  pmpHomogeneous_endsBeforeUpper_5; // @[PMP.scala 113:40]
  wire  _pmpHomogeneous_T_218; // @[PMP.scala 115:21]
  wire  _pmpHomogeneous_T_219; // @[PMP.scala 115:62]
  wire  _pmpHomogeneous_T_220; // @[PMP.scala 115:41]
  wire  _pmpHomogeneous_T_221; // @[PMP.scala 120:58]
  wire  _pmpHomogeneous_T_222; // @[PMP.scala 120:8]
  wire  _pmpHomogeneous_T_223; // @[PMP.scala 140:10]
  wire  _pmpHomogeneous_maskHomogeneous_T_52; // @[package.scala 32:76]
  wire  _pmpHomogeneous_maskHomogeneous_T_54; // @[package.scala 32:76]
  wire  pmpHomogeneous_maskHomogeneous_6; // @[package.scala 32:76]
  wire [31:0] _pmpHomogeneous_T_225; // @[PMP.scala 62:36]
  wire [31:0] _pmpHomogeneous_T_227; // @[PMP.scala 62:48]
  wire [65:0] _GEN_175; // @[PMP.scala 100:53]
  wire [65:0] _pmpHomogeneous_T_229; // @[PMP.scala 100:53]
  wire  _pmpHomogeneous_T_231; // @[PMP.scala 100:78]
  wire  _pmpHomogeneous_T_238; // @[PMP.scala 100:78]
  wire  _pmpHomogeneous_T_245; // @[PMP.scala 100:78]
  wire  _pmpHomogeneous_T_247; // @[package.scala 32:76]
  wire  _pmpHomogeneous_T_249; // @[package.scala 32:76]
  wire  _pmpHomogeneous_T_251; // @[package.scala 32:76]
  wire  _pmpHomogeneous_T_252; // @[PMP.scala 100:21]
  wire  _pmpHomogeneous_beginsAfterUpper_T_34; // @[PMP.scala 109:32]
  wire  pmpHomogeneous_beginsAfterUpper_6; // @[PMP.scala 109:28]
  wire [31:0] _pmpHomogeneous_endsBeforeUpper_T_41; // @[PMP.scala 113:53]
  wire [65:0] _GEN_183; // @[PMP.scala 113:40]
  wire  pmpHomogeneous_endsBeforeUpper_6; // @[PMP.scala 113:40]
  wire  _pmpHomogeneous_T_255; // @[PMP.scala 115:21]
  wire  _pmpHomogeneous_T_256; // @[PMP.scala 115:62]
  wire  _pmpHomogeneous_T_257; // @[PMP.scala 115:41]
  wire  _pmpHomogeneous_T_258; // @[PMP.scala 120:58]
  wire  _pmpHomogeneous_T_259; // @[PMP.scala 120:8]
  wire  _pmpHomogeneous_T_260; // @[PMP.scala 140:10]
  wire  _pmpHomogeneous_maskHomogeneous_T_60; // @[package.scala 32:76]
  wire  _pmpHomogeneous_maskHomogeneous_T_62; // @[package.scala 32:76]
  wire  pmpHomogeneous_maskHomogeneous_7; // @[package.scala 32:76]
  wire [31:0] _pmpHomogeneous_T_262; // @[PMP.scala 62:36]
  wire [31:0] _pmpHomogeneous_T_264; // @[PMP.scala 62:48]
  wire [65:0] _GEN_184; // @[PMP.scala 100:53]
  wire [65:0] _pmpHomogeneous_T_266; // @[PMP.scala 100:53]
  wire  _pmpHomogeneous_T_268; // @[PMP.scala 100:78]
  wire  _pmpHomogeneous_T_275; // @[PMP.scala 100:78]
  wire  _pmpHomogeneous_T_282; // @[PMP.scala 100:78]
  wire  _pmpHomogeneous_T_284; // @[package.scala 32:76]
  wire  _pmpHomogeneous_T_286; // @[package.scala 32:76]
  wire  _pmpHomogeneous_T_288; // @[package.scala 32:76]
  wire  _pmpHomogeneous_T_289; // @[PMP.scala 100:21]
  wire  _pmpHomogeneous_beginsAfterUpper_T_39; // @[PMP.scala 109:32]
  wire  pmpHomogeneous_beginsAfterUpper_7; // @[PMP.scala 109:28]
  wire [31:0] _pmpHomogeneous_endsBeforeUpper_T_47; // @[PMP.scala 113:53]
  wire [65:0] _GEN_192; // @[PMP.scala 113:40]
  wire  pmpHomogeneous_endsBeforeUpper_7; // @[PMP.scala 113:40]
  wire  _pmpHomogeneous_T_292; // @[PMP.scala 115:21]
  wire  _pmpHomogeneous_T_293; // @[PMP.scala 115:62]
  wire  _pmpHomogeneous_T_294; // @[PMP.scala 115:41]
  wire  _pmpHomogeneous_T_295; // @[PMP.scala 120:58]
  wire  _pmpHomogeneous_T_296; // @[PMP.scala 120:8]
  wire  pmpHomogeneous; // @[PMP.scala 140:10]
  wire  homogeneous; // @[PTW.scala 310:36]
  wire  _T_100; // @[Conditional.scala 37:30]
  wire [2:0] _next_state_T; // @[PTW.scala 332:26]
  wire [2:0] _GEN_40; // @[PTW.scala 331:32]
  wire  _count_T_1; // @[PTW.scala 334:39]
  wire  _T_102; // @[Conditional.scala 37:30]
  wire [1:0] _count_T_3; // @[PTW.scala 338:24]
  wire [2:0] _next_state_T_1; // @[PTW.scala 341:26]
  wire [2:0] _GEN_43; // @[PTW.scala 337:28]
  wire  _T_103; // @[Conditional.scala 37:30]
  wire  _T_104; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_47; // @[PTW.scala 351:35]
  wire  _GEN_48; // @[PTW.scala 351:35]
  wire  _GEN_49; // @[PTW.scala 351:35]
  wire  _T_107; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_54; // @[Conditional.scala 39:67]
  wire  _GEN_55; // @[Conditional.scala 39:67]
  wire  _GEN_56; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_60; // @[Conditional.scala 39:67]
  wire  _GEN_61; // @[Conditional.scala 39:67]
  wire  _GEN_62; // @[Conditional.scala 39:67]
  wire  _GEN_63; // @[Conditional.scala 39:67]
  wire  _GEN_64; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_67; // @[Conditional.scala 39:67]
  wire  _GEN_68; // @[Conditional.scala 39:67]
  wire  _GEN_70; // @[Conditional.scala 39:67]
  wire  _GEN_71; // @[Conditional.scala 39:67]
  wire  _GEN_75; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_76; // @[Conditional.scala 39:67]
  wire  _GEN_77; // @[Conditional.scala 39:67]
  wire  _GEN_79; // @[Conditional.scala 39:67]
  wire  _GEN_80; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_82; // @[Conditional.scala 40:58]
  wire  _GEN_87; // @[Conditional.scala 40:58]
  wire  _GEN_88; // @[Conditional.scala 40:58]
  wire  _r_pte_T_2; // @[PTW.scala 376:15]
  wire  _r_pte_T_4; // @[PTW.scala 376:40]
  wire  _r_pte_T_6; // @[PTW.scala 377:25]
  wire [53:0] pte_2_ppn; // @[PTW.scala 370:13]
  wire [53:0] _r_pte_T_8_ppn; // @[PTW.scala 378:8]
  wire [53:0] pte_1_ppn; // @[PTW.scala 370:13]
  wire [53:0] _r_pte_T_9_ppn; // @[PTW.scala 377:8]
  wire  _r_pte_T_9_d; // @[PTW.scala 377:8]
  wire  _r_pte_T_9_a; // @[PTW.scala 377:8]
  wire  _r_pte_T_9_g; // @[PTW.scala 377:8]
  wire  _r_pte_T_9_u; // @[PTW.scala 377:8]
  wire  _r_pte_T_9_x; // @[PTW.scala 377:8]
  wire  _r_pte_T_9_w; // @[PTW.scala 377:8]
  wire  _r_pte_T_9_r; // @[PTW.scala 377:8]
  wire  _r_pte_T_9_v; // @[PTW.scala 377:8]
  wire [53:0] _r_pte_T_10_ppn; // @[PTW.scala 376:8]
  wire  _r_pte_T_10_d; // @[PTW.scala 376:8]
  wire  _r_pte_T_10_a; // @[PTW.scala 376:8]
  wire  _r_pte_T_10_g; // @[PTW.scala 376:8]
  wire  _r_pte_T_10_u; // @[PTW.scala 376:8]
  wire  _r_pte_T_10_x; // @[PTW.scala 376:8]
  wire  _r_pte_T_10_w; // @[PTW.scala 376:8]
  wire  _r_pte_T_10_r; // @[PTW.scala 376:8]
  wire  _r_pte_T_10_v; // @[PTW.scala 376:8]
  wire  _GEN_90; // @[PTW.scala 384:28]
  wire  _GEN_91; // @[PTW.scala 384:28]
  wire  _T_121; // @[PTW.scala 389:18]
  wire  _T_123; // @[PTW.scala 389:11]
  wire  _l2_refill_T_1; // @[PTW.scala 394:26]
  wire  _l2_refill_T_3; // @[PTW.scala 394:44]
  wire  ae; // @[PTW.scala 395:22]
  wire [2:0] _GEN_102; // @[PTW.scala 390:21]
  wire  _GEN_104; // @[PTW.scala 390:21]
  wire [2:0] _GEN_108; // @[PTW.scala 388:25]
  wire  _T_131; // @[PTW.scala 406:18]
  wire  _T_133; // @[PTW.scala 406:11]
  reg [19:0] PTW_state; // @[Register tracking PTW state]
  reg [31:0] _RAND_39;
  reg  PTW_cov [0:1048575]; // @[Coverage map for PTW]
  reg [31:0] _RAND_40;
  wire  PTW_cov_read_data; // @[Coverage map for PTW]
  wire [19:0] PTW_cov_read_addr; // @[Coverage map for PTW]
  wire  PTW_cov_write_data; // @[Coverage map for PTW]
  wire [19:0] PTW_cov_write_addr; // @[Coverage map for PTW]
  wire  PTW_cov_write_mask; // @[Coverage map for PTW]
  wire  PTW_cov_write_en; // @[Coverage map for PTW]
  reg [29:0] PTW_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_41;
  wire [10:0] valid_shl;
  wire [19:0] valid_pad;
  wire [17:0] count_shl;
  wire [19:0] count_pad;
  wire [8:0] state_reg_shl;
  wire [19:0] state_reg_pad;
  wire [6:0] mem_resp_valid_shl;
  wire [19:0] mem_resp_valid_pad;
  wire [9:0] state_shl;
  wire [19:0] state_pad;
  wire [13:0] invalidated_shl;
  wire [19:0] invalidated_pad;
  wire [19:0] PTW_xor4;
  wire [19:0] PTW_xor1;
  wire [19:0] PTW_xor6;
  wire [19:0] PTW_xor2;
  wire [19:0] PTW_xor0;
  wire [29:0] arb_sum;
  wire [29:0] state_barrier_sum;
  wire [29:0] r_pte_barrier_sum;
  wire  stopEn0;
  wire  stopEn1;
  wire  stopEn2;
  wire  arb_metaAssert_wire;
  wire  state_barrier_metaAssert_wire;
  wire  r_pte_barrier_metaAssert_wire;
  wire  PTW_or4;
  wire  PTW_or1;
  wire  PTW_or6;
  wire  PTW_or2;
  wire  PTW_or0;
  reg  PTW_metaAssert;
  reg [31:0] _RAND_42;
  Arbiter arb ( // @[PTW.scala 112:19]
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_bits_addr(arb_io_in_0_bits_bits_addr),
    .io_in_1_ready(arb_io_in_1_ready),
    .io_in_1_valid(arb_io_in_1_valid),
    .io_in_1_bits_valid(arb_io_in_1_bits_valid),
    .io_in_1_bits_bits_addr(arb_io_in_1_bits_bits_addr),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_valid(arb_io_out_bits_valid),
    .io_out_bits_bits_addr(arb_io_out_bits_bits_addr),
    .io_chosen(arb_io_chosen),
    .io_covSum(arb_io_covSum),
    .metaAssert(arb_metaAssert)
  );
  OptimizationBarrier_42 state_barrier ( // @[package.scala 258:25]
    .io_x(state_barrier_io_x),
    .io_y(state_barrier_io_y),
    .io_covSum(state_barrier_io_covSum),
    .metaAssert(state_barrier_metaAssert)
  );
  OptimizationBarrier_43 r_pte_barrier ( // @[package.scala 258:25]
    .io_x_ppn(r_pte_barrier_io_x_ppn),
    .io_x_d(r_pte_barrier_io_x_d),
    .io_x_a(r_pte_barrier_io_x_a),
    .io_x_g(r_pte_barrier_io_x_g),
    .io_x_u(r_pte_barrier_io_x_u),
    .io_x_x(r_pte_barrier_io_x_x),
    .io_x_w(r_pte_barrier_io_x_w),
    .io_x_r(r_pte_barrier_io_x_r),
    .io_x_v(r_pte_barrier_io_x_v),
    .io_y_ppn(r_pte_barrier_io_y_ppn),
    .io_y_d(r_pte_barrier_io_y_d),
    .io_y_a(r_pte_barrier_io_y_a),
    .io_y_g(r_pte_barrier_io_y_g),
    .io_y_u(r_pte_barrier_io_y_u),
    .io_y_x(r_pte_barrier_io_y_x),
    .io_y_w(r_pte_barrier_io_y_w),
    .io_y_r(r_pte_barrier_io_y_r),
    .io_y_v(r_pte_barrier_io_y_v),
    .io_covSum(r_pte_barrier_io_covSum),
    .metaAssert(r_pte_barrier_metaAssert)
  );
  assign _arb_io_out_ready_T = state == 3'h0; // @[PTW.scala 114:30]
  assign _clock_en_T = state != 3'h0; // @[PTW.scala 118:24]
  assign tmp_v = mem_resp_data[0]; // @[PTW.scala 146:33]
  assign tmp_r = mem_resp_data[1]; // @[PTW.scala 146:33]
  assign tmp_w = mem_resp_data[2]; // @[PTW.scala 146:33]
  assign tmp_x = mem_resp_data[3]; // @[PTW.scala 146:33]
  assign tmp_u = mem_resp_data[4]; // @[PTW.scala 146:33]
  assign tmp_g = mem_resp_data[5]; // @[PTW.scala 146:33]
  assign tmp_a = mem_resp_data[6]; // @[PTW.scala 146:33]
  assign tmp_d = mem_resp_data[7]; // @[PTW.scala 146:33]
  assign tmp_ppn = mem_resp_data[63:10]; // @[PTW.scala 146:33]
  assign _T_11 = tmp_r | tmp_w; // @[PTW.scala 149:17]
  assign _T_12 = _T_11 | tmp_x; // @[PTW.scala 149:26]
  assign _T_13 = count <= 2'h0; // @[PTW.scala 152:21]
  assign _T_15 = tmp_ppn[17:9] != 9'h0; // @[PTW.scala 152:95]
  assign _T_16 = _T_13 & _T_15; // @[PTW.scala 152:26]
  assign _GEN_0 = _T_16 ? 1'h0 : tmp_v; // @[PTW.scala 152:102]
  assign _T_17 = count <= 2'h1; // @[PTW.scala 152:21]
  assign _T_19 = tmp_ppn[8:0] != 9'h0; // @[PTW.scala 152:95]
  assign _T_20 = _T_17 & _T_19; // @[PTW.scala 152:26]
  assign _GEN_1 = _T_20 ? 1'h0 : _GEN_0; // @[PTW.scala 152:102]
  assign res_v = _T_12 ? _GEN_1 : tmp_v; // @[PTW.scala 149:36]
  assign invalid_paddr = tmp_ppn[53:20] != 34'h0; // @[PTW.scala 154:32]
  assign _traverse_T_1 = res_v & ~tmp_r; // @[PTW.scala 72:33]
  assign _traverse_T_3 = _traverse_T_1 & ~tmp_w; // @[PTW.scala 72:39]
  assign _traverse_T_5 = _traverse_T_3 & ~tmp_x; // @[PTW.scala 72:45]
  assign _traverse_T_7 = _traverse_T_5 & ~invalid_paddr; // @[PTW.scala 156:30]
  assign _traverse_T_8 = count < 2'h2; // @[PTW.scala 156:57]
  assign traverse = _traverse_T_7 & _traverse_T_8; // @[PTW.scala 156:48]
  assign vpn_idxs_0 = r_req_addr[26:18]; // @[PTW.scala 158:60]
  assign vpn_idxs_1 = r_req_addr[17:9]; // @[PTW.scala 158:90]
  assign vpn_idxs_2 = r_req_addr[8:0]; // @[PTW.scala 158:90]
  assign _pte_addr_vpn_idx_T = count == 2'h1; // @[package.scala 32:86]
  assign _pte_addr_vpn_idx_T_1 = _pte_addr_vpn_idx_T ? vpn_idxs_1 : vpn_idxs_0; // @[package.scala 32:76]
  assign _pte_addr_vpn_idx_T_2 = count == 2'h2; // @[package.scala 32:86]
  assign _pte_addr_vpn_idx_T_3 = _pte_addr_vpn_idx_T_2 ? vpn_idxs_2 : _pte_addr_vpn_idx_T_1; // @[package.scala 32:76]
  assign _pte_addr_vpn_idx_T_4 = count == 2'h3; // @[package.scala 32:86]
  assign vpn_idx = _pte_addr_vpn_idx_T_4 ? vpn_idxs_2 : _pte_addr_vpn_idx_T_3; // @[package.scala 32:76]
  assign _pte_addr_T = {r_pte_ppn,vpn_idx}; // @[Cat.scala 30:58]
  assign pte_addr = {_pte_addr_T, 3'h0}; // @[PTW.scala 160:29]
  assign fragmented_superpage_ppn_choices_hi = r_pte_ppn[53:18]; // @[PTW.scala 163:69]
  assign fragmented_superpage_ppn_choices_lo = r_req_addr[17:0]; // @[PTW.scala 163:99]
  assign choices_0 = {fragmented_superpage_ppn_choices_hi,fragmented_superpage_ppn_choices_lo}; // @[Cat.scala 30:58]
  assign fragmented_superpage_ppn_choices_hi_1 = r_pte_ppn[53:9]; // @[PTW.scala 163:69]
  assign choices_1 = {fragmented_superpage_ppn_choices_hi_1,vpn_idxs_2}; // @[Cat.scala 30:58]
  assign fragmented_superpage_ppn_truncIdx = count[0]; // @[package.scala 31:49]
  assign fragmented_superpage_ppn = fragmented_superpage_ppn_truncIdx ? choices_1 : choices_0; // @[package.scala 32:76]
  assign _T_22 = arb_io_out_ready & arb_io_out_valid; // @[Decoupled.scala 40:37]
  assign _GEN_115 = {{34'd0}, tags_0}; // @[PTW.scala 179:27]
  assign lo_lo_lo = _GEN_115 == pte_addr; // @[PTW.scala 179:27]
  assign _GEN_116 = {{34'd0}, tags_1}; // @[PTW.scala 179:27]
  assign lo_lo_hi = _GEN_116 == pte_addr; // @[PTW.scala 179:27]
  assign _GEN_117 = {{34'd0}, tags_2}; // @[PTW.scala 179:27]
  assign lo_hi_lo = _GEN_117 == pte_addr; // @[PTW.scala 179:27]
  assign _GEN_118 = {{34'd0}, tags_3}; // @[PTW.scala 179:27]
  assign lo_hi_hi = _GEN_118 == pte_addr; // @[PTW.scala 179:27]
  assign _GEN_119 = {{34'd0}, tags_4}; // @[PTW.scala 179:27]
  assign hi_lo_lo = _GEN_119 == pte_addr; // @[PTW.scala 179:27]
  assign _GEN_120 = {{34'd0}, tags_5}; // @[PTW.scala 179:27]
  assign hi_lo_hi = _GEN_120 == pte_addr; // @[PTW.scala 179:27]
  assign _GEN_121 = {{34'd0}, tags_6}; // @[PTW.scala 179:27]
  assign hi_hi_lo = _GEN_121 == pte_addr; // @[PTW.scala 179:27]
  assign _GEN_122 = {{34'd0}, tags_7}; // @[PTW.scala 179:27]
  assign hi_hi_hi = _GEN_122 == pte_addr; // @[PTW.scala 179:27]
  assign _T_23 = {hi_hi_hi,hi_hi_lo,hi_lo_hi,hi_lo_lo,lo_hi_hi,lo_hi_lo,lo_lo_hi,lo_lo_lo}; // @[Cat.scala 30:58]
  assign hits = _T_23 & valid; // @[PTW.scala 179:48]
  assign hit = |hits; // @[PTW.scala 180:20]
  assign _T_24 = mem_resp_valid & traverse; // @[PTW.scala 181:26]
  assign _T_26 = _T_24 & ~hit; // @[PTW.scala 181:38]
  assign _T_28 = _T_26 & ~invalidated; // @[PTW.scala 181:46]
  assign _T_29 = &valid; // @[PTW.scala 182:25]
  assign hi_1 = state_reg[6]; // @[Replacement.scala 243:38]
  assign left_subtree_state = state_reg[5:3]; // @[package.scala 154:13]
  assign right_subtree_state = state_reg[2:0]; // @[Replacement.scala 245:38]
  assign hi_2 = left_subtree_state[2]; // @[Replacement.scala 243:38]
  assign left_subtree_state_1 = left_subtree_state[1]; // @[package.scala 154:13]
  assign right_subtree_state_1 = left_subtree_state[0]; // @[Replacement.scala 245:38]
  assign lo_1 = hi_2 ? left_subtree_state_1 : right_subtree_state_1; // @[Replacement.scala 250:16]
  assign _T_32 = {hi_2,lo_1}; // @[Cat.scala 30:58]
  assign hi_3 = right_subtree_state[2]; // @[Replacement.scala 243:38]
  assign left_subtree_state_2 = right_subtree_state[1]; // @[package.scala 154:13]
  assign right_subtree_state_2 = right_subtree_state[0]; // @[Replacement.scala 245:38]
  assign lo_2 = hi_3 ? left_subtree_state_2 : right_subtree_state_2; // @[Replacement.scala 250:16]
  assign _T_35 = {hi_3,lo_2}; // @[Cat.scala 30:58]
  assign lo_3 = hi_1 ? _T_32 : _T_35; // @[Replacement.scala 250:16]
  assign _T_36 = {hi_1,lo_3}; // @[Cat.scala 30:58]
  assign _T_38 = ~valid[0]; // @[OneHot.scala 47:40]
  assign _T_39 = ~valid[1]; // @[OneHot.scala 47:40]
  assign _T_40 = ~valid[2]; // @[OneHot.scala 47:40]
  assign _T_41 = ~valid[3]; // @[OneHot.scala 47:40]
  assign _T_42 = ~valid[4]; // @[OneHot.scala 47:40]
  assign _T_43 = ~valid[5]; // @[OneHot.scala 47:40]
  assign _T_44 = ~valid[6]; // @[OneHot.scala 47:40]
  assign _T_46 = _T_44 ? 3'h6 : 3'h7; // @[Mux.scala 47:69]
  assign _T_47 = _T_43 ? 3'h5 : _T_46; // @[Mux.scala 47:69]
  assign _T_48 = _T_42 ? 3'h4 : _T_47; // @[Mux.scala 47:69]
  assign _T_49 = _T_41 ? 3'h3 : _T_48; // @[Mux.scala 47:69]
  assign _T_50 = _T_40 ? 3'h2 : _T_49; // @[Mux.scala 47:69]
  assign _T_51 = _T_39 ? 3'h1 : _T_50; // @[Mux.scala 47:69]
  assign _T_52 = _T_38 ? 3'h0 : _T_51; // @[Mux.scala 47:69]
  assign r = _T_29 ? _T_36 : _T_52; // @[PTW.scala 182:18]
  assign _T_53 = 8'h1 << r; // @[OneHot.scala 58:35]
  assign _T_54 = valid | _T_53; // @[PTW.scala 183:22]
  assign res_ppn = {{34'd0}, tmp_ppn[19:0]}; // @[PTW.scala 148:13]
  assign _T_55 = state == 3'h1; // @[PTW.scala 187:24]
  assign _T_56 = hit & _T_55; // @[PTW.scala 187:15]
  assign hi_4 = hits[7:4]; // @[OneHot.scala 30:18]
  assign lo_4 = hits[3:0]; // @[OneHot.scala 31:18]
  assign hi_5 = |hi_4; // @[OneHot.scala 32:14]
  assign _T_57 = hi_4 | lo_4; // @[OneHot.scala 32:28]
  assign hi_6 = _T_57[3:2]; // @[OneHot.scala 30:18]
  assign lo_5 = _T_57[1:0]; // @[OneHot.scala 31:18]
  assign hi_7 = |hi_6; // @[OneHot.scala 32:14]
  assign _T_58 = hi_6 | lo_5; // @[OneHot.scala 32:28]
  assign lo_6 = _T_58[1]; // @[CircuitMath.scala 30:8]
  assign state_reg_touch_way_sized = {hi_5,hi_7,lo_6}; // @[Cat.scala 30:58]
  assign state_reg_hi_hi = ~state_reg_touch_way_sized[2]; // @[Replacement.scala 196:33]
  assign state_reg_hi_hi_1 = ~state_reg_touch_way_sized[1]; // @[Replacement.scala 196:33]
  assign state_reg_hi_lo = state_reg_hi_hi_1 ? left_subtree_state_1 : ~state_reg_touch_way_sized[0]; // @[Replacement.scala 203:16]
  assign state_reg_lo = state_reg_hi_hi_1 ? ~state_reg_touch_way_sized[0] : right_subtree_state_1; // @[Replacement.scala 206:16]
  assign _state_reg_T_7 = {state_reg_hi_hi_1,state_reg_hi_lo,state_reg_lo}; // @[Cat.scala 30:58]
  assign state_reg_hi_lo_1 = state_reg_hi_hi ? left_subtree_state : _state_reg_T_7; // @[Replacement.scala 203:16]
  assign state_reg_hi_lo_2 = state_reg_hi_hi_1 ? left_subtree_state_2 : ~state_reg_touch_way_sized[0]; // @[Replacement.scala 203:16]
  assign state_reg_lo_1 = state_reg_hi_hi_1 ? ~state_reg_touch_way_sized[0] : right_subtree_state_2; // @[Replacement.scala 206:16]
  assign _state_reg_T_15 = {state_reg_hi_hi_1,state_reg_hi_lo_2,state_reg_lo_1}; // @[Cat.scala 30:58]
  assign state_reg_lo_2 = state_reg_hi_hi ? _state_reg_T_15 : right_subtree_state; // @[Replacement.scala 206:16]
  assign _state_reg_T_16 = {state_reg_hi_hi,state_reg_hi_lo_1,state_reg_lo_2}; // @[Cat.scala 30:58]
  assign _T_61 = io_dpath_sfence_valid & ~io_dpath_sfence_bits_rs1; // @[PTW.scala 188:33]
  assign pte_cache_hit = hit & _traverse_T_8; // @[PTW.scala 193:10]
  assign _T_79 = hits[0] ? data_0 : 20'h0; // @[Mux.scala 27:72]
  assign _T_80 = hits[1] ? data_1 : 20'h0; // @[Mux.scala 27:72]
  assign _T_81 = hits[2] ? data_2 : 20'h0; // @[Mux.scala 27:72]
  assign _T_82 = hits[3] ? data_3 : 20'h0; // @[Mux.scala 27:72]
  assign _T_83 = hits[4] ? data_4 : 20'h0; // @[Mux.scala 27:72]
  assign _T_84 = hits[5] ? data_5 : 20'h0; // @[Mux.scala 27:72]
  assign _T_85 = hits[6] ? data_6 : 20'h0; // @[Mux.scala 27:72]
  assign _T_86 = hits[7] ? data_7 : 20'h0; // @[Mux.scala 27:72]
  assign _T_87 = _T_79 | _T_80; // @[Mux.scala 27:72]
  assign _T_88 = _T_87 | _T_81; // @[Mux.scala 27:72]
  assign _T_89 = _T_88 | _T_82; // @[Mux.scala 27:72]
  assign _T_90 = _T_89 | _T_83; // @[Mux.scala 27:72]
  assign _T_91 = _T_90 | _T_84; // @[Mux.scala 27:72]
  assign _T_92 = _T_91 | _T_85; // @[Mux.scala 27:72]
  assign pte_cache_data = _T_92 | _T_86; // @[Mux.scala 27:72]
  assign _io_dpath_perf_pte_hit_T_1 = pte_hit & _T_55; // @[PTW.scala 197:36]
  assign _T_94 = io_dpath_perf_pte_miss | io_dpath_perf_pte_hit; // @[PTW.scala 198:59]
  assign _T_95 = io_dpath_perf_l2hit & _T_94; // @[PTW.scala 198:32]
  assign _T_98 = ~_T_95 | reset; // @[PTW.scala 198:9]
  assign _invalidated_T_1 = invalidated & _clock_en_T; // @[PTW.scala 285:56]
  assign _io_mem_req_valid_T_1 = state == 3'h3; // @[PTW.scala 287:48]
  assign _pmaPgLevelHomogeneous_T_6 = pte_addr ^ 66'hc000000; // @[Parameters.scala 137:31]
  assign _pmaPgLevelHomogeneous_T_7 = {1'b0,$signed(_pmaPgLevelHomogeneous_T_6)}; // @[Parameters.scala 137:49]
  assign _pmaPgLevelHomogeneous_T_9 = $signed(_pmaPgLevelHomogeneous_T_7) & -67'sh4000000; // @[Parameters.scala 137:52]
  assign _pmaPgLevelHomogeneous_T_10 = $signed(_pmaPgLevelHomogeneous_T_9) == 67'sh0; // @[Parameters.scala 137:67]
  assign _pmaPgLevelHomogeneous_T_11 = pte_addr ^ 66'h60000000; // @[Parameters.scala 137:31]
  assign _pmaPgLevelHomogeneous_T_12 = {1'b0,$signed(_pmaPgLevelHomogeneous_T_11)}; // @[Parameters.scala 137:49]
  assign _pmaPgLevelHomogeneous_T_14 = $signed(_pmaPgLevelHomogeneous_T_12) & -67'sh20000000; // @[Parameters.scala 137:52]
  assign _pmaPgLevelHomogeneous_T_15 = $signed(_pmaPgLevelHomogeneous_T_14) == 67'sh0; // @[Parameters.scala 137:67]
  assign _pmaPgLevelHomogeneous_T_16 = pte_addr ^ 66'h80000000; // @[Parameters.scala 137:31]
  assign _pmaPgLevelHomogeneous_T_17 = {1'b0,$signed(_pmaPgLevelHomogeneous_T_16)}; // @[Parameters.scala 137:49]
  assign _pmaPgLevelHomogeneous_T_19 = $signed(_pmaPgLevelHomogeneous_T_17) & -67'sh10000000; // @[Parameters.scala 137:52]
  assign _pmaPgLevelHomogeneous_T_20 = $signed(_pmaPgLevelHomogeneous_T_19) == 67'sh0; // @[Parameters.scala 137:67]
  assign _pmaPgLevelHomogeneous_T_22 = _pmaPgLevelHomogeneous_T_10 | _pmaPgLevelHomogeneous_T_15; // @[TLBPermissions.scala 99:65]
  assign pmaPgLevelHomogeneous_1 = _pmaPgLevelHomogeneous_T_22 | _pmaPgLevelHomogeneous_T_20; // @[TLBPermissions.scala 99:65]
  assign _pmaPgLevelHomogeneous_T_26 = {1'b0,$signed(pte_addr)}; // @[Parameters.scala 137:49]
  assign _pmaPgLevelHomogeneous_T_53 = $signed(_pmaPgLevelHomogeneous_T_26) & -67'sh1000; // @[Parameters.scala 137:52]
  assign _pmaPgLevelHomogeneous_T_54 = $signed(_pmaPgLevelHomogeneous_T_53) == 67'sh0; // @[Parameters.scala 137:67]
  assign _pmaPgLevelHomogeneous_T_55 = pte_addr ^ 66'h3000; // @[Parameters.scala 137:31]
  assign _pmaPgLevelHomogeneous_T_56 = {1'b0,$signed(_pmaPgLevelHomogeneous_T_55)}; // @[Parameters.scala 137:49]
  assign _pmaPgLevelHomogeneous_T_58 = $signed(_pmaPgLevelHomogeneous_T_56) & -67'sh1000; // @[Parameters.scala 137:52]
  assign _pmaPgLevelHomogeneous_T_59 = $signed(_pmaPgLevelHomogeneous_T_58) == 67'sh0; // @[Parameters.scala 137:67]
  assign _pmaPgLevelHomogeneous_T_60 = pte_addr ^ 66'h10000; // @[Parameters.scala 137:31]
  assign _pmaPgLevelHomogeneous_T_61 = {1'b0,$signed(_pmaPgLevelHomogeneous_T_60)}; // @[Parameters.scala 137:49]
  assign _pmaPgLevelHomogeneous_T_63 = $signed(_pmaPgLevelHomogeneous_T_61) & -67'sh10000; // @[Parameters.scala 137:52]
  assign _pmaPgLevelHomogeneous_T_64 = $signed(_pmaPgLevelHomogeneous_T_63) == 67'sh0; // @[Parameters.scala 137:67]
  assign _pmaPgLevelHomogeneous_T_65 = pte_addr ^ 66'h2000000; // @[Parameters.scala 137:31]
  assign _pmaPgLevelHomogeneous_T_66 = {1'b0,$signed(_pmaPgLevelHomogeneous_T_65)}; // @[Parameters.scala 137:49]
  assign _pmaPgLevelHomogeneous_T_68 = $signed(_pmaPgLevelHomogeneous_T_66) & -67'sh10000; // @[Parameters.scala 137:52]
  assign _pmaPgLevelHomogeneous_T_69 = $signed(_pmaPgLevelHomogeneous_T_68) == 67'sh0; // @[Parameters.scala 137:67]
  assign _pmaPgLevelHomogeneous_T_86 = _pmaPgLevelHomogeneous_T_54 | _pmaPgLevelHomogeneous_T_59; // @[TLBPermissions.scala 99:65]
  assign _pmaPgLevelHomogeneous_T_87 = _pmaPgLevelHomogeneous_T_86 | _pmaPgLevelHomogeneous_T_64; // @[TLBPermissions.scala 99:65]
  assign _pmaPgLevelHomogeneous_T_88 = _pmaPgLevelHomogeneous_T_87 | _pmaPgLevelHomogeneous_T_69; // @[TLBPermissions.scala 99:65]
  assign _pmaPgLevelHomogeneous_T_89 = _pmaPgLevelHomogeneous_T_88 | _pmaPgLevelHomogeneous_T_10; // @[TLBPermissions.scala 99:65]
  assign _pmaPgLevelHomogeneous_T_90 = _pmaPgLevelHomogeneous_T_89 | _pmaPgLevelHomogeneous_T_15; // @[TLBPermissions.scala 99:65]
  assign pmaPgLevelHomogeneous_2 = _pmaPgLevelHomogeneous_T_90 | _pmaPgLevelHomogeneous_T_20; // @[TLBPermissions.scala 99:65]
  assign _pmaHomogeneous_T_1 = _pte_addr_vpn_idx_T & pmaPgLevelHomogeneous_1; // @[package.scala 32:76]
  assign _pmaHomogeneous_T_3 = _pte_addr_vpn_idx_T_2 ? pmaPgLevelHomogeneous_2 : _pmaHomogeneous_T_1; // @[package.scala 32:76]
  assign pmaHomogeneous = _pte_addr_vpn_idx_T_4 ? pmaPgLevelHomogeneous_2 : _pmaHomogeneous_T_3; // @[package.scala 32:76]
  assign _pmpHomogeneous_T_1 = {pte_addr[65:12], 12'h0}; // @[PTW.scala 309:92]
  assign _pmpHomogeneous_maskHomogeneous_T_4 = _pte_addr_vpn_idx_T ? io_dpath_pmp_0_mask[20] : io_dpath_pmp_0_mask[29]; // @[package.scala 32:76]
  assign _pmpHomogeneous_maskHomogeneous_T_6 = _pte_addr_vpn_idx_T_2 ? io_dpath_pmp_0_mask[11] : _pmpHomogeneous_maskHomogeneous_T_4; // @[package.scala 32:76]
  assign pmpHomogeneous_maskHomogeneous = _pte_addr_vpn_idx_T_4 ? io_dpath_pmp_0_mask[11] : _pmpHomogeneous_maskHomogeneous_T_6; // @[package.scala 32:76]
  assign _pmpHomogeneous_T_3 = {io_dpath_pmp_0_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _pmpHomogeneous_T_5 = ~_pmpHomogeneous_T_3 | 32'h3; // @[PMP.scala 62:48]
  assign _GEN_123 = {{34'd0}, ~_pmpHomogeneous_T_5}; // @[PMP.scala 100:53]
  assign _pmpHomogeneous_T_7 = _pmpHomogeneous_T_1 ^ _GEN_123; // @[PMP.scala 100:53]
  assign _pmpHomogeneous_T_9 = _pmpHomogeneous_T_7[65:30] != 36'h0; // @[PMP.scala 100:78]
  assign _pmpHomogeneous_T_16 = _pmpHomogeneous_T_7[65:21] != 45'h0; // @[PMP.scala 100:78]
  assign _pmpHomogeneous_T_23 = _pmpHomogeneous_T_7[65:12] != 54'h0; // @[PMP.scala 100:78]
  assign _pmpHomogeneous_T_25 = _pte_addr_vpn_idx_T ? _pmpHomogeneous_T_16 : _pmpHomogeneous_T_9; // @[package.scala 32:76]
  assign _pmpHomogeneous_T_27 = _pte_addr_vpn_idx_T_2 ? _pmpHomogeneous_T_23 : _pmpHomogeneous_T_25; // @[package.scala 32:76]
  assign _pmpHomogeneous_T_29 = _pte_addr_vpn_idx_T_4 ? _pmpHomogeneous_T_23 : _pmpHomogeneous_T_27; // @[package.scala 32:76]
  assign _pmpHomogeneous_T_30 = pmpHomogeneous_maskHomogeneous | _pmpHomogeneous_T_29; // @[PMP.scala 100:21]
  assign _pmpHomogeneous_beginsAfterUpper_T_4 = _pmpHomogeneous_T_1 < _GEN_123; // @[PMP.scala 109:32]
  assign pmpHomogeneous_beginsAfterUpper = ~_pmpHomogeneous_beginsAfterUpper_T_4; // @[PMP.scala 109:28]
  assign _pmpHomogeneous_pgMask_T_1 = _pte_addr_vpn_idx_T ? 32'hffe00000 : 32'hc0000000; // @[package.scala 32:76]
  assign _pmpHomogeneous_pgMask_T_3 = _pte_addr_vpn_idx_T_2 ? 32'hfffff000 : _pmpHomogeneous_pgMask_T_1; // @[package.scala 32:76]
  assign pmpHomogeneous_pgMask = _pte_addr_vpn_idx_T_4 ? 32'hfffff000 : _pmpHomogeneous_pgMask_T_3; // @[package.scala 32:76]
  assign _GEN_127 = {{34'd0}, pmpHomogeneous_pgMask}; // @[PMP.scala 112:30]
  assign _pmpHomogeneous_endsBeforeLower_T = _pmpHomogeneous_T_1 & _GEN_127; // @[PMP.scala 112:30]
  assign _pmpHomogeneous_endsBeforeUpper_T_5 = ~_pmpHomogeneous_T_5 & pmpHomogeneous_pgMask; // @[PMP.scala 113:53]
  assign _GEN_129 = {{34'd0}, _pmpHomogeneous_endsBeforeUpper_T_5}; // @[PMP.scala 113:40]
  assign pmpHomogeneous_endsBeforeUpper = _pmpHomogeneous_endsBeforeLower_T < _GEN_129; // @[PMP.scala 113:40]
  assign _pmpHomogeneous_T_35 = pmpHomogeneous_beginsAfterUpper | pmpHomogeneous_endsBeforeUpper; // @[PMP.scala 115:41]
  assign _pmpHomogeneous_T_36 = ~io_dpath_pmp_0_cfg_a[0] | _pmpHomogeneous_T_35; // @[PMP.scala 120:58]
  assign _pmpHomogeneous_T_37 = io_dpath_pmp_0_cfg_a[1] ? _pmpHomogeneous_T_30 : _pmpHomogeneous_T_36; // @[PMP.scala 120:8]
  assign _pmpHomogeneous_maskHomogeneous_T_12 = _pte_addr_vpn_idx_T ? io_dpath_pmp_1_mask[20] : io_dpath_pmp_1_mask[29]; // @[package.scala 32:76]
  assign _pmpHomogeneous_maskHomogeneous_T_14 = _pte_addr_vpn_idx_T_2 ? io_dpath_pmp_1_mask[11] : _pmpHomogeneous_maskHomogeneous_T_12; // @[package.scala 32:76]
  assign pmpHomogeneous_maskHomogeneous_1 = _pte_addr_vpn_idx_T_4 ? io_dpath_pmp_1_mask[11] : _pmpHomogeneous_maskHomogeneous_T_14; // @[package.scala 32:76]
  assign _pmpHomogeneous_T_40 = {io_dpath_pmp_1_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _pmpHomogeneous_T_42 = ~_pmpHomogeneous_T_40 | 32'h3; // @[PMP.scala 62:48]
  assign _GEN_130 = {{34'd0}, ~_pmpHomogeneous_T_42}; // @[PMP.scala 100:53]
  assign _pmpHomogeneous_T_44 = _pmpHomogeneous_T_1 ^ _GEN_130; // @[PMP.scala 100:53]
  assign _pmpHomogeneous_T_46 = _pmpHomogeneous_T_44[65:30] != 36'h0; // @[PMP.scala 100:78]
  assign _pmpHomogeneous_T_53 = _pmpHomogeneous_T_44[65:21] != 45'h0; // @[PMP.scala 100:78]
  assign _pmpHomogeneous_T_60 = _pmpHomogeneous_T_44[65:12] != 54'h0; // @[PMP.scala 100:78]
  assign _pmpHomogeneous_T_62 = _pte_addr_vpn_idx_T ? _pmpHomogeneous_T_53 : _pmpHomogeneous_T_46; // @[package.scala 32:76]
  assign _pmpHomogeneous_T_64 = _pte_addr_vpn_idx_T_2 ? _pmpHomogeneous_T_60 : _pmpHomogeneous_T_62; // @[package.scala 32:76]
  assign _pmpHomogeneous_T_66 = _pte_addr_vpn_idx_T_4 ? _pmpHomogeneous_T_60 : _pmpHomogeneous_T_64; // @[package.scala 32:76]
  assign _pmpHomogeneous_T_67 = pmpHomogeneous_maskHomogeneous_1 | _pmpHomogeneous_T_66; // @[PMP.scala 100:21]
  assign _pmpHomogeneous_beginsAfterUpper_T_9 = _pmpHomogeneous_T_1 < _GEN_130; // @[PMP.scala 109:32]
  assign pmpHomogeneous_beginsAfterUpper_1 = ~_pmpHomogeneous_beginsAfterUpper_T_9; // @[PMP.scala 109:28]
  assign _pmpHomogeneous_endsBeforeUpper_T_11 = ~_pmpHomogeneous_T_42 & pmpHomogeneous_pgMask; // @[PMP.scala 113:53]
  assign _GEN_138 = {{34'd0}, _pmpHomogeneous_endsBeforeUpper_T_11}; // @[PMP.scala 113:40]
  assign pmpHomogeneous_endsBeforeUpper_1 = _pmpHomogeneous_endsBeforeLower_T < _GEN_138; // @[PMP.scala 113:40]
  assign _pmpHomogeneous_T_70 = pmpHomogeneous_endsBeforeUpper | pmpHomogeneous_beginsAfterUpper_1; // @[PMP.scala 115:21]
  assign _pmpHomogeneous_T_71 = pmpHomogeneous_beginsAfterUpper & pmpHomogeneous_endsBeforeUpper_1; // @[PMP.scala 115:62]
  assign _pmpHomogeneous_T_72 = _pmpHomogeneous_T_70 | _pmpHomogeneous_T_71; // @[PMP.scala 115:41]
  assign _pmpHomogeneous_T_73 = ~io_dpath_pmp_1_cfg_a[0] | _pmpHomogeneous_T_72; // @[PMP.scala 120:58]
  assign _pmpHomogeneous_T_74 = io_dpath_pmp_1_cfg_a[1] ? _pmpHomogeneous_T_67 : _pmpHomogeneous_T_73; // @[PMP.scala 120:8]
  assign _pmpHomogeneous_T_75 = _pmpHomogeneous_T_37 & _pmpHomogeneous_T_74; // @[PMP.scala 140:10]
  assign _pmpHomogeneous_maskHomogeneous_T_20 = _pte_addr_vpn_idx_T ? io_dpath_pmp_2_mask[20] : io_dpath_pmp_2_mask[29]; // @[package.scala 32:76]
  assign _pmpHomogeneous_maskHomogeneous_T_22 = _pte_addr_vpn_idx_T_2 ? io_dpath_pmp_2_mask[11] : _pmpHomogeneous_maskHomogeneous_T_20; // @[package.scala 32:76]
  assign pmpHomogeneous_maskHomogeneous_2 = _pte_addr_vpn_idx_T_4 ? io_dpath_pmp_2_mask[11] : _pmpHomogeneous_maskHomogeneous_T_22; // @[package.scala 32:76]
  assign _pmpHomogeneous_T_77 = {io_dpath_pmp_2_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _pmpHomogeneous_T_79 = ~_pmpHomogeneous_T_77 | 32'h3; // @[PMP.scala 62:48]
  assign _GEN_139 = {{34'd0}, ~_pmpHomogeneous_T_79}; // @[PMP.scala 100:53]
  assign _pmpHomogeneous_T_81 = _pmpHomogeneous_T_1 ^ _GEN_139; // @[PMP.scala 100:53]
  assign _pmpHomogeneous_T_83 = _pmpHomogeneous_T_81[65:30] != 36'h0; // @[PMP.scala 100:78]
  assign _pmpHomogeneous_T_90 = _pmpHomogeneous_T_81[65:21] != 45'h0; // @[PMP.scala 100:78]
  assign _pmpHomogeneous_T_97 = _pmpHomogeneous_T_81[65:12] != 54'h0; // @[PMP.scala 100:78]
  assign _pmpHomogeneous_T_99 = _pte_addr_vpn_idx_T ? _pmpHomogeneous_T_90 : _pmpHomogeneous_T_83; // @[package.scala 32:76]
  assign _pmpHomogeneous_T_101 = _pte_addr_vpn_idx_T_2 ? _pmpHomogeneous_T_97 : _pmpHomogeneous_T_99; // @[package.scala 32:76]
  assign _pmpHomogeneous_T_103 = _pte_addr_vpn_idx_T_4 ? _pmpHomogeneous_T_97 : _pmpHomogeneous_T_101; // @[package.scala 32:76]
  assign _pmpHomogeneous_T_104 = pmpHomogeneous_maskHomogeneous_2 | _pmpHomogeneous_T_103; // @[PMP.scala 100:21]
  assign _pmpHomogeneous_beginsAfterUpper_T_14 = _pmpHomogeneous_T_1 < _GEN_139; // @[PMP.scala 109:32]
  assign pmpHomogeneous_beginsAfterUpper_2 = ~_pmpHomogeneous_beginsAfterUpper_T_14; // @[PMP.scala 109:28]
  assign _pmpHomogeneous_endsBeforeUpper_T_17 = ~_pmpHomogeneous_T_79 & pmpHomogeneous_pgMask; // @[PMP.scala 113:53]
  assign _GEN_147 = {{34'd0}, _pmpHomogeneous_endsBeforeUpper_T_17}; // @[PMP.scala 113:40]
  assign pmpHomogeneous_endsBeforeUpper_2 = _pmpHomogeneous_endsBeforeLower_T < _GEN_147; // @[PMP.scala 113:40]
  assign _pmpHomogeneous_T_107 = pmpHomogeneous_endsBeforeUpper_1 | pmpHomogeneous_beginsAfterUpper_2; // @[PMP.scala 115:21]
  assign _pmpHomogeneous_T_108 = pmpHomogeneous_beginsAfterUpper_1 & pmpHomogeneous_endsBeforeUpper_2; // @[PMP.scala 115:62]
  assign _pmpHomogeneous_T_109 = _pmpHomogeneous_T_107 | _pmpHomogeneous_T_108; // @[PMP.scala 115:41]
  assign _pmpHomogeneous_T_110 = ~io_dpath_pmp_2_cfg_a[0] | _pmpHomogeneous_T_109; // @[PMP.scala 120:58]
  assign _pmpHomogeneous_T_111 = io_dpath_pmp_2_cfg_a[1] ? _pmpHomogeneous_T_104 : _pmpHomogeneous_T_110; // @[PMP.scala 120:8]
  assign _pmpHomogeneous_T_112 = _pmpHomogeneous_T_75 & _pmpHomogeneous_T_111; // @[PMP.scala 140:10]
  assign _pmpHomogeneous_maskHomogeneous_T_28 = _pte_addr_vpn_idx_T ? io_dpath_pmp_3_mask[20] : io_dpath_pmp_3_mask[29]; // @[package.scala 32:76]
  assign _pmpHomogeneous_maskHomogeneous_T_30 = _pte_addr_vpn_idx_T_2 ? io_dpath_pmp_3_mask[11] : _pmpHomogeneous_maskHomogeneous_T_28; // @[package.scala 32:76]
  assign pmpHomogeneous_maskHomogeneous_3 = _pte_addr_vpn_idx_T_4 ? io_dpath_pmp_3_mask[11] : _pmpHomogeneous_maskHomogeneous_T_30; // @[package.scala 32:76]
  assign _pmpHomogeneous_T_114 = {io_dpath_pmp_3_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _pmpHomogeneous_T_116 = ~_pmpHomogeneous_T_114 | 32'h3; // @[PMP.scala 62:48]
  assign _GEN_148 = {{34'd0}, ~_pmpHomogeneous_T_116}; // @[PMP.scala 100:53]
  assign _pmpHomogeneous_T_118 = _pmpHomogeneous_T_1 ^ _GEN_148; // @[PMP.scala 100:53]
  assign _pmpHomogeneous_T_120 = _pmpHomogeneous_T_118[65:30] != 36'h0; // @[PMP.scala 100:78]
  assign _pmpHomogeneous_T_127 = _pmpHomogeneous_T_118[65:21] != 45'h0; // @[PMP.scala 100:78]
  assign _pmpHomogeneous_T_134 = _pmpHomogeneous_T_118[65:12] != 54'h0; // @[PMP.scala 100:78]
  assign _pmpHomogeneous_T_136 = _pte_addr_vpn_idx_T ? _pmpHomogeneous_T_127 : _pmpHomogeneous_T_120; // @[package.scala 32:76]
  assign _pmpHomogeneous_T_138 = _pte_addr_vpn_idx_T_2 ? _pmpHomogeneous_T_134 : _pmpHomogeneous_T_136; // @[package.scala 32:76]
  assign _pmpHomogeneous_T_140 = _pte_addr_vpn_idx_T_4 ? _pmpHomogeneous_T_134 : _pmpHomogeneous_T_138; // @[package.scala 32:76]
  assign _pmpHomogeneous_T_141 = pmpHomogeneous_maskHomogeneous_3 | _pmpHomogeneous_T_140; // @[PMP.scala 100:21]
  assign _pmpHomogeneous_beginsAfterUpper_T_19 = _pmpHomogeneous_T_1 < _GEN_148; // @[PMP.scala 109:32]
  assign pmpHomogeneous_beginsAfterUpper_3 = ~_pmpHomogeneous_beginsAfterUpper_T_19; // @[PMP.scala 109:28]
  assign _pmpHomogeneous_endsBeforeUpper_T_23 = ~_pmpHomogeneous_T_116 & pmpHomogeneous_pgMask; // @[PMP.scala 113:53]
  assign _GEN_156 = {{34'd0}, _pmpHomogeneous_endsBeforeUpper_T_23}; // @[PMP.scala 113:40]
  assign pmpHomogeneous_endsBeforeUpper_3 = _pmpHomogeneous_endsBeforeLower_T < _GEN_156; // @[PMP.scala 113:40]
  assign _pmpHomogeneous_T_144 = pmpHomogeneous_endsBeforeUpper_2 | pmpHomogeneous_beginsAfterUpper_3; // @[PMP.scala 115:21]
  assign _pmpHomogeneous_T_145 = pmpHomogeneous_beginsAfterUpper_2 & pmpHomogeneous_endsBeforeUpper_3; // @[PMP.scala 115:62]
  assign _pmpHomogeneous_T_146 = _pmpHomogeneous_T_144 | _pmpHomogeneous_T_145; // @[PMP.scala 115:41]
  assign _pmpHomogeneous_T_147 = ~io_dpath_pmp_3_cfg_a[0] | _pmpHomogeneous_T_146; // @[PMP.scala 120:58]
  assign _pmpHomogeneous_T_148 = io_dpath_pmp_3_cfg_a[1] ? _pmpHomogeneous_T_141 : _pmpHomogeneous_T_147; // @[PMP.scala 120:8]
  assign _pmpHomogeneous_T_149 = _pmpHomogeneous_T_112 & _pmpHomogeneous_T_148; // @[PMP.scala 140:10]
  assign _pmpHomogeneous_maskHomogeneous_T_36 = _pte_addr_vpn_idx_T ? io_dpath_pmp_4_mask[20] : io_dpath_pmp_4_mask[29]; // @[package.scala 32:76]
  assign _pmpHomogeneous_maskHomogeneous_T_38 = _pte_addr_vpn_idx_T_2 ? io_dpath_pmp_4_mask[11] : _pmpHomogeneous_maskHomogeneous_T_36; // @[package.scala 32:76]
  assign pmpHomogeneous_maskHomogeneous_4 = _pte_addr_vpn_idx_T_4 ? io_dpath_pmp_4_mask[11] : _pmpHomogeneous_maskHomogeneous_T_38; // @[package.scala 32:76]
  assign _pmpHomogeneous_T_151 = {io_dpath_pmp_4_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _pmpHomogeneous_T_153 = ~_pmpHomogeneous_T_151 | 32'h3; // @[PMP.scala 62:48]
  assign _GEN_157 = {{34'd0}, ~_pmpHomogeneous_T_153}; // @[PMP.scala 100:53]
  assign _pmpHomogeneous_T_155 = _pmpHomogeneous_T_1 ^ _GEN_157; // @[PMP.scala 100:53]
  assign _pmpHomogeneous_T_157 = _pmpHomogeneous_T_155[65:30] != 36'h0; // @[PMP.scala 100:78]
  assign _pmpHomogeneous_T_164 = _pmpHomogeneous_T_155[65:21] != 45'h0; // @[PMP.scala 100:78]
  assign _pmpHomogeneous_T_171 = _pmpHomogeneous_T_155[65:12] != 54'h0; // @[PMP.scala 100:78]
  assign _pmpHomogeneous_T_173 = _pte_addr_vpn_idx_T ? _pmpHomogeneous_T_164 : _pmpHomogeneous_T_157; // @[package.scala 32:76]
  assign _pmpHomogeneous_T_175 = _pte_addr_vpn_idx_T_2 ? _pmpHomogeneous_T_171 : _pmpHomogeneous_T_173; // @[package.scala 32:76]
  assign _pmpHomogeneous_T_177 = _pte_addr_vpn_idx_T_4 ? _pmpHomogeneous_T_171 : _pmpHomogeneous_T_175; // @[package.scala 32:76]
  assign _pmpHomogeneous_T_178 = pmpHomogeneous_maskHomogeneous_4 | _pmpHomogeneous_T_177; // @[PMP.scala 100:21]
  assign _pmpHomogeneous_beginsAfterUpper_T_24 = _pmpHomogeneous_T_1 < _GEN_157; // @[PMP.scala 109:32]
  assign pmpHomogeneous_beginsAfterUpper_4 = ~_pmpHomogeneous_beginsAfterUpper_T_24; // @[PMP.scala 109:28]
  assign _pmpHomogeneous_endsBeforeUpper_T_29 = ~_pmpHomogeneous_T_153 & pmpHomogeneous_pgMask; // @[PMP.scala 113:53]
  assign _GEN_165 = {{34'd0}, _pmpHomogeneous_endsBeforeUpper_T_29}; // @[PMP.scala 113:40]
  assign pmpHomogeneous_endsBeforeUpper_4 = _pmpHomogeneous_endsBeforeLower_T < _GEN_165; // @[PMP.scala 113:40]
  assign _pmpHomogeneous_T_181 = pmpHomogeneous_endsBeforeUpper_3 | pmpHomogeneous_beginsAfterUpper_4; // @[PMP.scala 115:21]
  assign _pmpHomogeneous_T_182 = pmpHomogeneous_beginsAfterUpper_3 & pmpHomogeneous_endsBeforeUpper_4; // @[PMP.scala 115:62]
  assign _pmpHomogeneous_T_183 = _pmpHomogeneous_T_181 | _pmpHomogeneous_T_182; // @[PMP.scala 115:41]
  assign _pmpHomogeneous_T_184 = ~io_dpath_pmp_4_cfg_a[0] | _pmpHomogeneous_T_183; // @[PMP.scala 120:58]
  assign _pmpHomogeneous_T_185 = io_dpath_pmp_4_cfg_a[1] ? _pmpHomogeneous_T_178 : _pmpHomogeneous_T_184; // @[PMP.scala 120:8]
  assign _pmpHomogeneous_T_186 = _pmpHomogeneous_T_149 & _pmpHomogeneous_T_185; // @[PMP.scala 140:10]
  assign _pmpHomogeneous_maskHomogeneous_T_44 = _pte_addr_vpn_idx_T ? io_dpath_pmp_5_mask[20] : io_dpath_pmp_5_mask[29]; // @[package.scala 32:76]
  assign _pmpHomogeneous_maskHomogeneous_T_46 = _pte_addr_vpn_idx_T_2 ? io_dpath_pmp_5_mask[11] : _pmpHomogeneous_maskHomogeneous_T_44; // @[package.scala 32:76]
  assign pmpHomogeneous_maskHomogeneous_5 = _pte_addr_vpn_idx_T_4 ? io_dpath_pmp_5_mask[11] : _pmpHomogeneous_maskHomogeneous_T_46; // @[package.scala 32:76]
  assign _pmpHomogeneous_T_188 = {io_dpath_pmp_5_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _pmpHomogeneous_T_190 = ~_pmpHomogeneous_T_188 | 32'h3; // @[PMP.scala 62:48]
  assign _GEN_166 = {{34'd0}, ~_pmpHomogeneous_T_190}; // @[PMP.scala 100:53]
  assign _pmpHomogeneous_T_192 = _pmpHomogeneous_T_1 ^ _GEN_166; // @[PMP.scala 100:53]
  assign _pmpHomogeneous_T_194 = _pmpHomogeneous_T_192[65:30] != 36'h0; // @[PMP.scala 100:78]
  assign _pmpHomogeneous_T_201 = _pmpHomogeneous_T_192[65:21] != 45'h0; // @[PMP.scala 100:78]
  assign _pmpHomogeneous_T_208 = _pmpHomogeneous_T_192[65:12] != 54'h0; // @[PMP.scala 100:78]
  assign _pmpHomogeneous_T_210 = _pte_addr_vpn_idx_T ? _pmpHomogeneous_T_201 : _pmpHomogeneous_T_194; // @[package.scala 32:76]
  assign _pmpHomogeneous_T_212 = _pte_addr_vpn_idx_T_2 ? _pmpHomogeneous_T_208 : _pmpHomogeneous_T_210; // @[package.scala 32:76]
  assign _pmpHomogeneous_T_214 = _pte_addr_vpn_idx_T_4 ? _pmpHomogeneous_T_208 : _pmpHomogeneous_T_212; // @[package.scala 32:76]
  assign _pmpHomogeneous_T_215 = pmpHomogeneous_maskHomogeneous_5 | _pmpHomogeneous_T_214; // @[PMP.scala 100:21]
  assign _pmpHomogeneous_beginsAfterUpper_T_29 = _pmpHomogeneous_T_1 < _GEN_166; // @[PMP.scala 109:32]
  assign pmpHomogeneous_beginsAfterUpper_5 = ~_pmpHomogeneous_beginsAfterUpper_T_29; // @[PMP.scala 109:28]
  assign _pmpHomogeneous_endsBeforeUpper_T_35 = ~_pmpHomogeneous_T_190 & pmpHomogeneous_pgMask; // @[PMP.scala 113:53]
  assign _GEN_174 = {{34'd0}, _pmpHomogeneous_endsBeforeUpper_T_35}; // @[PMP.scala 113:40]
  assign pmpHomogeneous_endsBeforeUpper_5 = _pmpHomogeneous_endsBeforeLower_T < _GEN_174; // @[PMP.scala 113:40]
  assign _pmpHomogeneous_T_218 = pmpHomogeneous_endsBeforeUpper_4 | pmpHomogeneous_beginsAfterUpper_5; // @[PMP.scala 115:21]
  assign _pmpHomogeneous_T_219 = pmpHomogeneous_beginsAfterUpper_4 & pmpHomogeneous_endsBeforeUpper_5; // @[PMP.scala 115:62]
  assign _pmpHomogeneous_T_220 = _pmpHomogeneous_T_218 | _pmpHomogeneous_T_219; // @[PMP.scala 115:41]
  assign _pmpHomogeneous_T_221 = ~io_dpath_pmp_5_cfg_a[0] | _pmpHomogeneous_T_220; // @[PMP.scala 120:58]
  assign _pmpHomogeneous_T_222 = io_dpath_pmp_5_cfg_a[1] ? _pmpHomogeneous_T_215 : _pmpHomogeneous_T_221; // @[PMP.scala 120:8]
  assign _pmpHomogeneous_T_223 = _pmpHomogeneous_T_186 & _pmpHomogeneous_T_222; // @[PMP.scala 140:10]
  assign _pmpHomogeneous_maskHomogeneous_T_52 = _pte_addr_vpn_idx_T ? io_dpath_pmp_6_mask[20] : io_dpath_pmp_6_mask[29]; // @[package.scala 32:76]
  assign _pmpHomogeneous_maskHomogeneous_T_54 = _pte_addr_vpn_idx_T_2 ? io_dpath_pmp_6_mask[11] : _pmpHomogeneous_maskHomogeneous_T_52; // @[package.scala 32:76]
  assign pmpHomogeneous_maskHomogeneous_6 = _pte_addr_vpn_idx_T_4 ? io_dpath_pmp_6_mask[11] : _pmpHomogeneous_maskHomogeneous_T_54; // @[package.scala 32:76]
  assign _pmpHomogeneous_T_225 = {io_dpath_pmp_6_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _pmpHomogeneous_T_227 = ~_pmpHomogeneous_T_225 | 32'h3; // @[PMP.scala 62:48]
  assign _GEN_175 = {{34'd0}, ~_pmpHomogeneous_T_227}; // @[PMP.scala 100:53]
  assign _pmpHomogeneous_T_229 = _pmpHomogeneous_T_1 ^ _GEN_175; // @[PMP.scala 100:53]
  assign _pmpHomogeneous_T_231 = _pmpHomogeneous_T_229[65:30] != 36'h0; // @[PMP.scala 100:78]
  assign _pmpHomogeneous_T_238 = _pmpHomogeneous_T_229[65:21] != 45'h0; // @[PMP.scala 100:78]
  assign _pmpHomogeneous_T_245 = _pmpHomogeneous_T_229[65:12] != 54'h0; // @[PMP.scala 100:78]
  assign _pmpHomogeneous_T_247 = _pte_addr_vpn_idx_T ? _pmpHomogeneous_T_238 : _pmpHomogeneous_T_231; // @[package.scala 32:76]
  assign _pmpHomogeneous_T_249 = _pte_addr_vpn_idx_T_2 ? _pmpHomogeneous_T_245 : _pmpHomogeneous_T_247; // @[package.scala 32:76]
  assign _pmpHomogeneous_T_251 = _pte_addr_vpn_idx_T_4 ? _pmpHomogeneous_T_245 : _pmpHomogeneous_T_249; // @[package.scala 32:76]
  assign _pmpHomogeneous_T_252 = pmpHomogeneous_maskHomogeneous_6 | _pmpHomogeneous_T_251; // @[PMP.scala 100:21]
  assign _pmpHomogeneous_beginsAfterUpper_T_34 = _pmpHomogeneous_T_1 < _GEN_175; // @[PMP.scala 109:32]
  assign pmpHomogeneous_beginsAfterUpper_6 = ~_pmpHomogeneous_beginsAfterUpper_T_34; // @[PMP.scala 109:28]
  assign _pmpHomogeneous_endsBeforeUpper_T_41 = ~_pmpHomogeneous_T_227 & pmpHomogeneous_pgMask; // @[PMP.scala 113:53]
  assign _GEN_183 = {{34'd0}, _pmpHomogeneous_endsBeforeUpper_T_41}; // @[PMP.scala 113:40]
  assign pmpHomogeneous_endsBeforeUpper_6 = _pmpHomogeneous_endsBeforeLower_T < _GEN_183; // @[PMP.scala 113:40]
  assign _pmpHomogeneous_T_255 = pmpHomogeneous_endsBeforeUpper_5 | pmpHomogeneous_beginsAfterUpper_6; // @[PMP.scala 115:21]
  assign _pmpHomogeneous_T_256 = pmpHomogeneous_beginsAfterUpper_5 & pmpHomogeneous_endsBeforeUpper_6; // @[PMP.scala 115:62]
  assign _pmpHomogeneous_T_257 = _pmpHomogeneous_T_255 | _pmpHomogeneous_T_256; // @[PMP.scala 115:41]
  assign _pmpHomogeneous_T_258 = ~io_dpath_pmp_6_cfg_a[0] | _pmpHomogeneous_T_257; // @[PMP.scala 120:58]
  assign _pmpHomogeneous_T_259 = io_dpath_pmp_6_cfg_a[1] ? _pmpHomogeneous_T_252 : _pmpHomogeneous_T_258; // @[PMP.scala 120:8]
  assign _pmpHomogeneous_T_260 = _pmpHomogeneous_T_223 & _pmpHomogeneous_T_259; // @[PMP.scala 140:10]
  assign _pmpHomogeneous_maskHomogeneous_T_60 = _pte_addr_vpn_idx_T ? io_dpath_pmp_7_mask[20] : io_dpath_pmp_7_mask[29]; // @[package.scala 32:76]
  assign _pmpHomogeneous_maskHomogeneous_T_62 = _pte_addr_vpn_idx_T_2 ? io_dpath_pmp_7_mask[11] : _pmpHomogeneous_maskHomogeneous_T_60; // @[package.scala 32:76]
  assign pmpHomogeneous_maskHomogeneous_7 = _pte_addr_vpn_idx_T_4 ? io_dpath_pmp_7_mask[11] : _pmpHomogeneous_maskHomogeneous_T_62; // @[package.scala 32:76]
  assign _pmpHomogeneous_T_262 = {io_dpath_pmp_7_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _pmpHomogeneous_T_264 = ~_pmpHomogeneous_T_262 | 32'h3; // @[PMP.scala 62:48]
  assign _GEN_184 = {{34'd0}, ~_pmpHomogeneous_T_264}; // @[PMP.scala 100:53]
  assign _pmpHomogeneous_T_266 = _pmpHomogeneous_T_1 ^ _GEN_184; // @[PMP.scala 100:53]
  assign _pmpHomogeneous_T_268 = _pmpHomogeneous_T_266[65:30] != 36'h0; // @[PMP.scala 100:78]
  assign _pmpHomogeneous_T_275 = _pmpHomogeneous_T_266[65:21] != 45'h0; // @[PMP.scala 100:78]
  assign _pmpHomogeneous_T_282 = _pmpHomogeneous_T_266[65:12] != 54'h0; // @[PMP.scala 100:78]
  assign _pmpHomogeneous_T_284 = _pte_addr_vpn_idx_T ? _pmpHomogeneous_T_275 : _pmpHomogeneous_T_268; // @[package.scala 32:76]
  assign _pmpHomogeneous_T_286 = _pte_addr_vpn_idx_T_2 ? _pmpHomogeneous_T_282 : _pmpHomogeneous_T_284; // @[package.scala 32:76]
  assign _pmpHomogeneous_T_288 = _pte_addr_vpn_idx_T_4 ? _pmpHomogeneous_T_282 : _pmpHomogeneous_T_286; // @[package.scala 32:76]
  assign _pmpHomogeneous_T_289 = pmpHomogeneous_maskHomogeneous_7 | _pmpHomogeneous_T_288; // @[PMP.scala 100:21]
  assign _pmpHomogeneous_beginsAfterUpper_T_39 = _pmpHomogeneous_T_1 < _GEN_184; // @[PMP.scala 109:32]
  assign pmpHomogeneous_beginsAfterUpper_7 = ~_pmpHomogeneous_beginsAfterUpper_T_39; // @[PMP.scala 109:28]
  assign _pmpHomogeneous_endsBeforeUpper_T_47 = ~_pmpHomogeneous_T_264 & pmpHomogeneous_pgMask; // @[PMP.scala 113:53]
  assign _GEN_192 = {{34'd0}, _pmpHomogeneous_endsBeforeUpper_T_47}; // @[PMP.scala 113:40]
  assign pmpHomogeneous_endsBeforeUpper_7 = _pmpHomogeneous_endsBeforeLower_T < _GEN_192; // @[PMP.scala 113:40]
  assign _pmpHomogeneous_T_292 = pmpHomogeneous_endsBeforeUpper_6 | pmpHomogeneous_beginsAfterUpper_7; // @[PMP.scala 115:21]
  assign _pmpHomogeneous_T_293 = pmpHomogeneous_beginsAfterUpper_6 & pmpHomogeneous_endsBeforeUpper_7; // @[PMP.scala 115:62]
  assign _pmpHomogeneous_T_294 = _pmpHomogeneous_T_292 | _pmpHomogeneous_T_293; // @[PMP.scala 115:41]
  assign _pmpHomogeneous_T_295 = ~io_dpath_pmp_7_cfg_a[0] | _pmpHomogeneous_T_294; // @[PMP.scala 120:58]
  assign _pmpHomogeneous_T_296 = io_dpath_pmp_7_cfg_a[1] ? _pmpHomogeneous_T_289 : _pmpHomogeneous_T_295; // @[PMP.scala 120:8]
  assign pmpHomogeneous = _pmpHomogeneous_T_260 & _pmpHomogeneous_T_296; // @[PMP.scala 140:10]
  assign homogeneous = pmaHomogeneous & pmpHomogeneous; // @[PTW.scala 310:36]
  assign _T_100 = 3'h0 == state; // @[Conditional.scala 37:30]
  assign _next_state_T = arb_io_out_bits_valid ? 3'h1 : 3'h0; // @[PTW.scala 332:26]
  assign _GEN_40 = _T_22 ? _next_state_T : state; // @[PTW.scala 331:32]
  assign _count_T_1 = 1'h0 - 1'h0; // @[PTW.scala 334:39]
  assign _T_102 = 3'h1 == state; // @[Conditional.scala 37:30]
  assign _count_T_3 = count + 2'h1; // @[PTW.scala 338:24]
  assign _next_state_T_1 = io_mem_req_ready ? 3'h2 : 3'h1; // @[PTW.scala 341:26]
  assign _GEN_43 = pte_cache_hit ? state : _next_state_T_1; // @[PTW.scala 337:28]
  assign _T_103 = 3'h2 == state; // @[Conditional.scala 37:30]
  assign _T_104 = 3'h4 == state; // @[Conditional.scala 37:30]
  assign _GEN_47 = io_mem_s2_xcpt_ae_ld ? 3'h0 : 3'h5; // @[PTW.scala 351:35]
  assign _GEN_48 = io_mem_s2_xcpt_ae_ld & ~r_req_dest; // @[PTW.scala 351:35]
  assign _GEN_49 = io_mem_s2_xcpt_ae_ld & r_req_dest; // @[PTW.scala 351:35]
  assign _T_107 = 3'h7 == state; // @[Conditional.scala 37:30]
  assign _GEN_54 = _T_107 ? 3'h0 : state; // @[Conditional.scala 39:67]
  assign _GEN_55 = _T_107 & ~r_req_dest; // @[Conditional.scala 39:67]
  assign _GEN_56 = _T_107 & r_req_dest; // @[Conditional.scala 39:67]
  assign _GEN_60 = _T_104 ? _GEN_47 : _GEN_54; // @[Conditional.scala 39:67]
  assign _GEN_61 = _T_104 & _traverse_T_8; // @[Conditional.scala 39:67]
  assign _GEN_62 = _T_104 & io_mem_s2_xcpt_ae_ld; // @[Conditional.scala 39:67]
  assign _GEN_63 = _T_104 ? _GEN_48 : _GEN_55; // @[Conditional.scala 39:67]
  assign _GEN_64 = _T_104 ? _GEN_49 : _GEN_56; // @[Conditional.scala 39:67]
  assign _GEN_67 = _T_103 ? 3'h4 : _GEN_60; // @[Conditional.scala 39:67]
  assign _GEN_68 = _T_103 ? 1'h0 : _GEN_61; // @[Conditional.scala 39:67]
  assign _GEN_70 = _T_103 ? 1'h0 : _GEN_63; // @[Conditional.scala 39:67]
  assign _GEN_71 = _T_103 ? 1'h0 : _GEN_64; // @[Conditional.scala 39:67]
  assign _GEN_75 = _T_102 & pte_cache_hit; // @[Conditional.scala 39:67]
  assign _GEN_76 = _T_102 ? _GEN_43 : _GEN_67; // @[Conditional.scala 39:67]
  assign _GEN_77 = _T_102 ? 1'h0 : _GEN_68; // @[Conditional.scala 39:67]
  assign _GEN_79 = _T_102 ? 1'h0 : _GEN_70; // @[Conditional.scala 39:67]
  assign _GEN_80 = _T_102 ? 1'h0 : _GEN_71; // @[Conditional.scala 39:67]
  assign _GEN_82 = _T_100 ? _GEN_40 : _GEN_76; // @[Conditional.scala 40:58]
  assign _GEN_87 = _T_100 ? 1'h0 : _GEN_79; // @[Conditional.scala 40:58]
  assign _GEN_88 = _T_100 ? 1'h0 : _GEN_80; // @[Conditional.scala 40:58]
  assign _r_pte_T_2 = state == 3'h7; // @[PTW.scala 376:15]
  assign _r_pte_T_4 = _r_pte_T_2 & ~homogeneous; // @[PTW.scala 376:40]
  assign _r_pte_T_6 = _T_55 & pte_cache_hit; // @[PTW.scala 377:25]
  assign pte_2_ppn = {{10'd0}, io_dpath_ptbr_ppn}; // @[PTW.scala 370:13]
  assign _r_pte_T_8_ppn = _T_22 ? pte_2_ppn : r_pte_ppn; // @[PTW.scala 378:8]
  assign pte_1_ppn = {{34'd0}, pte_cache_data}; // @[PTW.scala 370:13]
  assign _r_pte_T_9_ppn = _r_pte_T_6 ? pte_1_ppn : _r_pte_T_8_ppn; // @[PTW.scala 377:8]
  assign _r_pte_T_9_d = _r_pte_T_6 ? 1'h0 : r_pte_d; // @[PTW.scala 377:8]
  assign _r_pte_T_9_a = _r_pte_T_6 ? 1'h0 : r_pte_a; // @[PTW.scala 377:8]
  assign _r_pte_T_9_g = _r_pte_T_6 ? 1'h0 : r_pte_g; // @[PTW.scala 377:8]
  assign _r_pte_T_9_u = _r_pte_T_6 ? 1'h0 : r_pte_u; // @[PTW.scala 377:8]
  assign _r_pte_T_9_x = _r_pte_T_6 ? 1'h0 : r_pte_x; // @[PTW.scala 377:8]
  assign _r_pte_T_9_w = _r_pte_T_6 ? 1'h0 : r_pte_w; // @[PTW.scala 377:8]
  assign _r_pte_T_9_r = _r_pte_T_6 ? 1'h0 : r_pte_r; // @[PTW.scala 377:8]
  assign _r_pte_T_9_v = _r_pte_T_6 ? 1'h0 : r_pte_v; // @[PTW.scala 377:8]
  assign _r_pte_T_10_ppn = _r_pte_T_4 ? fragmented_superpage_ppn : _r_pte_T_9_ppn; // @[PTW.scala 376:8]
  assign _r_pte_T_10_d = _r_pte_T_4 ? r_pte_d : _r_pte_T_9_d; // @[PTW.scala 376:8]
  assign _r_pte_T_10_a = _r_pte_T_4 ? r_pte_a : _r_pte_T_9_a; // @[PTW.scala 376:8]
  assign _r_pte_T_10_g = _r_pte_T_4 ? r_pte_g : _r_pte_T_9_g; // @[PTW.scala 376:8]
  assign _r_pte_T_10_u = _r_pte_T_4 ? r_pte_u : _r_pte_T_9_u; // @[PTW.scala 376:8]
  assign _r_pte_T_10_x = _r_pte_T_4 ? r_pte_x : _r_pte_T_9_x; // @[PTW.scala 376:8]
  assign _r_pte_T_10_w = _r_pte_T_4 ? r_pte_w : _r_pte_T_9_w; // @[PTW.scala 376:8]
  assign _r_pte_T_10_r = _r_pte_T_4 ? r_pte_r : _r_pte_T_9_r; // @[PTW.scala 376:8]
  assign _r_pte_T_10_v = _r_pte_T_4 ? r_pte_v : _r_pte_T_9_v; // @[PTW.scala 376:8]
  assign _GEN_90 = ~r_req_dest | _GEN_87; // @[PTW.scala 384:28]
  assign _GEN_91 = r_req_dest | _GEN_88; // @[PTW.scala 384:28]
  assign _T_121 = state == 3'h5; // @[PTW.scala 389:18]
  assign _T_123 = _T_121 | reset; // @[PTW.scala 389:11]
  assign _l2_refill_T_1 = res_v & ~invalid_paddr; // @[PTW.scala 394:26]
  assign _l2_refill_T_3 = _l2_refill_T_1 & _pte_addr_vpn_idx_T_2; // @[PTW.scala 394:44]
  assign ae = res_v & invalid_paddr; // @[PTW.scala 395:22]
  assign _GEN_102 = traverse ? 3'h1 : 3'h0; // @[PTW.scala 390:21]
  assign _GEN_104 = traverse ? 1'h0 : _l2_refill_T_3; // @[PTW.scala 390:21]
  assign _GEN_108 = mem_resp_valid ? _GEN_102 : _GEN_82; // @[PTW.scala 388:25]
  assign _T_131 = state == 3'h4; // @[PTW.scala 406:18]
  assign _T_133 = _T_131 | reset; // @[PTW.scala 406:11]
  assign io_requestor_0_req_ready = arb_io_in_0_ready; // @[PTW.scala 113:13]
  assign io_requestor_0_resp_valid = resp_valid_0; // @[PTW.scala 313:32]
  assign io_requestor_0_resp_bits_ae = resp_ae; // @[PTW.scala 314:34]
  assign io_requestor_0_resp_bits_pte_ppn = r_pte_ppn; // @[PTW.scala 315:35]
  assign io_requestor_0_resp_bits_pte_d = r_pte_d; // @[PTW.scala 315:35]
  assign io_requestor_0_resp_bits_pte_a = r_pte_a; // @[PTW.scala 315:35]
  assign io_requestor_0_resp_bits_pte_g = r_pte_g; // @[PTW.scala 315:35]
  assign io_requestor_0_resp_bits_pte_u = r_pte_u; // @[PTW.scala 315:35]
  assign io_requestor_0_resp_bits_pte_x = r_pte_x; // @[PTW.scala 315:35]
  assign io_requestor_0_resp_bits_pte_w = r_pte_w; // @[PTW.scala 315:35]
  assign io_requestor_0_resp_bits_pte_r = r_pte_r; // @[PTW.scala 315:35]
  assign io_requestor_0_resp_bits_pte_v = r_pte_v; // @[PTW.scala 315:35]
  assign io_requestor_0_resp_bits_level = count; // @[PTW.scala 316:37]
  assign io_requestor_0_resp_bits_homogeneous = pmaHomogeneous & pmpHomogeneous; // @[PTW.scala 317:43]
  assign io_requestor_0_ptbr_mode = io_dpath_ptbr_mode; // @[PTW.scala 319:26]
  assign io_requestor_0_status_debug = io_dpath_status_debug; // @[PTW.scala 321:28]
  assign io_requestor_0_status_dprv = io_dpath_status_dprv; // @[PTW.scala 321:28]
  assign io_requestor_0_status_mxr = io_dpath_status_mxr; // @[PTW.scala 321:28]
  assign io_requestor_0_status_sum = io_dpath_status_sum; // @[PTW.scala 321:28]
  assign io_requestor_0_pmp_0_cfg_l = io_dpath_pmp_0_cfg_l; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_0_cfg_a = io_dpath_pmp_0_cfg_a; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_0_cfg_x = io_dpath_pmp_0_cfg_x; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_0_cfg_w = io_dpath_pmp_0_cfg_w; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_0_cfg_r = io_dpath_pmp_0_cfg_r; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_0_addr = io_dpath_pmp_0_addr; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_0_mask = io_dpath_pmp_0_mask; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_1_cfg_l = io_dpath_pmp_1_cfg_l; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_1_cfg_a = io_dpath_pmp_1_cfg_a; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_1_cfg_x = io_dpath_pmp_1_cfg_x; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_1_cfg_w = io_dpath_pmp_1_cfg_w; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_1_cfg_r = io_dpath_pmp_1_cfg_r; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_1_addr = io_dpath_pmp_1_addr; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_1_mask = io_dpath_pmp_1_mask; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_2_cfg_l = io_dpath_pmp_2_cfg_l; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_2_cfg_a = io_dpath_pmp_2_cfg_a; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_2_cfg_x = io_dpath_pmp_2_cfg_x; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_2_cfg_w = io_dpath_pmp_2_cfg_w; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_2_cfg_r = io_dpath_pmp_2_cfg_r; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_2_addr = io_dpath_pmp_2_addr; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_2_mask = io_dpath_pmp_2_mask; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_3_cfg_l = io_dpath_pmp_3_cfg_l; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_3_cfg_a = io_dpath_pmp_3_cfg_a; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_3_cfg_x = io_dpath_pmp_3_cfg_x; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_3_cfg_w = io_dpath_pmp_3_cfg_w; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_3_cfg_r = io_dpath_pmp_3_cfg_r; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_3_addr = io_dpath_pmp_3_addr; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_3_mask = io_dpath_pmp_3_mask; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_4_cfg_l = io_dpath_pmp_4_cfg_l; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_4_cfg_a = io_dpath_pmp_4_cfg_a; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_4_cfg_x = io_dpath_pmp_4_cfg_x; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_4_cfg_w = io_dpath_pmp_4_cfg_w; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_4_cfg_r = io_dpath_pmp_4_cfg_r; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_4_addr = io_dpath_pmp_4_addr; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_4_mask = io_dpath_pmp_4_mask; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_5_cfg_l = io_dpath_pmp_5_cfg_l; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_5_cfg_a = io_dpath_pmp_5_cfg_a; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_5_cfg_x = io_dpath_pmp_5_cfg_x; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_5_cfg_w = io_dpath_pmp_5_cfg_w; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_5_cfg_r = io_dpath_pmp_5_cfg_r; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_5_addr = io_dpath_pmp_5_addr; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_5_mask = io_dpath_pmp_5_mask; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_6_cfg_l = io_dpath_pmp_6_cfg_l; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_6_cfg_a = io_dpath_pmp_6_cfg_a; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_6_cfg_x = io_dpath_pmp_6_cfg_x; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_6_cfg_w = io_dpath_pmp_6_cfg_w; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_6_cfg_r = io_dpath_pmp_6_cfg_r; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_6_addr = io_dpath_pmp_6_addr; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_6_mask = io_dpath_pmp_6_mask; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_7_cfg_l = io_dpath_pmp_7_cfg_l; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_7_cfg_a = io_dpath_pmp_7_cfg_a; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_7_cfg_x = io_dpath_pmp_7_cfg_x; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_7_cfg_w = io_dpath_pmp_7_cfg_w; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_7_cfg_r = io_dpath_pmp_7_cfg_r; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_7_addr = io_dpath_pmp_7_addr; // @[PTW.scala 322:25]
  assign io_requestor_0_pmp_7_mask = io_dpath_pmp_7_mask; // @[PTW.scala 322:25]
  assign io_requestor_1_req_ready = arb_io_in_1_ready; // @[PTW.scala 113:13]
  assign io_requestor_1_resp_valid = resp_valid_1; // @[PTW.scala 313:32]
  assign io_requestor_1_resp_bits_ae = resp_ae; // @[PTW.scala 314:34]
  assign io_requestor_1_resp_bits_pte_ppn = r_pte_ppn; // @[PTW.scala 315:35]
  assign io_requestor_1_resp_bits_pte_d = r_pte_d; // @[PTW.scala 315:35]
  assign io_requestor_1_resp_bits_pte_a = r_pte_a; // @[PTW.scala 315:35]
  assign io_requestor_1_resp_bits_pte_g = r_pte_g; // @[PTW.scala 315:35]
  assign io_requestor_1_resp_bits_pte_u = r_pte_u; // @[PTW.scala 315:35]
  assign io_requestor_1_resp_bits_pte_x = r_pte_x; // @[PTW.scala 315:35]
  assign io_requestor_1_resp_bits_pte_w = r_pte_w; // @[PTW.scala 315:35]
  assign io_requestor_1_resp_bits_pte_r = r_pte_r; // @[PTW.scala 315:35]
  assign io_requestor_1_resp_bits_pte_v = r_pte_v; // @[PTW.scala 315:35]
  assign io_requestor_1_resp_bits_level = count; // @[PTW.scala 316:37]
  assign io_requestor_1_resp_bits_homogeneous = pmaHomogeneous & pmpHomogeneous; // @[PTW.scala 317:43]
  assign io_requestor_1_ptbr_mode = io_dpath_ptbr_mode; // @[PTW.scala 319:26]
  assign io_requestor_1_status_debug = io_dpath_status_debug; // @[PTW.scala 321:28]
  assign io_requestor_1_status_prv = io_dpath_status_prv; // @[PTW.scala 321:28]
  assign io_requestor_1_pmp_0_cfg_l = io_dpath_pmp_0_cfg_l; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_0_cfg_a = io_dpath_pmp_0_cfg_a; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_0_cfg_x = io_dpath_pmp_0_cfg_x; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_0_cfg_w = io_dpath_pmp_0_cfg_w; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_0_cfg_r = io_dpath_pmp_0_cfg_r; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_0_addr = io_dpath_pmp_0_addr; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_0_mask = io_dpath_pmp_0_mask; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_1_cfg_l = io_dpath_pmp_1_cfg_l; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_1_cfg_a = io_dpath_pmp_1_cfg_a; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_1_cfg_x = io_dpath_pmp_1_cfg_x; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_1_cfg_w = io_dpath_pmp_1_cfg_w; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_1_cfg_r = io_dpath_pmp_1_cfg_r; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_1_addr = io_dpath_pmp_1_addr; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_1_mask = io_dpath_pmp_1_mask; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_2_cfg_l = io_dpath_pmp_2_cfg_l; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_2_cfg_a = io_dpath_pmp_2_cfg_a; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_2_cfg_x = io_dpath_pmp_2_cfg_x; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_2_cfg_w = io_dpath_pmp_2_cfg_w; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_2_cfg_r = io_dpath_pmp_2_cfg_r; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_2_addr = io_dpath_pmp_2_addr; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_2_mask = io_dpath_pmp_2_mask; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_3_cfg_l = io_dpath_pmp_3_cfg_l; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_3_cfg_a = io_dpath_pmp_3_cfg_a; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_3_cfg_x = io_dpath_pmp_3_cfg_x; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_3_cfg_w = io_dpath_pmp_3_cfg_w; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_3_cfg_r = io_dpath_pmp_3_cfg_r; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_3_addr = io_dpath_pmp_3_addr; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_3_mask = io_dpath_pmp_3_mask; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_4_cfg_l = io_dpath_pmp_4_cfg_l; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_4_cfg_a = io_dpath_pmp_4_cfg_a; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_4_cfg_x = io_dpath_pmp_4_cfg_x; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_4_cfg_w = io_dpath_pmp_4_cfg_w; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_4_cfg_r = io_dpath_pmp_4_cfg_r; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_4_addr = io_dpath_pmp_4_addr; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_4_mask = io_dpath_pmp_4_mask; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_5_cfg_l = io_dpath_pmp_5_cfg_l; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_5_cfg_a = io_dpath_pmp_5_cfg_a; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_5_cfg_x = io_dpath_pmp_5_cfg_x; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_5_cfg_w = io_dpath_pmp_5_cfg_w; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_5_cfg_r = io_dpath_pmp_5_cfg_r; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_5_addr = io_dpath_pmp_5_addr; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_5_mask = io_dpath_pmp_5_mask; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_6_cfg_l = io_dpath_pmp_6_cfg_l; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_6_cfg_a = io_dpath_pmp_6_cfg_a; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_6_cfg_x = io_dpath_pmp_6_cfg_x; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_6_cfg_w = io_dpath_pmp_6_cfg_w; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_6_cfg_r = io_dpath_pmp_6_cfg_r; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_6_addr = io_dpath_pmp_6_addr; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_6_mask = io_dpath_pmp_6_mask; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_7_cfg_l = io_dpath_pmp_7_cfg_l; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_7_cfg_a = io_dpath_pmp_7_cfg_a; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_7_cfg_x = io_dpath_pmp_7_cfg_x; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_7_cfg_w = io_dpath_pmp_7_cfg_w; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_7_cfg_r = io_dpath_pmp_7_cfg_r; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_7_addr = io_dpath_pmp_7_addr; // @[PTW.scala 322:25]
  assign io_requestor_1_pmp_7_mask = io_dpath_pmp_7_mask; // @[PTW.scala 322:25]
  assign io_requestor_1_customCSRs_csrs_0_value = io_dpath_customCSRs_csrs_0_value; // @[PTW.scala 320:32]
  assign io_mem_req_valid = _T_55 | _io_mem_req_valid_T_1; // @[PTW.scala 287:20]
  assign io_mem_req_bits_addr = pte_addr[39:0]; // @[PTW.scala 292:24]
  assign io_mem_s1_kill = state != 3'h2; // @[PTW.scala 295:18]
  assign io_dpath_perf_l2hit = 1'h0; // @[PTW.scala 204:23]
  assign io_dpath_perf_pte_miss = _T_100 ? 1'h0 : _GEN_77; // @[PTW.scala 196:26 PTW.scala 350:30]
  assign io_dpath_perf_pte_hit = _io_dpath_perf_pte_hit_T_1 & ~io_dpath_perf_l2hit; // @[PTW.scala 197:25]
  assign arb_io_in_0_valid = io_requestor_0_req_valid; // @[PTW.scala 113:13]
  assign arb_io_in_0_bits_bits_addr = io_requestor_0_req_bits_bits_addr; // @[PTW.scala 113:13]
  assign arb_io_in_1_valid = io_requestor_1_req_valid; // @[PTW.scala 113:13]
  assign arb_io_in_1_bits_valid = io_requestor_1_req_bits_valid; // @[PTW.scala 113:13]
  assign arb_io_in_1_bits_bits_addr = io_requestor_1_req_bits_bits_addr; // @[PTW.scala 113:13]
  assign arb_io_out_ready = _arb_io_out_ready_T & ~l2_refill; // @[PTW.scala 114:20]
  assign state_barrier_io_x = io_mem_s2_nack ? 3'h1 : _GEN_108; // @[package.scala 266:18]
  assign r_pte_barrier_io_x_ppn = mem_resp_valid ? res_ppn : _r_pte_T_10_ppn; // @[package.scala 266:18]
  assign r_pte_barrier_io_x_d = mem_resp_valid ? tmp_d : _r_pte_T_10_d; // @[package.scala 266:18]
  assign r_pte_barrier_io_x_a = mem_resp_valid ? tmp_a : _r_pte_T_10_a; // @[package.scala 266:18]
  assign r_pte_barrier_io_x_g = mem_resp_valid ? tmp_g : _r_pte_T_10_g; // @[package.scala 266:18]
  assign r_pte_barrier_io_x_u = mem_resp_valid ? tmp_u : _r_pte_T_10_u; // @[package.scala 266:18]
  assign r_pte_barrier_io_x_x = mem_resp_valid ? tmp_x : _r_pte_T_10_x; // @[package.scala 266:18]
  assign r_pte_barrier_io_x_w = mem_resp_valid ? tmp_w : _r_pte_T_10_w; // @[package.scala 266:18]
  assign r_pte_barrier_io_x_r = mem_resp_valid ? tmp_r : _r_pte_T_10_r; // @[package.scala 266:18]
  assign r_pte_barrier_io_x_v = mem_resp_valid ? res_v : _r_pte_T_10_v; // @[package.scala 266:18]
  assign PTW_cov_read_addr = PTW_state;
  assign PTW_cov_read_data = PTW_cov[PTW_cov_read_addr]; // @[Coverage map for PTW]
  assign PTW_cov_write_data = 1'h1;
  assign PTW_cov_write_addr = PTW_state;
  assign PTW_cov_write_mask = 1'h1;
  assign PTW_cov_write_en = 1'h1;
  assign valid_shl = {valid, 3'h0};
  assign valid_pad = {9'h0,valid_shl};
  assign count_shl = {count, 16'h0};
  assign count_pad = {2'h0,count_shl};
  assign state_reg_shl = {state_reg, 2'h0};
  assign state_reg_pad = {11'h0,state_reg_shl};
  assign mem_resp_valid_shl = {mem_resp_valid, 6'h0};
  assign mem_resp_valid_pad = {13'h0,mem_resp_valid_shl};
  assign state_shl = {state, 7'h0};
  assign state_pad = {10'h0,state_shl};
  assign invalidated_shl = {invalidated, 13'h0};
  assign invalidated_pad = {6'h0,invalidated_shl};
  assign PTW_xor4 = count_pad ^ state_reg_pad;
  assign PTW_xor1 = valid_pad ^ PTW_xor4;
  assign PTW_xor6 = state_pad ^ invalidated_pad;
  assign PTW_xor2 = mem_resp_valid_pad ^ PTW_xor6;
  assign PTW_xor0 = PTW_xor1 ^ PTW_xor2;
  assign arb_sum = PTW_covSum + arb_io_covSum;
  assign state_barrier_sum = arb_sum + state_barrier_io_covSum;
  assign r_pte_barrier_sum = state_barrier_sum + r_pte_barrier_io_covSum;
  assign io_covSum = r_pte_barrier_sum;
  assign stopEn0 = ~_T_98;
  assign stopEn1 = mem_resp_valid & ~_T_123;
  assign stopEn2 = io_mem_s2_nack & ~_T_133;
  assign arb_metaAssert_wire = arb_metaAssert;
  assign state_barrier_metaAssert_wire = state_barrier_metaAssert;
  assign r_pte_barrier_metaAssert_wire = r_pte_barrier_metaAssert;
  assign PTW_or4 = stopEn1 | stopEn2;
  assign PTW_or1 = stopEn0 | PTW_or4;
  assign PTW_or6 = state_barrier_metaAssert_wire | r_pte_barrier_metaAssert_wire;
  assign PTW_or2 = arb_metaAssert_wire | PTW_or6;
  assign PTW_or0 = PTW_or1 | PTW_or2;
  assign metaAssert = PTW_metaAssert;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  l2_refill = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  resp_valid_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  resp_valid_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  invalidated = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  count = _RAND_5[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  resp_ae = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  r_req_addr = _RAND_7[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  r_req_dest = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {2{`RANDOM}};
  r_pte_ppn = _RAND_9[53:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  r_pte_d = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  r_pte_a = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  r_pte_g = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  r_pte_u = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  r_pte_x = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  r_pte_w = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  r_pte_r = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  r_pte_v = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  mem_resp_valid = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {2{`RANDOM}};
  mem_resp_data = _RAND_19[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  state_reg = _RAND_20[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  valid = _RAND_21[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  tags_0 = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  tags_1 = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  tags_2 = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  tags_3 = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  tags_4 = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  tags_5 = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  tags_6 = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  tags_7 = _RAND_29[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  data_0 = _RAND_30[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  data_1 = _RAND_31[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  data_2 = _RAND_32[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  data_3 = _RAND_33[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  data_4 = _RAND_34[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  data_5 = _RAND_35[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  data_6 = _RAND_36[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  data_7 = _RAND_37[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  pte_hit = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  PTW_state = _RAND_39[19:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1048576; initvar = initvar+1)
    PTW_cov[initvar] = _RAND_40[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  PTW_covSum = _RAND_41[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  PTW_metaAssert = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      state <= 3'h0;
    end else if (reset) begin
      state <= 3'h0;
    end else begin
      state <= state_barrier_io_y;
    end
    if (metaReset) begin
      l2_refill <= 1'h0;
    end else begin
      l2_refill <= mem_resp_valid & _GEN_104;
    end
    if (metaReset) begin
      resp_valid_0 <= 1'h0;
    end else if (mem_resp_valid) begin
      if (traverse) begin
        if (_T_100) begin
          resp_valid_0 <= 1'h0;
        end else if (_T_102) begin
          resp_valid_0 <= 1'h0;
        end else if (_T_103) begin
          resp_valid_0 <= 1'h0;
        end else if (_T_104) begin
          resp_valid_0 <= _GEN_48;
        end else begin
          resp_valid_0 <= _GEN_55;
        end
      end else begin
        resp_valid_0 <= _GEN_90;
      end
    end else if (_T_100) begin
      resp_valid_0 <= 1'h0;
    end else if (_T_102) begin
      resp_valid_0 <= 1'h0;
    end else if (_T_103) begin
      resp_valid_0 <= 1'h0;
    end else if (_T_104) begin
      resp_valid_0 <= _GEN_48;
    end else begin
      resp_valid_0 <= _GEN_55;
    end
    if (metaReset) begin
      resp_valid_1 <= 1'h0;
    end else if (mem_resp_valid) begin
      if (traverse) begin
        if (_T_100) begin
          resp_valid_1 <= 1'h0;
        end else if (_T_102) begin
          resp_valid_1 <= 1'h0;
        end else if (_T_103) begin
          resp_valid_1 <= 1'h0;
        end else if (_T_104) begin
          resp_valid_1 <= _GEN_49;
        end else begin
          resp_valid_1 <= _GEN_56;
        end
      end else begin
        resp_valid_1 <= _GEN_91;
      end
    end else if (_T_100) begin
      resp_valid_1 <= 1'h0;
    end else if (_T_102) begin
      resp_valid_1 <= 1'h0;
    end else if (_T_103) begin
      resp_valid_1 <= 1'h0;
    end else if (_T_104) begin
      resp_valid_1 <= _GEN_49;
    end else begin
      resp_valid_1 <= _GEN_56;
    end
    if (metaReset) begin
      invalidated <= 1'h0;
    end else begin
      invalidated <= io_dpath_sfence_valid | _invalidated_T_1;
    end
    if (metaReset) begin
      count <= 2'h0;
    end else if (mem_resp_valid) begin
      if (traverse) begin
        count <= _count_T_3;
      end else if (_T_100) begin
        count <= {{1'd0}, _count_T_1};
      end else if (_T_102) begin
        if (pte_cache_hit) begin
          count <= _count_T_3;
        end
      end else if (!(_T_103)) begin
        if (!(_T_104)) begin
          if (_T_107) begin
            if (~homogeneous) begin
              count <= 2'h2;
            end
          end
        end
      end
    end else if (_T_100) begin
      count <= {{1'd0}, _count_T_1};
    end else if (_T_102) begin
      if (pte_cache_hit) begin
        count <= _count_T_3;
      end
    end else if (!(_T_103)) begin
      if (!(_T_104)) begin
        if (_T_107) begin
          if (~homogeneous) begin
            count <= 2'h2;
          end
        end
      end
    end
    if (metaReset) begin
      resp_ae <= 1'h0;
    end else if (mem_resp_valid) begin
      if (traverse) begin
        if (_T_100) begin
          resp_ae <= 1'h0;
        end else if (_T_102) begin
          resp_ae <= 1'h0;
        end else if (_T_103) begin
          resp_ae <= 1'h0;
        end else begin
          resp_ae <= _GEN_62;
        end
      end else begin
        resp_ae <= ae;
      end
    end else if (_T_100) begin
      resp_ae <= 1'h0;
    end else if (_T_102) begin
      resp_ae <= 1'h0;
    end else if (_T_103) begin
      resp_ae <= 1'h0;
    end else begin
      resp_ae <= _GEN_62;
    end
    if (metaReset) begin
      r_req_addr <= 27'h0;
    end else if (_T_22) begin
      r_req_addr <= arb_io_out_bits_bits_addr;
    end
    if (metaReset) begin
      r_req_dest <= 1'h0;
    end else if (_T_22) begin
      r_req_dest <= arb_io_chosen;
    end
    if (metaReset) begin
      r_pte_ppn <= 54'h0;
    end else begin
      r_pte_ppn <= r_pte_barrier_io_y_ppn;
    end
    if (metaReset) begin
      r_pte_d <= 1'h0;
    end else begin
      r_pte_d <= r_pte_barrier_io_y_d;
    end
    if (metaReset) begin
      r_pte_a <= 1'h0;
    end else begin
      r_pte_a <= r_pte_barrier_io_y_a;
    end
    if (metaReset) begin
      r_pte_g <= 1'h0;
    end else begin
      r_pte_g <= r_pte_barrier_io_y_g;
    end
    if (metaReset) begin
      r_pte_u <= 1'h0;
    end else begin
      r_pte_u <= r_pte_barrier_io_y_u;
    end
    if (metaReset) begin
      r_pte_x <= 1'h0;
    end else begin
      r_pte_x <= r_pte_barrier_io_y_x;
    end
    if (metaReset) begin
      r_pte_w <= 1'h0;
    end else begin
      r_pte_w <= r_pte_barrier_io_y_w;
    end
    if (metaReset) begin
      r_pte_r <= 1'h0;
    end else begin
      r_pte_r <= r_pte_barrier_io_y_r;
    end
    if (metaReset) begin
      r_pte_v <= 1'h0;
    end else begin
      r_pte_v <= r_pte_barrier_io_y_v;
    end
    if (metaReset) begin
      mem_resp_valid <= 1'h0;
    end else begin
      mem_resp_valid <= io_mem_resp_valid;
    end
    if (metaReset) begin
      mem_resp_data <= 64'h0;
    end else begin
      mem_resp_data <= io_mem_resp_bits_data;
    end
    if (metaReset) begin
      state_reg <= 7'h0;
    end else if (reset) begin
      state_reg <= 7'h0;
    end else if (_T_56) begin
      state_reg <= _state_reg_T_16;
    end
    if (metaReset) begin
      valid <= 8'h0;
    end else if (reset) begin
      valid <= 8'h0;
    end else if (_T_61) begin
      valid <= 8'h0;
    end else if (_T_28) begin
      valid <= _T_54;
    end
    if (metaReset) begin
      tags_0 <= 32'h0;
    end else if (_T_28) begin
      if (3'h0 == r) begin
        tags_0 <= pte_addr[31:0];
      end
    end
    if (metaReset) begin
      tags_1 <= 32'h0;
    end else if (_T_28) begin
      if (3'h1 == r) begin
        tags_1 <= pte_addr[31:0];
      end
    end
    if (metaReset) begin
      tags_2 <= 32'h0;
    end else if (_T_28) begin
      if (3'h2 == r) begin
        tags_2 <= pte_addr[31:0];
      end
    end
    if (metaReset) begin
      tags_3 <= 32'h0;
    end else if (_T_28) begin
      if (3'h3 == r) begin
        tags_3 <= pte_addr[31:0];
      end
    end
    if (metaReset) begin
      tags_4 <= 32'h0;
    end else if (_T_28) begin
      if (3'h4 == r) begin
        tags_4 <= pte_addr[31:0];
      end
    end
    if (metaReset) begin
      tags_5 <= 32'h0;
    end else if (_T_28) begin
      if (3'h5 == r) begin
        tags_5 <= pte_addr[31:0];
      end
    end
    if (metaReset) begin
      tags_6 <= 32'h0;
    end else if (_T_28) begin
      if (3'h6 == r) begin
        tags_6 <= pte_addr[31:0];
      end
    end
    if (metaReset) begin
      tags_7 <= 32'h0;
    end else if (_T_28) begin
      if (3'h7 == r) begin
        tags_7 <= pte_addr[31:0];
      end
    end
    if (metaReset) begin
      data_0 <= 20'h0;
    end else if (_T_28) begin
      if (3'h0 == r) begin
        data_0 <= res_ppn[19:0];
      end
    end
    if (metaReset) begin
      data_1 <= 20'h0;
    end else if (_T_28) begin
      if (3'h1 == r) begin
        data_1 <= res_ppn[19:0];
      end
    end
    if (metaReset) begin
      data_2 <= 20'h0;
    end else if (_T_28) begin
      if (3'h2 == r) begin
        data_2 <= res_ppn[19:0];
      end
    end
    if (metaReset) begin
      data_3 <= 20'h0;
    end else if (_T_28) begin
      if (3'h3 == r) begin
        data_3 <= res_ppn[19:0];
      end
    end
    if (metaReset) begin
      data_4 <= 20'h0;
    end else if (_T_28) begin
      if (3'h4 == r) begin
        data_4 <= res_ppn[19:0];
      end
    end
    if (metaReset) begin
      data_5 <= 20'h0;
    end else if (_T_28) begin
      if (3'h5 == r) begin
        data_5 <= res_ppn[19:0];
      end
    end
    if (metaReset) begin
      data_6 <= 20'h0;
    end else if (_T_28) begin
      if (3'h6 == r) begin
        data_6 <= res_ppn[19:0];
      end
    end
    if (metaReset) begin
      data_7 <= 20'h0;
    end else if (_T_28) begin
      if (3'h7 == r) begin
        data_7 <= res_ppn[19:0];
      end
    end
    if (metaReset) begin
      pte_hit <= 1'h0;
    end else if (_T_100) begin
      pte_hit <= 1'h0;
    end else begin
      pte_hit <= _GEN_75;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_98) begin
          $fwrite(32'h80000002,"Assertion failed: PTE Cache Hit/Miss Performance Monitor Events are lower priority than L2TLB Hit event\n    at PTW.scala:198 assert(!(io.dpath.perf.l2hit && (io.dpath.perf.pte_miss || io.dpath.perf.pte_hit)),\n"); // @[PTW.scala 198:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_98) begin
          $fatal; // @[PTW.scala 198:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (mem_resp_valid & ~_T_123) begin
          $fwrite(32'h80000002,"Assertion failed\n    at PTW.scala:389 assert(state === s_wait3)\n"); // @[PTW.scala 389:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (mem_resp_valid & ~_T_123) begin
          $fatal; // @[PTW.scala 389:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_mem_s2_nack & ~_T_133) begin
          $fwrite(32'h80000002,"Assertion failed\n    at PTW.scala:406 assert(state === s_wait2)\n"); // @[PTW.scala 406:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_mem_s2_nack & ~_T_133) begin
          $fatal; // @[PTW.scala 406:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    PTW_state <= PTW_xor0;
    if (!(PTW_cov_read_data)) begin
      PTW_covSum <= PTW_covSum + 1'h1;
    end
    if (metaReset) begin
      PTW_metaAssert <= 1'h0;
    end else begin
      PTW_metaAssert <= PTW_metaAssert | PTW_or0;
    end
  end
  always @(posedge clock) begin
    if(PTW_cov_write_en & PTW_cov_write_mask) begin
      PTW_cov[PTW_cov_write_addr] <= PTW_cov_write_data; // @[Coverage map for PTW]
    end
  end
endmodule
module Rocket(
  input         clock,
  input         reset,
  input         io_hartid,
  input         io_interrupts_debug,
  input         io_interrupts_mtip,
  input         io_interrupts_msip,
  input         io_interrupts_meip,
  input         io_interrupts_seip,
  output        io_imem_might_request,
  output        io_imem_req_valid,
  output [39:0] io_imem_req_bits_pc,
  output        io_imem_req_bits_speculative,
  output        io_imem_sfence_valid,
  output        io_imem_sfence_bits_rs1,
  output        io_imem_sfence_bits_rs2,
  output [38:0] io_imem_sfence_bits_addr,
  output        io_imem_resp_ready,
  input         io_imem_resp_valid,
  input         io_imem_resp_bits_btb_taken,
  input         io_imem_resp_bits_btb_bridx,
  input  [4:0]  io_imem_resp_bits_btb_entry,
  input  [7:0]  io_imem_resp_bits_btb_bht_history,
  input  [39:0] io_imem_resp_bits_pc,
  input  [31:0] io_imem_resp_bits_data,
  input         io_imem_resp_bits_xcpt_pf_inst,
  input         io_imem_resp_bits_xcpt_ae_inst,
  input         io_imem_resp_bits_replay,
  output        io_imem_btb_update_valid,
  output [4:0]  io_imem_btb_update_bits_prediction_entry,
  output [38:0] io_imem_btb_update_bits_pc,
  output        io_imem_btb_update_bits_isValid,
  output [38:0] io_imem_btb_update_bits_br_pc,
  output [1:0]  io_imem_btb_update_bits_cfiType,
  output        io_imem_bht_update_valid,
  output [7:0]  io_imem_bht_update_bits_prediction_history,
  output [38:0] io_imem_bht_update_bits_pc,
  output        io_imem_bht_update_bits_branch,
  output        io_imem_bht_update_bits_taken,
  output        io_imem_bht_update_bits_mispredict,
  output        io_imem_flush_icache,
  input         io_dmem_req_ready,
  output        io_dmem_req_valid,
  output [39:0] io_dmem_req_bits_addr,
  output [6:0]  io_dmem_req_bits_tag,
  output [4:0]  io_dmem_req_bits_cmd,
  output [1:0]  io_dmem_req_bits_size,
  output        io_dmem_req_bits_signed,
  output        io_dmem_s1_kill,
  output [63:0] io_dmem_s1_data_data,
  input         io_dmem_s2_nack,
  input         io_dmem_resp_valid,
  input  [6:0]  io_dmem_resp_bits_tag,
  input  [1:0]  io_dmem_resp_bits_size,
  input  [63:0] io_dmem_resp_bits_data,
  input         io_dmem_resp_bits_replay,
  input         io_dmem_resp_bits_has_data,
  input  [63:0] io_dmem_resp_bits_data_word_bypass,
  input         io_dmem_replay_next,
  input         io_dmem_s2_xcpt_ma_ld,
  input         io_dmem_s2_xcpt_ma_st,
  input         io_dmem_s2_xcpt_pf_ld,
  input         io_dmem_s2_xcpt_pf_st,
  input         io_dmem_s2_xcpt_ae_ld,
  input         io_dmem_s2_xcpt_ae_st,
  input         io_dmem_ordered,
  input         io_dmem_perf_release,
  input         io_dmem_perf_grant,
  output [3:0]  io_ptw_ptbr_mode,
  output [43:0] io_ptw_ptbr_ppn,
  output        io_ptw_sfence_valid,
  output        io_ptw_sfence_bits_rs1,
  output        io_ptw_status_debug,
  output [1:0]  io_ptw_status_dprv,
  output [1:0]  io_ptw_status_prv,
  output        io_ptw_status_mxr,
  output        io_ptw_status_sum,
  output        io_ptw_pmp_0_cfg_l,
  output [1:0]  io_ptw_pmp_0_cfg_a,
  output        io_ptw_pmp_0_cfg_x,
  output        io_ptw_pmp_0_cfg_w,
  output        io_ptw_pmp_0_cfg_r,
  output [29:0] io_ptw_pmp_0_addr,
  output [31:0] io_ptw_pmp_0_mask,
  output        io_ptw_pmp_1_cfg_l,
  output [1:0]  io_ptw_pmp_1_cfg_a,
  output        io_ptw_pmp_1_cfg_x,
  output        io_ptw_pmp_1_cfg_w,
  output        io_ptw_pmp_1_cfg_r,
  output [29:0] io_ptw_pmp_1_addr,
  output [31:0] io_ptw_pmp_1_mask,
  output        io_ptw_pmp_2_cfg_l,
  output [1:0]  io_ptw_pmp_2_cfg_a,
  output        io_ptw_pmp_2_cfg_x,
  output        io_ptw_pmp_2_cfg_w,
  output        io_ptw_pmp_2_cfg_r,
  output [29:0] io_ptw_pmp_2_addr,
  output [31:0] io_ptw_pmp_2_mask,
  output        io_ptw_pmp_3_cfg_l,
  output [1:0]  io_ptw_pmp_3_cfg_a,
  output        io_ptw_pmp_3_cfg_x,
  output        io_ptw_pmp_3_cfg_w,
  output        io_ptw_pmp_3_cfg_r,
  output [29:0] io_ptw_pmp_3_addr,
  output [31:0] io_ptw_pmp_3_mask,
  output        io_ptw_pmp_4_cfg_l,
  output [1:0]  io_ptw_pmp_4_cfg_a,
  output        io_ptw_pmp_4_cfg_x,
  output        io_ptw_pmp_4_cfg_w,
  output        io_ptw_pmp_4_cfg_r,
  output [29:0] io_ptw_pmp_4_addr,
  output [31:0] io_ptw_pmp_4_mask,
  output        io_ptw_pmp_5_cfg_l,
  output [1:0]  io_ptw_pmp_5_cfg_a,
  output        io_ptw_pmp_5_cfg_x,
  output        io_ptw_pmp_5_cfg_w,
  output        io_ptw_pmp_5_cfg_r,
  output [29:0] io_ptw_pmp_5_addr,
  output [31:0] io_ptw_pmp_5_mask,
  output        io_ptw_pmp_6_cfg_l,
  output [1:0]  io_ptw_pmp_6_cfg_a,
  output        io_ptw_pmp_6_cfg_x,
  output        io_ptw_pmp_6_cfg_w,
  output        io_ptw_pmp_6_cfg_r,
  output [29:0] io_ptw_pmp_6_addr,
  output [31:0] io_ptw_pmp_6_mask,
  output        io_ptw_pmp_7_cfg_l,
  output [1:0]  io_ptw_pmp_7_cfg_a,
  output        io_ptw_pmp_7_cfg_x,
  output        io_ptw_pmp_7_cfg_w,
  output        io_ptw_pmp_7_cfg_r,
  output [29:0] io_ptw_pmp_7_addr,
  output [31:0] io_ptw_pmp_7_mask,
  output [63:0] io_ptw_customCSRs_csrs_0_value,
  output [31:0] io_fpu_inst,
  output [63:0] io_fpu_fromint_data,
  output [2:0]  io_fpu_fcsr_rm,
  input         io_fpu_fcsr_flags_valid,
  input  [4:0]  io_fpu_fcsr_flags_bits,
  input  [63:0] io_fpu_store_data,
  input  [63:0] io_fpu_toint_data,
  output        io_fpu_dmem_resp_val,
  output [2:0]  io_fpu_dmem_resp_type,
  output [4:0]  io_fpu_dmem_resp_tag,
  output [63:0] io_fpu_dmem_resp_data,
  output        io_fpu_valid,
  input         io_fpu_fcsr_rdy,
  input         io_fpu_nack_mem,
  input         io_fpu_illegal_rm,
  output        io_fpu_killx,
  output        io_fpu_killm,
  input         io_fpu_dec_wen,
  input         io_fpu_dec_ren1,
  input         io_fpu_dec_ren2,
  input         io_fpu_dec_ren3,
  input         io_fpu_sboard_set,
  input         io_fpu_sboard_clr,
  input  [4:0]  io_fpu_sboard_clra,
  output        io_trace_0_valid,
  output [39:0] io_trace_0_iaddr,
  output [31:0] io_trace_0_insn,
  output [2:0]  io_trace_0_priv,
  output        io_trace_0_exception,
  output        io_trace_0_interrupt,
  output [63:0] io_trace_0_cause,
  output [39:0] io_trace_0_tval,
  output        io_wfi,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset,
  input         PlusArgTimeout_halt,
  input         csr_halt,
  input         ibuf_halt,
  input         div_halt
);
  wire  ibuf_clock; // @[RocketCore.scala 254:20]
  wire  ibuf_reset; // @[RocketCore.scala 254:20]
  wire  ibuf_io_imem_ready; // @[RocketCore.scala 254:20]
  wire  ibuf_io_imem_valid; // @[RocketCore.scala 254:20]
  wire  ibuf_io_imem_bits_btb_taken; // @[RocketCore.scala 254:20]
  wire  ibuf_io_imem_bits_btb_bridx; // @[RocketCore.scala 254:20]
  wire [4:0] ibuf_io_imem_bits_btb_entry; // @[RocketCore.scala 254:20]
  wire [7:0] ibuf_io_imem_bits_btb_bht_history; // @[RocketCore.scala 254:20]
  wire [39:0] ibuf_io_imem_bits_pc; // @[RocketCore.scala 254:20]
  wire [31:0] ibuf_io_imem_bits_data; // @[RocketCore.scala 254:20]
  wire  ibuf_io_imem_bits_xcpt_pf_inst; // @[RocketCore.scala 254:20]
  wire  ibuf_io_imem_bits_xcpt_ae_inst; // @[RocketCore.scala 254:20]
  wire  ibuf_io_imem_bits_replay; // @[RocketCore.scala 254:20]
  wire  ibuf_io_kill; // @[RocketCore.scala 254:20]
  wire [39:0] ibuf_io_pc; // @[RocketCore.scala 254:20]
  wire [4:0] ibuf_io_btb_resp_entry; // @[RocketCore.scala 254:20]
  wire [7:0] ibuf_io_btb_resp_bht_history; // @[RocketCore.scala 254:20]
  wire  ibuf_io_inst_0_ready; // @[RocketCore.scala 254:20]
  wire  ibuf_io_inst_0_valid; // @[RocketCore.scala 254:20]
  wire  ibuf_io_inst_0_bits_xcpt0_pf_inst; // @[RocketCore.scala 254:20]
  wire  ibuf_io_inst_0_bits_xcpt0_ae_inst; // @[RocketCore.scala 254:20]
  wire  ibuf_io_inst_0_bits_xcpt1_pf_inst; // @[RocketCore.scala 254:20]
  wire  ibuf_io_inst_0_bits_xcpt1_ae_inst; // @[RocketCore.scala 254:20]
  wire  ibuf_io_inst_0_bits_replay; // @[RocketCore.scala 254:20]
  wire  ibuf_io_inst_0_bits_rvc; // @[RocketCore.scala 254:20]
  wire [31:0] ibuf_io_inst_0_bits_inst_bits; // @[RocketCore.scala 254:20]
  wire [4:0] ibuf_io_inst_0_bits_inst_rd; // @[RocketCore.scala 254:20]
  wire [4:0] ibuf_io_inst_0_bits_inst_rs1; // @[RocketCore.scala 254:20]
  wire [4:0] ibuf_io_inst_0_bits_inst_rs2; // @[RocketCore.scala 254:20]
  wire [4:0] ibuf_io_inst_0_bits_inst_rs3; // @[RocketCore.scala 254:20]
  wire [31:0] ibuf_io_inst_0_bits_raw; // @[RocketCore.scala 254:20]
  wire [29:0] ibuf_io_covSum; // @[RocketCore.scala 254:20]
  wire  ibuf_metaAssert; // @[RocketCore.scala 254:20]
  wire  ibuf_metaReset; // @[RocketCore.scala 254:20]
  reg [63:0] rf [0:30]; // @[RocketCore.scala 1015:15]
  reg [63:0] _RAND_0;
  wire [63:0] rf_id_rs_MPORT_data; // @[RocketCore.scala 1015:15]
  wire [4:0] rf_id_rs_MPORT_addr; // @[RocketCore.scala 1015:15]
  reg [63:0] _RAND_1;
  wire [63:0] rf_id_rs_MPORT_1_data; // @[RocketCore.scala 1015:15]
  wire [4:0] rf_id_rs_MPORT_1_addr; // @[RocketCore.scala 1015:15]
  reg [63:0] _RAND_2;
  wire [63:0] rf_MPORT_data; // @[RocketCore.scala 1015:15]
  wire [4:0] rf_MPORT_addr; // @[RocketCore.scala 1015:15]
  wire  rf_MPORT_mask; // @[RocketCore.scala 1015:15]
  wire  rf_MPORT_en; // @[RocketCore.scala 1015:15]
  wire  csr_clock; // @[RocketCore.scala 282:19]
  wire  csr_reset; // @[RocketCore.scala 282:19]
  wire  csr_io_ungated_clock; // @[RocketCore.scala 282:19]
  wire  csr_io_interrupts_debug; // @[RocketCore.scala 282:19]
  wire  csr_io_interrupts_mtip; // @[RocketCore.scala 282:19]
  wire  csr_io_interrupts_msip; // @[RocketCore.scala 282:19]
  wire  csr_io_interrupts_meip; // @[RocketCore.scala 282:19]
  wire  csr_io_interrupts_seip; // @[RocketCore.scala 282:19]
  wire  csr_io_hartid; // @[RocketCore.scala 282:19]
  wire [11:0] csr_io_rw_addr; // @[RocketCore.scala 282:19]
  wire [2:0] csr_io_rw_cmd; // @[RocketCore.scala 282:19]
  wire [63:0] csr_io_rw_rdata; // @[RocketCore.scala 282:19]
  wire [63:0] csr_io_rw_wdata; // @[RocketCore.scala 282:19]
  wire [11:0] csr_io_decode_0_csr; // @[RocketCore.scala 282:19]
  wire  csr_io_decode_0_fp_illegal; // @[RocketCore.scala 282:19]
  wire  csr_io_decode_0_fp_csr; // @[RocketCore.scala 282:19]
  wire  csr_io_decode_0_read_illegal; // @[RocketCore.scala 282:19]
  wire  csr_io_decode_0_write_illegal; // @[RocketCore.scala 282:19]
  wire  csr_io_decode_0_write_flush; // @[RocketCore.scala 282:19]
  wire  csr_io_decode_0_system_illegal; // @[RocketCore.scala 282:19]
  wire  csr_io_csr_stall; // @[RocketCore.scala 282:19]
  wire  csr_io_eret; // @[RocketCore.scala 282:19]
  wire  csr_io_singleStep; // @[RocketCore.scala 282:19]
  wire  csr_io_status_debug; // @[RocketCore.scala 282:19]
  wire  csr_io_status_cease; // @[RocketCore.scala 282:19]
  wire  csr_io_status_wfi; // @[RocketCore.scala 282:19]
  wire [31:0] csr_io_status_isa; // @[RocketCore.scala 282:19]
  wire [1:0] csr_io_status_dprv; // @[RocketCore.scala 282:19]
  wire [1:0] csr_io_status_prv; // @[RocketCore.scala 282:19]
  wire  csr_io_status_sd; // @[RocketCore.scala 282:19]
  wire [26:0] csr_io_status_zero2; // @[RocketCore.scala 282:19]
  wire [1:0] csr_io_status_sxl; // @[RocketCore.scala 282:19]
  wire [1:0] csr_io_status_uxl; // @[RocketCore.scala 282:19]
  wire  csr_io_status_sd_rv32; // @[RocketCore.scala 282:19]
  wire [7:0] csr_io_status_zero1; // @[RocketCore.scala 282:19]
  wire  csr_io_status_tsr; // @[RocketCore.scala 282:19]
  wire  csr_io_status_tw; // @[RocketCore.scala 282:19]
  wire  csr_io_status_tvm; // @[RocketCore.scala 282:19]
  wire  csr_io_status_mxr; // @[RocketCore.scala 282:19]
  wire  csr_io_status_sum; // @[RocketCore.scala 282:19]
  wire  csr_io_status_mprv; // @[RocketCore.scala 282:19]
  wire [1:0] csr_io_status_xs; // @[RocketCore.scala 282:19]
  wire [1:0] csr_io_status_fs; // @[RocketCore.scala 282:19]
  wire [1:0] csr_io_status_mpp; // @[RocketCore.scala 282:19]
  wire [1:0] csr_io_status_vs; // @[RocketCore.scala 282:19]
  wire  csr_io_status_spp; // @[RocketCore.scala 282:19]
  wire  csr_io_status_mpie; // @[RocketCore.scala 282:19]
  wire  csr_io_status_hpie; // @[RocketCore.scala 282:19]
  wire  csr_io_status_spie; // @[RocketCore.scala 282:19]
  wire  csr_io_status_upie; // @[RocketCore.scala 282:19]
  wire  csr_io_status_mie; // @[RocketCore.scala 282:19]
  wire  csr_io_status_hie; // @[RocketCore.scala 282:19]
  wire  csr_io_status_sie; // @[RocketCore.scala 282:19]
  wire  csr_io_status_uie; // @[RocketCore.scala 282:19]
  wire [3:0] csr_io_ptbr_mode; // @[RocketCore.scala 282:19]
  wire [43:0] csr_io_ptbr_ppn; // @[RocketCore.scala 282:19]
  wire [39:0] csr_io_evec; // @[RocketCore.scala 282:19]
  wire  csr_io_exception; // @[RocketCore.scala 282:19]
  wire  csr_io_retire; // @[RocketCore.scala 282:19]
  wire [63:0] csr_io_cause; // @[RocketCore.scala 282:19]
  wire [39:0] csr_io_pc; // @[RocketCore.scala 282:19]
  wire [39:0] csr_io_tval; // @[RocketCore.scala 282:19]
  wire [63:0] csr_io_time; // @[RocketCore.scala 282:19]
  wire [2:0] csr_io_fcsr_rm; // @[RocketCore.scala 282:19]
  wire  csr_io_fcsr_flags_valid; // @[RocketCore.scala 282:19]
  wire [4:0] csr_io_fcsr_flags_bits; // @[RocketCore.scala 282:19]
  wire  csr_io_interrupt; // @[RocketCore.scala 282:19]
  wire [63:0] csr_io_interrupt_cause; // @[RocketCore.scala 282:19]
  wire  csr_io_bp_0_control_action; // @[RocketCore.scala 282:19]
  wire [1:0] csr_io_bp_0_control_tmatch; // @[RocketCore.scala 282:19]
  wire  csr_io_bp_0_control_m; // @[RocketCore.scala 282:19]
  wire  csr_io_bp_0_control_s; // @[RocketCore.scala 282:19]
  wire  csr_io_bp_0_control_u; // @[RocketCore.scala 282:19]
  wire  csr_io_bp_0_control_x; // @[RocketCore.scala 282:19]
  wire  csr_io_bp_0_control_w; // @[RocketCore.scala 282:19]
  wire  csr_io_bp_0_control_r; // @[RocketCore.scala 282:19]
  wire [38:0] csr_io_bp_0_address; // @[RocketCore.scala 282:19]
  wire  csr_io_pmp_0_cfg_l; // @[RocketCore.scala 282:19]
  wire [1:0] csr_io_pmp_0_cfg_a; // @[RocketCore.scala 282:19]
  wire  csr_io_pmp_0_cfg_x; // @[RocketCore.scala 282:19]
  wire  csr_io_pmp_0_cfg_w; // @[RocketCore.scala 282:19]
  wire  csr_io_pmp_0_cfg_r; // @[RocketCore.scala 282:19]
  wire [29:0] csr_io_pmp_0_addr; // @[RocketCore.scala 282:19]
  wire [31:0] csr_io_pmp_0_mask; // @[RocketCore.scala 282:19]
  wire  csr_io_pmp_1_cfg_l; // @[RocketCore.scala 282:19]
  wire [1:0] csr_io_pmp_1_cfg_a; // @[RocketCore.scala 282:19]
  wire  csr_io_pmp_1_cfg_x; // @[RocketCore.scala 282:19]
  wire  csr_io_pmp_1_cfg_w; // @[RocketCore.scala 282:19]
  wire  csr_io_pmp_1_cfg_r; // @[RocketCore.scala 282:19]
  wire [29:0] csr_io_pmp_1_addr; // @[RocketCore.scala 282:19]
  wire [31:0] csr_io_pmp_1_mask; // @[RocketCore.scala 282:19]
  wire  csr_io_pmp_2_cfg_l; // @[RocketCore.scala 282:19]
  wire [1:0] csr_io_pmp_2_cfg_a; // @[RocketCore.scala 282:19]
  wire  csr_io_pmp_2_cfg_x; // @[RocketCore.scala 282:19]
  wire  csr_io_pmp_2_cfg_w; // @[RocketCore.scala 282:19]
  wire  csr_io_pmp_2_cfg_r; // @[RocketCore.scala 282:19]
  wire [29:0] csr_io_pmp_2_addr; // @[RocketCore.scala 282:19]
  wire [31:0] csr_io_pmp_2_mask; // @[RocketCore.scala 282:19]
  wire  csr_io_pmp_3_cfg_l; // @[RocketCore.scala 282:19]
  wire [1:0] csr_io_pmp_3_cfg_a; // @[RocketCore.scala 282:19]
  wire  csr_io_pmp_3_cfg_x; // @[RocketCore.scala 282:19]
  wire  csr_io_pmp_3_cfg_w; // @[RocketCore.scala 282:19]
  wire  csr_io_pmp_3_cfg_r; // @[RocketCore.scala 282:19]
  wire [29:0] csr_io_pmp_3_addr; // @[RocketCore.scala 282:19]
  wire [31:0] csr_io_pmp_3_mask; // @[RocketCore.scala 282:19]
  wire  csr_io_pmp_4_cfg_l; // @[RocketCore.scala 282:19]
  wire [1:0] csr_io_pmp_4_cfg_a; // @[RocketCore.scala 282:19]
  wire  csr_io_pmp_4_cfg_x; // @[RocketCore.scala 282:19]
  wire  csr_io_pmp_4_cfg_w; // @[RocketCore.scala 282:19]
  wire  csr_io_pmp_4_cfg_r; // @[RocketCore.scala 282:19]
  wire [29:0] csr_io_pmp_4_addr; // @[RocketCore.scala 282:19]
  wire [31:0] csr_io_pmp_4_mask; // @[RocketCore.scala 282:19]
  wire  csr_io_pmp_5_cfg_l; // @[RocketCore.scala 282:19]
  wire [1:0] csr_io_pmp_5_cfg_a; // @[RocketCore.scala 282:19]
  wire  csr_io_pmp_5_cfg_x; // @[RocketCore.scala 282:19]
  wire  csr_io_pmp_5_cfg_w; // @[RocketCore.scala 282:19]
  wire  csr_io_pmp_5_cfg_r; // @[RocketCore.scala 282:19]
  wire [29:0] csr_io_pmp_5_addr; // @[RocketCore.scala 282:19]
  wire [31:0] csr_io_pmp_5_mask; // @[RocketCore.scala 282:19]
  wire  csr_io_pmp_6_cfg_l; // @[RocketCore.scala 282:19]
  wire [1:0] csr_io_pmp_6_cfg_a; // @[RocketCore.scala 282:19]
  wire  csr_io_pmp_6_cfg_x; // @[RocketCore.scala 282:19]
  wire  csr_io_pmp_6_cfg_w; // @[RocketCore.scala 282:19]
  wire  csr_io_pmp_6_cfg_r; // @[RocketCore.scala 282:19]
  wire [29:0] csr_io_pmp_6_addr; // @[RocketCore.scala 282:19]
  wire [31:0] csr_io_pmp_6_mask; // @[RocketCore.scala 282:19]
  wire  csr_io_pmp_7_cfg_l; // @[RocketCore.scala 282:19]
  wire [1:0] csr_io_pmp_7_cfg_a; // @[RocketCore.scala 282:19]
  wire  csr_io_pmp_7_cfg_x; // @[RocketCore.scala 282:19]
  wire  csr_io_pmp_7_cfg_w; // @[RocketCore.scala 282:19]
  wire  csr_io_pmp_7_cfg_r; // @[RocketCore.scala 282:19]
  wire [29:0] csr_io_pmp_7_addr; // @[RocketCore.scala 282:19]
  wire [31:0] csr_io_pmp_7_mask; // @[RocketCore.scala 282:19]
  wire  csr_io_inhibit_cycle; // @[RocketCore.scala 282:19]
  wire [31:0] csr_io_inst_0; // @[RocketCore.scala 282:19]
  wire  csr_io_trace_0_valid; // @[RocketCore.scala 282:19]
  wire [39:0] csr_io_trace_0_iaddr; // @[RocketCore.scala 282:19]
  wire [31:0] csr_io_trace_0_insn; // @[RocketCore.scala 282:19]
  wire [2:0] csr_io_trace_0_priv; // @[RocketCore.scala 282:19]
  wire  csr_io_trace_0_exception; // @[RocketCore.scala 282:19]
  wire  csr_io_trace_0_interrupt; // @[RocketCore.scala 282:19]
  wire [63:0] csr_io_trace_0_cause; // @[RocketCore.scala 282:19]
  wire [39:0] csr_io_trace_0_tval; // @[RocketCore.scala 282:19]
  wire [63:0] csr_io_customCSRs_0_value; // @[RocketCore.scala 282:19]
  wire [29:0] csr_io_covSum; // @[RocketCore.scala 282:19]
  wire  csr_metaAssert; // @[RocketCore.scala 282:19]
  wire  csr_metaReset; // @[RocketCore.scala 282:19]
  wire  bpu_io_status_debug; // @[RocketCore.scala 323:19]
  wire [1:0] bpu_io_status_prv; // @[RocketCore.scala 323:19]
  wire  bpu_io_bp_0_control_action; // @[RocketCore.scala 323:19]
  wire [1:0] bpu_io_bp_0_control_tmatch; // @[RocketCore.scala 323:19]
  wire  bpu_io_bp_0_control_m; // @[RocketCore.scala 323:19]
  wire  bpu_io_bp_0_control_s; // @[RocketCore.scala 323:19]
  wire  bpu_io_bp_0_control_u; // @[RocketCore.scala 323:19]
  wire  bpu_io_bp_0_control_x; // @[RocketCore.scala 323:19]
  wire  bpu_io_bp_0_control_w; // @[RocketCore.scala 323:19]
  wire  bpu_io_bp_0_control_r; // @[RocketCore.scala 323:19]
  wire [38:0] bpu_io_bp_0_address; // @[RocketCore.scala 323:19]
  wire [38:0] bpu_io_pc; // @[RocketCore.scala 323:19]
  wire [38:0] bpu_io_ea; // @[RocketCore.scala 323:19]
  wire  bpu_io_xcpt_if; // @[RocketCore.scala 323:19]
  wire  bpu_io_xcpt_ld; // @[RocketCore.scala 323:19]
  wire  bpu_io_xcpt_st; // @[RocketCore.scala 323:19]
  wire  bpu_io_debug_if; // @[RocketCore.scala 323:19]
  wire  bpu_io_debug_ld; // @[RocketCore.scala 323:19]
  wire  bpu_io_debug_st; // @[RocketCore.scala 323:19]
  wire [29:0] bpu_io_covSum; // @[RocketCore.scala 323:19]
  wire  bpu_metaAssert; // @[RocketCore.scala 323:19]
  wire  alu_io_dw; // @[RocketCore.scala 385:19]
  wire [3:0] alu_io_fn; // @[RocketCore.scala 385:19]
  wire [63:0] alu_io_in2; // @[RocketCore.scala 385:19]
  wire [63:0] alu_io_in1; // @[RocketCore.scala 385:19]
  wire [63:0] alu_io_out; // @[RocketCore.scala 385:19]
  wire [63:0] alu_io_adder_out; // @[RocketCore.scala 385:19]
  wire  alu_io_cmp_out; // @[RocketCore.scala 385:19]
  wire [29:0] alu_io_covSum; // @[RocketCore.scala 385:19]
  wire  alu_metaAssert; // @[RocketCore.scala 385:19]
  wire  div_clock; // @[RocketCore.scala 409:19]
  wire  div_reset; // @[RocketCore.scala 409:19]
  wire  div_io_req_ready; // @[RocketCore.scala 409:19]
  wire  div_io_req_valid; // @[RocketCore.scala 409:19]
  wire [3:0] div_io_req_bits_fn; // @[RocketCore.scala 409:19]
  wire  div_io_req_bits_dw; // @[RocketCore.scala 409:19]
  wire [63:0] div_io_req_bits_in1; // @[RocketCore.scala 409:19]
  wire [63:0] div_io_req_bits_in2; // @[RocketCore.scala 409:19]
  wire [4:0] div_io_req_bits_tag; // @[RocketCore.scala 409:19]
  wire  div_io_kill; // @[RocketCore.scala 409:19]
  wire  div_io_resp_ready; // @[RocketCore.scala 409:19]
  wire  div_io_resp_valid; // @[RocketCore.scala 409:19]
  wire [63:0] div_io_resp_bits_data; // @[RocketCore.scala 409:19]
  wire [4:0] div_io_resp_bits_tag; // @[RocketCore.scala 409:19]
  wire [29:0] div_io_covSum; // @[RocketCore.scala 409:19]
  wire  div_metaAssert; // @[RocketCore.scala 409:19]
  wire  div_metaReset; // @[RocketCore.scala 409:19]
  wire  PlusArgTimeout_clock; // @[PlusArg.scala 89:11]
  wire  PlusArgTimeout_reset; // @[PlusArg.scala 89:11]
  wire [31:0] PlusArgTimeout_io_count; // @[PlusArg.scala 89:11]
  wire [29:0] PlusArgTimeout_io_covSum; // @[PlusArg.scala 89:11]
  wire  PlusArgTimeout_metaAssert; // @[PlusArg.scala 89:11]
  wire  PlusArgTimeout_metaReset; // @[PlusArg.scala 89:11]
  reg  id_reg_pause; // @[RocketCore.scala 114:25]
  reg [31:0] _RAND_3;
  reg  imem_might_request_reg; // @[RocketCore.scala 115:35]
  reg [31:0] _RAND_4;
  reg  ex_ctrl_fp; // @[RocketCore.scala 190:20]
  reg [31:0] _RAND_5;
  reg  ex_ctrl_branch; // @[RocketCore.scala 190:20]
  reg [31:0] _RAND_6;
  reg  ex_ctrl_jal; // @[RocketCore.scala 190:20]
  reg [31:0] _RAND_7;
  reg  ex_ctrl_jalr; // @[RocketCore.scala 190:20]
  reg [31:0] _RAND_8;
  reg  ex_ctrl_rxs2; // @[RocketCore.scala 190:20]
  reg [31:0] _RAND_9;
  reg [1:0] ex_ctrl_sel_alu2; // @[RocketCore.scala 190:20]
  reg [31:0] _RAND_10;
  reg [1:0] ex_ctrl_sel_alu1; // @[RocketCore.scala 190:20]
  reg [31:0] _RAND_11;
  reg [2:0] ex_ctrl_sel_imm; // @[RocketCore.scala 190:20]
  reg [31:0] _RAND_12;
  reg  ex_ctrl_alu_dw; // @[RocketCore.scala 190:20]
  reg [31:0] _RAND_13;
  reg [3:0] ex_ctrl_alu_fn; // @[RocketCore.scala 190:20]
  reg [31:0] _RAND_14;
  reg  ex_ctrl_mem; // @[RocketCore.scala 190:20]
  reg [31:0] _RAND_15;
  reg [4:0] ex_ctrl_mem_cmd; // @[RocketCore.scala 190:20]
  reg [31:0] _RAND_16;
  reg  ex_ctrl_wfd; // @[RocketCore.scala 190:20]
  reg [31:0] _RAND_17;
  reg  ex_ctrl_div; // @[RocketCore.scala 190:20]
  reg [31:0] _RAND_18;
  reg  ex_ctrl_wxd; // @[RocketCore.scala 190:20]
  reg [31:0] _RAND_19;
  reg [2:0] ex_ctrl_csr; // @[RocketCore.scala 190:20]
  reg [31:0] _RAND_20;
  reg  ex_ctrl_fence_i; // @[RocketCore.scala 190:20]
  reg [31:0] _RAND_21;
  reg  mem_ctrl_fp; // @[RocketCore.scala 191:21]
  reg [31:0] _RAND_22;
  reg  mem_ctrl_branch; // @[RocketCore.scala 191:21]
  reg [31:0] _RAND_23;
  reg  mem_ctrl_jal; // @[RocketCore.scala 191:21]
  reg [31:0] _RAND_24;
  reg  mem_ctrl_jalr; // @[RocketCore.scala 191:21]
  reg [31:0] _RAND_25;
  reg  mem_ctrl_mem; // @[RocketCore.scala 191:21]
  reg [31:0] _RAND_26;
  reg  mem_ctrl_wfd; // @[RocketCore.scala 191:21]
  reg [31:0] _RAND_27;
  reg  mem_ctrl_div; // @[RocketCore.scala 191:21]
  reg [31:0] _RAND_28;
  reg  mem_ctrl_wxd; // @[RocketCore.scala 191:21]
  reg [31:0] _RAND_29;
  reg [2:0] mem_ctrl_csr; // @[RocketCore.scala 191:21]
  reg [31:0] _RAND_30;
  reg  mem_ctrl_fence_i; // @[RocketCore.scala 191:21]
  reg [31:0] _RAND_31;
  reg  wb_ctrl_mem; // @[RocketCore.scala 192:20]
  reg [31:0] _RAND_32;
  reg  wb_ctrl_wfd; // @[RocketCore.scala 192:20]
  reg [31:0] _RAND_33;
  reg  wb_ctrl_div; // @[RocketCore.scala 192:20]
  reg [31:0] _RAND_34;
  reg  wb_ctrl_wxd; // @[RocketCore.scala 192:20]
  reg [31:0] _RAND_35;
  reg [2:0] wb_ctrl_csr; // @[RocketCore.scala 192:20]
  reg [31:0] _RAND_36;
  reg  wb_ctrl_fence_i; // @[RocketCore.scala 192:20]
  reg [31:0] _RAND_37;
  reg  ex_reg_xcpt_interrupt; // @[RocketCore.scala 194:35]
  reg [31:0] _RAND_38;
  reg  ex_reg_valid; // @[RocketCore.scala 195:35]
  reg [31:0] _RAND_39;
  reg  ex_reg_rvc; // @[RocketCore.scala 196:35]
  reg [31:0] _RAND_40;
  reg [4:0] ex_reg_btb_resp_entry; // @[RocketCore.scala 197:35]
  reg [31:0] _RAND_41;
  reg [7:0] ex_reg_btb_resp_bht_history; // @[RocketCore.scala 197:35]
  reg [31:0] _RAND_42;
  reg  ex_reg_xcpt; // @[RocketCore.scala 198:35]
  reg [31:0] _RAND_43;
  reg  ex_reg_flush_pipe; // @[RocketCore.scala 199:35]
  reg [31:0] _RAND_44;
  reg  ex_reg_load_use; // @[RocketCore.scala 200:35]
  reg [31:0] _RAND_45;
  reg [63:0] ex_reg_cause; // @[RocketCore.scala 201:35]
  reg [63:0] _RAND_46;
  reg  ex_reg_replay; // @[RocketCore.scala 202:26]
  reg [31:0] _RAND_47;
  reg [39:0] ex_reg_pc; // @[RocketCore.scala 203:22]
  reg [63:0] _RAND_48;
  reg [1:0] ex_reg_mem_size; // @[RocketCore.scala 204:28]
  reg [31:0] _RAND_49;
  reg [31:0] ex_reg_inst; // @[RocketCore.scala 205:24]
  reg [31:0] _RAND_50;
  reg [31:0] ex_reg_raw_inst; // @[RocketCore.scala 206:28]
  reg [31:0] _RAND_51;
  reg  mem_reg_xcpt_interrupt; // @[RocketCore.scala 211:36]
  reg [31:0] _RAND_52;
  reg  mem_reg_valid; // @[RocketCore.scala 212:36]
  reg [31:0] _RAND_53;
  reg  mem_reg_rvc; // @[RocketCore.scala 213:36]
  reg [31:0] _RAND_54;
  reg [4:0] mem_reg_btb_resp_entry; // @[RocketCore.scala 214:36]
  reg [31:0] _RAND_55;
  reg [7:0] mem_reg_btb_resp_bht_history; // @[RocketCore.scala 214:36]
  reg [31:0] _RAND_56;
  reg  mem_reg_xcpt; // @[RocketCore.scala 215:36]
  reg [31:0] _RAND_57;
  reg  mem_reg_replay; // @[RocketCore.scala 216:36]
  reg [31:0] _RAND_58;
  reg  mem_reg_flush_pipe; // @[RocketCore.scala 217:36]
  reg [31:0] _RAND_59;
  reg [63:0] mem_reg_cause; // @[RocketCore.scala 218:36]
  reg [63:0] _RAND_60;
  reg  mem_reg_slow_bypass; // @[RocketCore.scala 219:36]
  reg [31:0] _RAND_61;
  reg  mem_reg_load; // @[RocketCore.scala 220:36]
  reg [31:0] _RAND_62;
  reg  mem_reg_store; // @[RocketCore.scala 221:36]
  reg [31:0] _RAND_63;
  reg  mem_reg_sfence; // @[RocketCore.scala 222:27]
  reg [31:0] _RAND_64;
  reg [39:0] mem_reg_pc; // @[RocketCore.scala 223:23]
  reg [63:0] _RAND_65;
  reg [31:0] mem_reg_inst; // @[RocketCore.scala 224:25]
  reg [31:0] _RAND_66;
  reg [1:0] mem_reg_mem_size; // @[RocketCore.scala 225:29]
  reg [31:0] _RAND_67;
  reg [31:0] mem_reg_raw_inst; // @[RocketCore.scala 226:29]
  reg [31:0] _RAND_68;
  reg [63:0] mem_reg_wdata; // @[RocketCore.scala 229:26]
  reg [63:0] _RAND_69;
  reg [63:0] mem_reg_rs2; // @[RocketCore.scala 230:24]
  reg [63:0] _RAND_70;
  reg  mem_br_taken; // @[RocketCore.scala 231:25]
  reg [31:0] _RAND_71;
  reg  wb_reg_valid; // @[RocketCore.scala 235:35]
  reg [31:0] _RAND_72;
  reg  wb_reg_xcpt; // @[RocketCore.scala 236:35]
  reg [31:0] _RAND_73;
  reg  wb_reg_replay; // @[RocketCore.scala 237:35]
  reg [31:0] _RAND_74;
  reg  wb_reg_flush_pipe; // @[RocketCore.scala 238:35]
  reg [31:0] _RAND_75;
  reg [63:0] wb_reg_cause; // @[RocketCore.scala 239:35]
  reg [63:0] _RAND_76;
  reg  wb_reg_sfence; // @[RocketCore.scala 240:26]
  reg [31:0] _RAND_77;
  reg [39:0] wb_reg_pc; // @[RocketCore.scala 241:22]
  reg [63:0] _RAND_78;
  reg [1:0] wb_reg_mem_size; // @[RocketCore.scala 242:28]
  reg [31:0] _RAND_79;
  reg [31:0] wb_reg_inst; // @[RocketCore.scala 243:24]
  reg [31:0] _RAND_80;
  reg [31:0] wb_reg_raw_inst; // @[RocketCore.scala 244:28]
  reg [31:0] _RAND_81;
  reg [63:0] wb_reg_wdata; // @[RocketCore.scala 245:25]
  reg [63:0] _RAND_82;
  wire  replay_wb_common; // @[RocketCore.scala 637:42]
  wire  _T_83; // @[RocketCore.scala 615:19]
  wire  _T_84; // @[RocketCore.scala 615:34]
  wire  _T_95; // @[RocketCore.scala 975:26]
  wire  _T_86; // @[RocketCore.scala 616:34]
  wire  _T_96; // @[RocketCore.scala 975:26]
  wire  _T_88; // @[RocketCore.scala 617:34]
  wire  _T_97; // @[RocketCore.scala 975:26]
  wire  _T_90; // @[RocketCore.scala 618:34]
  wire  _T_98; // @[RocketCore.scala 975:26]
  wire  _T_92; // @[RocketCore.scala 619:34]
  wire  _T_99; // @[RocketCore.scala 975:26]
  wire  _T_94; // @[RocketCore.scala 620:34]
  wire  wb_xcpt; // @[RocketCore.scala 975:26]
  wire  _take_pc_wb_T; // @[RocketCore.scala 640:27]
  wire  _take_pc_wb_T_1; // @[RocketCore.scala 640:38]
  wire  take_pc_wb; // @[RocketCore.scala 640:53]
  wire  _ex_pc_valid_T; // @[RocketCore.scala 490:34]
  wire  ex_pc_valid; // @[RocketCore.scala 490:51]
  wire  _mem_npc_T; // @[RocketCore.scala 513:36]
  wire [24:0] a; // @[RocketCore.scala 989:23]
  wire  _mem_npc_msb_T; // @[RocketCore.scala 990:21]
  wire  _mem_npc_msb_T_1; // @[RocketCore.scala 990:34]
  wire  _mem_npc_msb_T_2; // @[RocketCore.scala 990:29]
  wire  msb; // @[RocketCore.scala 990:18]
  wire [38:0] mem_npc_lo; // @[RocketCore.scala 991:16]
  wire [39:0] _mem_npc_T_2; // @[RocketCore.scala 513:106]
  wire  _mem_br_target_T_1; // @[RocketCore.scala 510:25]
  wire  mem_br_target_sign; // @[RocketCore.scala 1037:53]
  wire  mem_br_target_hi_hi_hi; // @[Cat.scala 30:58]
  wire [10:0] mem_br_target_hi_hi_lo; // @[Cat.scala 30:58]
  wire [7:0] mem_br_target_hi_lo_hi; // @[Cat.scala 30:58]
  wire  mem_br_target_hi_lo_lo; // @[Cat.scala 30:58]
  wire [5:0] mem_br_target_lo_hi_hi; // @[RocketCore.scala 1043:66]
  wire [3:0] mem_br_target_lo_hi_lo; // @[RocketCore.scala 1045:57]
  wire [31:0] _mem_br_target_T_3; // @[RocketCore.scala 1051:53]
  wire [7:0] mem_br_target_hi_lo_hi_1; // @[Cat.scala 30:58]
  wire  mem_br_target_hi_lo_lo_1; // @[Cat.scala 30:58]
  wire [31:0] _mem_br_target_T_5; // @[RocketCore.scala 1051:53]
  wire [3:0] _mem_br_target_T_6; // @[RocketCore.scala 512:8]
  wire [31:0] _mem_br_target_T_7; // @[RocketCore.scala 511:8]
  wire [31:0] _mem_br_target_T_8; // @[RocketCore.scala 510:8]
  wire [39:0] _GEN_248; // @[RocketCore.scala 509:41]
  wire [39:0] mem_br_target; // @[RocketCore.scala 509:41]
  wire [39:0] _mem_npc_T_3; // @[RocketCore.scala 513:21]
  wire [39:0] mem_npc; // @[RocketCore.scala 513:141]
  wire  _mem_wrong_npc_T; // @[RocketCore.scala 515:30]
  wire  _mem_wrong_npc_T_1; // @[RocketCore.scala 516:31]
  wire  _mem_wrong_npc_T_2; // @[RocketCore.scala 516:62]
  wire  _mem_wrong_npc_T_3; // @[RocketCore.scala 516:8]
  wire  mem_wrong_npc; // @[RocketCore.scala 515:8]
  wire  _take_pc_mem_T; // @[RocketCore.scala 523:54]
  wire  take_pc_mem; // @[RocketCore.scala 523:32]
  wire  take_pc_mem_wb; // @[RocketCore.scala 250:35]
  wire [31:0] _id_ctrl_decoder_bit_T; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_bit_T_1; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_3; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_5; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_7; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_9; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_11; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_13; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_15; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_17; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_19; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_21; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_23; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_25; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_bit_T_26; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_bit_T_27; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_29; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_31; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_33; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_35; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_37; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_39; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_41; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_43; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_bit_T_44; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_bit_T_45; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_47; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_49; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_51; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_53; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_55; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_57; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_59; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_61; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_63; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_65; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_67; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_69; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_71; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_73; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_75; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_77; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_79; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_bit_T_80; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_bit_T_81; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_83; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_85; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_bit_T_86; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_bit_T_87; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_89; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_91; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_93; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_bit_T_94; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_bit_T_95; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_97; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_bit_T_98; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_bit_T_99; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_101; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_103; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_105; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_107; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_109; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_111; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_113; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_bit_T_114; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_bit_T_115; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_117; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_119; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_121; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_123; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_125; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_127; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_129; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_131; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_133; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_135; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_137; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_139; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_141; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_143; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_145; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_147; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_149; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_151; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_153; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_155; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_157; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_159; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_161; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_163; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_165; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_167; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_169; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_171; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_173; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_175; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_177; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_179; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_181; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_183; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_185; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_187; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_189; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_191; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_193; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_195; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_197; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_199; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_bit_T_200; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_bit_T_201; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_203; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_205; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_207; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_209; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_211; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_213; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_215; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_217; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_219; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_221; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_223; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_bit_T_224; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_bit_T_225; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_226; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_227; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_229; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_231; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_233; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_235; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_237; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_239; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_241; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_bit_T_242; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_bit_T_243; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_245; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_247; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_249; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_251; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_253; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_255; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_257; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_259; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_261; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_263; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_265; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_267; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_269; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_271; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_273; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_275; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_277; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_279; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_281; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_283; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_285; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_287; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_289; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_291; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_293; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_295; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_297; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_299; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_300; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_301; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_302; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_303; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_304; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_306; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_308; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_310; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_312; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_314; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_316; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_bit_T_318; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_319; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_320; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_321; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_322; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_323; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_324; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_325; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_326; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_327; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_328; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_329; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_330; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_331; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_332; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_333; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_334; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_335; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_336; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_337; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_338; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_339; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_340; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_341; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_342; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_343; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_344; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_345; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_346; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_347; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_348; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_349; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_350; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_351; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_352; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_353; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_354; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_355; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_356; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_357; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_358; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_359; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_360; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_361; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_362; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_363; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_364; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_365; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_366; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_367; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_368; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_369; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_370; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_371; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_372; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_373; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_374; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_375; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_376; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_377; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_378; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_379; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_380; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_381; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_382; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_383; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_384; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_385; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_386; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_387; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_388; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_389; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_390; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_391; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_392; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_393; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_394; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_395; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_396; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_397; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_398; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_399; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_400; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_401; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_402; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_403; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_404; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_405; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_406; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_407; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_408; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_409; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_410; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_411; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_412; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_413; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_414; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_415; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_416; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_417; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_418; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_419; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_420; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_421; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_422; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_423; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_424; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_425; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_426; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_427; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_428; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_429; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_430; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_431; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_432; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_433; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_434; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_435; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_436; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_437; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_438; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_439; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_440; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_441; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_442; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_443; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_444; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_445; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_446; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_447; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_448; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_449; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_450; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_451; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_452; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_453; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_454; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_455; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_456; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_457; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_458; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_459; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_460; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_461; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_462; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_463; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_464; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_465; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_466; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_467; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_468; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_469; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_470; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_471; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_472; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_473; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_474; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_475; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_476; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_477; // @[Decode.scala 15:30]
  wire  id_ctrl_decoder_0; // @[Decode.scala 15:30]
  wire [31:0] _id_ctrl_decoder_T; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_1; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_2; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_3; // @[Decode.scala 14:121]
  wire  id_ctrl_decoder_1; // @[Decode.scala 15:30]
  wire [31:0] _id_ctrl_decoder_T_5; // @[Decode.scala 14:65]
  wire  id_ctrl_decoder_3; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_7; // @[Decode.scala 14:65]
  wire  id_ctrl_decoder_4; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_9; // @[Decode.scala 14:65]
  wire  id_ctrl_decoder_5; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_11; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_12; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_13; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_14; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_15; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_16; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_17; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_18; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_T_20; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_T_21; // @[Decode.scala 15:30]
  wire  id_ctrl_decoder_6; // @[Decode.scala 15:30]
  wire [31:0] _id_ctrl_decoder_T_22; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_23; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_24; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_25; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_26; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_27; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_28; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_29; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_30; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_31; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_T_33; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_T_34; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_T_35; // @[Decode.scala 15:30]
  wire  id_ctrl_decoder_7; // @[Decode.scala 15:30]
  wire [31:0] _id_ctrl_decoder_T_36; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_37; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_38; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_39; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_40; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_41; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_42; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_43; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_44; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_45; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_T_47; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_T_48; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_T_49; // @[Decode.scala 15:30]
  wire  id_ctrl_decoder_lo; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_T_51; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_52; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_53; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_54; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_55; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_T_57; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_T_58; // @[Decode.scala 15:30]
  wire  id_ctrl_decoder_hi; // @[Decode.scala 15:30]
  wire [1:0] id_ctrl_decoder_9; // @[Cat.scala 30:58]
  wire [31:0] _id_ctrl_decoder_T_59; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_60; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_61; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_62; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_63; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_64; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_T_66; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_T_67; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_T_68; // @[Decode.scala 15:30]
  wire  id_ctrl_decoder_lo_1; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_T_70; // @[Decode.scala 14:121]
  wire  id_ctrl_decoder_hi_1; // @[Decode.scala 15:30]
  wire [1:0] id_ctrl_decoder_10; // @[Cat.scala 30:58]
  wire  _id_ctrl_decoder_T_73; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_T_75; // @[Decode.scala 14:121]
  wire  id_ctrl_decoder_lo_2; // @[Decode.scala 15:30]
  wire [31:0] _id_ctrl_decoder_T_77; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_78; // @[Decode.scala 14:121]
  wire  id_ctrl_decoder_hi_lo; // @[Decode.scala 15:30]
  wire [31:0] _id_ctrl_decoder_T_80; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_81; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_82; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_83; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_T_85; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_T_87; // @[Decode.scala 15:30]
  wire  id_ctrl_decoder_hi_hi; // @[Decode.scala 15:30]
  wire [2:0] id_ctrl_decoder_11; // @[Cat.scala 30:58]
  wire [31:0] _id_ctrl_decoder_T_88; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_89; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_90; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_91; // @[Decode.scala 14:121]
  wire  id_ctrl_decoder_12; // @[Decode.scala 15:30]
  wire [31:0] _id_ctrl_decoder_T_93; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_94; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_95; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_96; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_97; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_98; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_99; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_100; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_T_102; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_T_103; // @[Decode.scala 15:30]
  wire  id_ctrl_decoder_lo_lo; // @[Decode.scala 15:30]
  wire [31:0] _id_ctrl_decoder_T_104; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_105; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_106; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_107; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_T_109; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_110; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_111; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_112; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_113; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_114; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_115; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_116; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_117; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_T_119; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_T_120; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_T_121; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_T_122; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_T_123; // @[Decode.scala 15:30]
  wire  id_ctrl_decoder_lo_hi; // @[Decode.scala 15:30]
  wire [31:0] _id_ctrl_decoder_T_124; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_125; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_126; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_127; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_128; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_129; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_130; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_131; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_132; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_133; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_T_135; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_T_136; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_T_137; // @[Decode.scala 15:30]
  wire  id_ctrl_decoder_hi_lo_1; // @[Decode.scala 15:30]
  wire [31:0] _id_ctrl_decoder_T_138; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_139; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_140; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_141; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_142; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_143; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_T_145; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_T_146; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_T_147; // @[Decode.scala 15:30]
  wire  id_ctrl_decoder_hi_hi_1; // @[Decode.scala 15:30]
  wire [3:0] id_ctrl_decoder_13; // @[Cat.scala 30:58]
  wire  _id_ctrl_decoder_bit_T_479; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_480; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_481; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_482; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_483; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_484; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_485; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_486; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_487; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_488; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_489; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_490; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_491; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_492; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_493; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_494; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_495; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_496; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_497; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_498; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_499; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_500; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_501; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_502; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_503; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_504; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_505; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_506; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_507; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_508; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_509; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_510; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_511; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_512; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_513; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_bit_T_514; // @[Decode.scala 15:30]
  wire  id_ctrl_decoder_14; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_T_149; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_150; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_151; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_152; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_153; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_T_155; // @[Decode.scala 15:30]
  wire  id_ctrl_decoder_lo_lo_1; // @[Decode.scala 15:30]
  wire [31:0] _id_ctrl_decoder_T_156; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_157; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_158; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_159; // @[Decode.scala 14:121]
  wire  id_ctrl_decoder_lo_hi_1; // @[Decode.scala 15:30]
  wire [31:0] _id_ctrl_decoder_T_161; // @[Decode.scala 14:65]
  wire  id_ctrl_decoder_hi_hi_hi; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_163; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_164; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_165; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_166; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_T_168; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_T_169; // @[Decode.scala 15:30]
  wire  id_ctrl_decoder_hi_lo_2; // @[Decode.scala 15:30]
  wire [31:0] _id_ctrl_decoder_T_170; // @[Decode.scala 14:65]
  wire  id_ctrl_decoder_hi_hi_lo; // @[Decode.scala 14:121]
  wire [4:0] id_ctrl_decoder_15; // @[Cat.scala 30:58]
  wire [31:0] _id_ctrl_decoder_T_172; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_173; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_174; // @[Decode.scala 14:65]
  wire [31:0] _id_ctrl_decoder_T_176; // @[Decode.scala 14:65]
  wire  id_ctrl_decoder_18; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_189; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_190; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_T_192; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_T_194; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_T_195; // @[Decode.scala 15:30]
  wire  id_ctrl_decoder_19; // @[Decode.scala 15:30]
  wire [31:0] _id_ctrl_decoder_T_196; // @[Decode.scala 14:65]
  wire  id_ctrl_decoder_21; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_T_199; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_T_201; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_202; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_203; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_204; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_205; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_206; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_207; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_208; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_209; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_210; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_211; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_T_213; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_T_214; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_T_215; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_T_216; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_T_217; // @[Decode.scala 15:30]
  wire  id_ctrl_decoder_22; // @[Decode.scala 15:30]
  wire [31:0] _id_ctrl_decoder_T_218; // @[Decode.scala 14:65]
  wire  id_ctrl_decoder_lo_5; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_220; // @[Decode.scala 14:65]
  wire  id_ctrl_decoder_hi_lo_3; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_222; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_223; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_224; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_225; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_226; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_227; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_T_229; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_T_230; // @[Decode.scala 15:30]
  wire  _id_ctrl_decoder_T_231; // @[Decode.scala 15:30]
  wire  id_ctrl_decoder_hi_hi_3; // @[Decode.scala 15:30]
  wire [2:0] id_ctrl_decoder_23; // @[Cat.scala 30:58]
  wire [31:0] _id_ctrl_decoder_T_232; // @[Decode.scala 14:65]
  wire  id_ctrl_decoder_24; // @[Decode.scala 14:121]
  wire  id_ctrl_decoder_25; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_236; // @[Decode.scala 14:65]
  wire  id_ctrl_decoder_26; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_238; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_239; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_240; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_241; // @[Decode.scala 14:121]
  wire [31:0] _id_ctrl_decoder_T_242; // @[Decode.scala 14:65]
  wire  _id_ctrl_decoder_T_243; // @[Decode.scala 14:121]
  wire  _id_ctrl_decoder_T_245; // @[Decode.scala 15:30]
  wire  id_ctrl_decoder_27; // @[Decode.scala 15:30]
  wire [4:0] id_raddr3; // @[RocketCore.scala 267:72]
  wire [4:0] id_raddr2; // @[RocketCore.scala 267:72]
  wire [4:0] id_raddr1; // @[RocketCore.scala 267:72]
  wire [4:0] id_waddr; // @[RocketCore.scala 267:72]
  reg  id_reg_fence; // @[RocketCore.scala 274:25]
  reg [31:0] _RAND_83;
  wire [63:0] _id_rs_T_4; // @[RocketCore.scala 1022:25]
  wire [63:0] _id_rs_T_9; // @[RocketCore.scala 1022:25]
  wire  _id_csr_en_T; // @[package.scala 15:47]
  wire  _id_csr_en_T_1; // @[package.scala 15:47]
  wire  _id_csr_en_T_2; // @[package.scala 15:47]
  wire  _id_csr_en_T_3; // @[package.scala 72:59]
  wire  id_csr_en; // @[package.scala 72:59]
  wire  id_system_insn; // @[RocketCore.scala 284:36]
  wire  _id_csr_ren_T_3; // @[RocketCore.scala 285:81]
  wire  id_csr_ren; // @[RocketCore.scala 285:54]
  wire  _id_sfence_T; // @[RocketCore.scala 287:50]
  wire  id_sfence; // @[RocketCore.scala 287:31]
  wire  _id_csr_flush_T; // @[RocketCore.scala 288:32]
  wire  _id_csr_flush_T_2; // @[RocketCore.scala 288:64]
  wire  _id_csr_flush_T_3; // @[RocketCore.scala 288:79]
  wire  id_csr_flush; // @[RocketCore.scala 288:50]
  wire  _id_illegal_insn_T_4; // @[RocketCore.scala 297:34]
  wire  _id_illegal_insn_T_5; // @[RocketCore.scala 296:40]
  wire  _id_illegal_insn_T_8; // @[RocketCore.scala 298:17]
  wire  _id_illegal_insn_T_9; // @[RocketCore.scala 297:65]
  wire  _id_illegal_insn_T_10; // @[RocketCore.scala 299:48]
  wire  _id_illegal_insn_T_11; // @[RocketCore.scala 299:16]
  wire  _id_illegal_insn_T_12; // @[RocketCore.scala 298:48]
  wire  _id_illegal_insn_T_15; // @[RocketCore.scala 300:16]
  wire  _id_illegal_insn_T_16; // @[RocketCore.scala 299:70]
  wire  _id_illegal_insn_T_19; // @[RocketCore.scala 301:30]
  wire  _id_illegal_insn_T_20; // @[RocketCore.scala 300:47]
  wire  _id_illegal_insn_T_40; // @[RocketCore.scala 307:64]
  wire  _id_illegal_insn_T_41; // @[RocketCore.scala 307:49]
  wire  _id_illegal_insn_T_42; // @[RocketCore.scala 307:15]
  wire  _id_illegal_insn_T_43; // @[RocketCore.scala 306:81]
  wire  _id_illegal_insn_T_46; // @[RocketCore.scala 308:65]
  wire  _id_illegal_insn_T_47; // @[RocketCore.scala 308:31]
  wire  id_illegal_insn; // @[RocketCore.scala 307:99]
  wire  id_amo_aq; // @[RocketCore.scala 310:29]
  wire  id_amo_rl; // @[RocketCore.scala 311:29]
  wire [3:0] id_fence_succ; // @[RocketCore.scala 313:33]
  wire  _id_fence_next_T; // @[RocketCore.scala 314:52]
  wire  id_fence_next; // @[RocketCore.scala 314:37]
  wire  id_mem_busy; // @[RocketCore.scala 315:38]
  wire  _GEN_0; // @[RocketCore.scala 316:23]
  wire  _id_do_fence_x8_T_1; // @[RocketCore.scala 321:33]
  wire  _id_do_fence_x8_T_2; // @[RocketCore.scala 321:46]
  wire  _id_do_fence_x8_T_4; // @[RocketCore.scala 321:81]
  wire  _id_do_fence_x8_T_5; // @[RocketCore.scala 321:65]
  wire  id_do_fence_x8; // @[RocketCore.scala 321:17]
  wire  _T_1; // @[RocketCore.scala 975:26]
  wire  _T_2; // @[RocketCore.scala 975:26]
  wire  _T_3; // @[RocketCore.scala 975:26]
  wire  _T_4; // @[RocketCore.scala 975:26]
  wire  _T_5; // @[RocketCore.scala 975:26]
  wire  _T_6; // @[RocketCore.scala 975:26]
  wire  id_xcpt; // @[RocketCore.scala 975:26]
  wire [1:0] _T_7; // @[Mux.scala 47:69]
  wire [3:0] _T_8; // @[Mux.scala 47:69]
  wire [3:0] _T_9; // @[Mux.scala 47:69]
  wire [3:0] _T_10; // @[Mux.scala 47:69]
  wire [3:0] _T_11; // @[Mux.scala 47:69]
  wire [3:0] _T_12; // @[Mux.scala 47:69]
  wire [4:0] ex_waddr; // @[RocketCore.scala 359:29]
  wire [4:0] mem_waddr; // @[RocketCore.scala 360:31]
  wire [4:0] wb_waddr; // @[RocketCore.scala 361:29]
  wire  _T_23; // @[RocketCore.scala 364:19]
  wire  _T_24; // @[RocketCore.scala 365:20]
  wire  _T_26; // @[RocketCore.scala 365:36]
  wire  id_bypass_src_0_0; // @[RocketCore.scala 367:82]
  wire  _id_bypass_src_T_1; // @[RocketCore.scala 367:82]
  wire  id_bypass_src_0_1; // @[RocketCore.scala 367:74]
  wire  _id_bypass_src_T_2; // @[RocketCore.scala 367:82]
  wire  id_bypass_src_0_2; // @[RocketCore.scala 367:74]
  wire  id_bypass_src_0_3; // @[RocketCore.scala 367:74]
  wire  id_bypass_src_1_0; // @[RocketCore.scala 367:82]
  wire  _id_bypass_src_T_5; // @[RocketCore.scala 367:82]
  wire  id_bypass_src_1_1; // @[RocketCore.scala 367:74]
  wire  _id_bypass_src_T_6; // @[RocketCore.scala 367:82]
  wire  id_bypass_src_1_2; // @[RocketCore.scala 367:74]
  wire  id_bypass_src_1_3; // @[RocketCore.scala 367:74]
  reg  ex_reg_rs_bypass_0; // @[RocketCore.scala 371:29]
  reg [31:0] _RAND_84;
  reg  ex_reg_rs_bypass_1; // @[RocketCore.scala 371:29]
  reg [31:0] _RAND_85;
  reg [1:0] ex_reg_rs_lsb_0; // @[RocketCore.scala 372:26]
  reg [31:0] _RAND_86;
  reg [1:0] ex_reg_rs_lsb_1; // @[RocketCore.scala 372:26]
  reg [31:0] _RAND_87;
  reg [61:0] ex_reg_rs_msb_0; // @[RocketCore.scala 373:26]
  reg [63:0] _RAND_88;
  reg [61:0] ex_reg_rs_msb_1; // @[RocketCore.scala 373:26]
  reg [63:0] _RAND_89;
  wire  _ex_rs_T; // @[package.scala 32:86]
  wire [63:0] _ex_rs_T_1; // @[package.scala 32:76]
  wire  _ex_rs_T_2; // @[package.scala 32:86]
  wire [63:0] _ex_rs_T_3; // @[package.scala 32:76]
  wire  _ex_rs_T_4; // @[package.scala 32:86]
  wire [63:0] _ex_rs_T_5; // @[package.scala 32:76]
  wire [63:0] _ex_rs_T_6; // @[Cat.scala 30:58]
  wire  _ex_rs_T_7; // @[package.scala 32:86]
  wire [63:0] _ex_rs_T_8; // @[package.scala 32:76]
  wire  _ex_rs_T_9; // @[package.scala 32:86]
  wire [63:0] _ex_rs_T_10; // @[package.scala 32:76]
  wire  _ex_rs_T_11; // @[package.scala 32:86]
  wire [63:0] _ex_rs_T_12; // @[package.scala 32:76]
  wire [63:0] _ex_rs_T_13; // @[Cat.scala 30:58]
  wire [63:0] ex_rs_1; // @[RocketCore.scala 375:14]
  wire  _ex_imm_sign_T; // @[RocketCore.scala 1037:24]
  wire  _ex_imm_sign_T_2; // @[RocketCore.scala 1037:53]
  wire  ex_imm_sign; // @[RocketCore.scala 1037:19]
  wire  _ex_imm_b30_20_T; // @[RocketCore.scala 1038:26]
  wire [10:0] _ex_imm_b30_20_T_2; // @[RocketCore.scala 1038:49]
  wire  _ex_imm_b19_12_T; // @[RocketCore.scala 1039:26]
  wire  _ex_imm_b19_12_T_1; // @[RocketCore.scala 1039:43]
  wire  _ex_imm_b19_12_T_2; // @[RocketCore.scala 1039:36]
  wire [7:0] _ex_imm_b19_12_T_4; // @[RocketCore.scala 1039:73]
  wire  _ex_imm_b11_T_2; // @[RocketCore.scala 1040:33]
  wire  _ex_imm_b11_T_3; // @[RocketCore.scala 1041:23]
  wire  _ex_imm_b11_T_5; // @[RocketCore.scala 1041:44]
  wire  _ex_imm_b11_T_6; // @[RocketCore.scala 1042:23]
  wire  _ex_imm_b11_T_8; // @[RocketCore.scala 1042:43]
  wire  _ex_imm_b11_T_9; // @[RocketCore.scala 1042:18]
  wire  _ex_imm_b11_T_10; // @[RocketCore.scala 1041:18]
  wire [5:0] ex_imm_lo_hi_hi; // @[RocketCore.scala 1043:20]
  wire  _ex_imm_b4_1_T_1; // @[RocketCore.scala 1045:24]
  wire  _ex_imm_b4_1_T_3; // @[RocketCore.scala 1045:34]
  wire [3:0] _ex_imm_b4_1_T_8; // @[RocketCore.scala 1046:19]
  wire [3:0] _ex_imm_b4_1_T_9; // @[RocketCore.scala 1045:19]
  wire [3:0] ex_imm_lo_hi_lo; // @[RocketCore.scala 1044:19]
  wire  _ex_imm_b0_T_2; // @[RocketCore.scala 1048:22]
  wire  _ex_imm_b0_T_6; // @[RocketCore.scala 1049:17]
  wire  _ex_imm_b0_T_7; // @[RocketCore.scala 1048:17]
  wire  ex_imm_lo_lo; // @[RocketCore.scala 1047:17]
  wire  ex_imm_hi_lo_lo; // @[Cat.scala 30:58]
  wire [7:0] ex_imm_hi_lo_hi; // @[Cat.scala 30:58]
  wire [10:0] ex_imm_hi_hi_lo; // @[Cat.scala 30:58]
  wire  ex_imm_hi_hi_hi; // @[Cat.scala 30:58]
  wire [31:0] ex_imm; // @[RocketCore.scala 1051:53]
  wire [63:0] _ex_op1_T; // @[RocketCore.scala 378:24]
  wire  _ex_op1_T_2; // @[Mux.scala 80:60]
  wire [63:0] _ex_op1_T_3; // @[Mux.scala 80:57]
  wire  _ex_op1_T_4; // @[Mux.scala 80:60]
  wire [63:0] _ex_op2_T; // @[RocketCore.scala 381:24]
  wire [3:0] _ex_op2_T_1; // @[RocketCore.scala 383:19]
  wire  _ex_op2_T_2; // @[Mux.scala 80:60]
  wire [63:0] _ex_op2_T_3; // @[Mux.scala 80:57]
  wire  _ex_op2_T_4; // @[Mux.scala 80:60]
  wire [63:0] _ex_op2_T_5; // @[Mux.scala 80:57]
  wire  _ex_op2_T_6; // @[Mux.scala 80:60]
  wire  _ctrl_killd_T_1; // @[RocketCore.scala 784:40]
  wire  _ctrl_killd_T_2; // @[RocketCore.scala 784:71]
  wire  _T_123; // @[RocketCore.scala 714:55]
  wire  _T_124; // @[RocketCore.scala 714:42]
  wire  _data_hazard_ex_T; // @[RocketCore.scala 734:70]
  wire  _data_hazard_ex_T_1; // @[RocketCore.scala 984:27]
  wire  _T_125; // @[RocketCore.scala 715:55]
  wire  _T_126; // @[RocketCore.scala 715:42]
  wire  _data_hazard_ex_T_2; // @[RocketCore.scala 734:70]
  wire  _data_hazard_ex_T_3; // @[RocketCore.scala 984:27]
  wire  _data_hazard_ex_T_6; // @[RocketCore.scala 984:50]
  wire  _T_127; // @[RocketCore.scala 716:55]
  wire  _T_128; // @[RocketCore.scala 716:42]
  wire  _data_hazard_ex_T_4; // @[RocketCore.scala 734:70]
  wire  _data_hazard_ex_T_5; // @[RocketCore.scala 984:27]
  wire  _data_hazard_ex_T_7; // @[RocketCore.scala 984:50]
  wire  data_hazard_ex; // @[RocketCore.scala 734:36]
  wire  _ex_cannot_bypass_T; // @[RocketCore.scala 733:38]
  wire  _ex_cannot_bypass_T_1; // @[RocketCore.scala 733:48]
  wire  _ex_cannot_bypass_T_2; // @[RocketCore.scala 733:64]
  wire  _ex_cannot_bypass_T_4; // @[RocketCore.scala 733:94]
  wire  ex_cannot_bypass; // @[RocketCore.scala 733:109]
  wire  _id_ex_hazard_T; // @[RocketCore.scala 736:54]
  wire  _fp_data_hazard_ex_T_1; // @[RocketCore.scala 984:27]
  wire  _fp_data_hazard_ex_T_3; // @[RocketCore.scala 984:27]
  wire  _fp_data_hazard_ex_T_8; // @[RocketCore.scala 984:50]
  wire  _fp_data_hazard_ex_T_4; // @[RocketCore.scala 735:76]
  wire  _fp_data_hazard_ex_T_5; // @[RocketCore.scala 984:27]
  wire  _fp_data_hazard_ex_T_9; // @[RocketCore.scala 984:50]
  wire  _fp_data_hazard_ex_T_7; // @[RocketCore.scala 984:27]
  wire  _fp_data_hazard_ex_T_10; // @[RocketCore.scala 984:50]
  wire  fp_data_hazard_ex; // @[RocketCore.scala 735:39]
  wire  _id_ex_hazard_T_1; // @[RocketCore.scala 736:74]
  wire  id_ex_hazard; // @[RocketCore.scala 736:35]
  wire  _data_hazard_mem_T; // @[RocketCore.scala 743:72]
  wire  _data_hazard_mem_T_1; // @[RocketCore.scala 984:27]
  wire  _data_hazard_mem_T_2; // @[RocketCore.scala 743:72]
  wire  _data_hazard_mem_T_3; // @[RocketCore.scala 984:27]
  wire  _data_hazard_mem_T_6; // @[RocketCore.scala 984:50]
  wire  _data_hazard_mem_T_4; // @[RocketCore.scala 743:72]
  wire  _data_hazard_mem_T_5; // @[RocketCore.scala 984:27]
  wire  _data_hazard_mem_T_7; // @[RocketCore.scala 984:50]
  wire  data_hazard_mem; // @[RocketCore.scala 743:38]
  wire  _mem_cannot_bypass_T; // @[RocketCore.scala 742:40]
  wire  _mem_cannot_bypass_T_1; // @[RocketCore.scala 742:66]
  wire  _mem_cannot_bypass_T_2; // @[RocketCore.scala 742:50]
  wire  _mem_cannot_bypass_T_4; // @[RocketCore.scala 742:100]
  wire  mem_cannot_bypass; // @[RocketCore.scala 742:116]
  wire  _id_mem_hazard_T; // @[RocketCore.scala 745:57]
  wire  _fp_data_hazard_mem_T_1; // @[RocketCore.scala 984:27]
  wire  _fp_data_hazard_mem_T_3; // @[RocketCore.scala 984:27]
  wire  _fp_data_hazard_mem_T_8; // @[RocketCore.scala 984:50]
  wire  _fp_data_hazard_mem_T_4; // @[RocketCore.scala 744:78]
  wire  _fp_data_hazard_mem_T_5; // @[RocketCore.scala 984:27]
  wire  _fp_data_hazard_mem_T_9; // @[RocketCore.scala 984:50]
  wire  _fp_data_hazard_mem_T_7; // @[RocketCore.scala 984:27]
  wire  _fp_data_hazard_mem_T_10; // @[RocketCore.scala 984:50]
  wire  fp_data_hazard_mem; // @[RocketCore.scala 744:41]
  wire  _id_mem_hazard_T_1; // @[RocketCore.scala 745:78]
  wire  id_mem_hazard; // @[RocketCore.scala 745:37]
  wire  _ctrl_stalld_T; // @[RocketCore.scala 772:18]
  wire  _data_hazard_wb_T; // @[RocketCore.scala 749:70]
  wire  _data_hazard_wb_T_1; // @[RocketCore.scala 984:27]
  wire  _data_hazard_wb_T_2; // @[RocketCore.scala 749:70]
  wire  _data_hazard_wb_T_3; // @[RocketCore.scala 984:27]
  wire  _data_hazard_wb_T_6; // @[RocketCore.scala 984:50]
  wire  _data_hazard_wb_T_4; // @[RocketCore.scala 749:70]
  wire  _data_hazard_wb_T_5; // @[RocketCore.scala 984:27]
  wire  _data_hazard_wb_T_7; // @[RocketCore.scala 984:50]
  wire  data_hazard_wb; // @[RocketCore.scala 749:36]
  wire  wb_dcache_miss; // @[RocketCore.scala 491:36]
  wire  wb_set_sboard; // @[RocketCore.scala 636:35]
  wire  _id_wb_hazard_T; // @[RocketCore.scala 751:54]
  wire  _fp_data_hazard_wb_T_1; // @[RocketCore.scala 984:27]
  wire  _fp_data_hazard_wb_T_3; // @[RocketCore.scala 984:27]
  wire  _fp_data_hazard_wb_T_8; // @[RocketCore.scala 984:50]
  wire  _fp_data_hazard_wb_T_4; // @[RocketCore.scala 750:76]
  wire  _fp_data_hazard_wb_T_5; // @[RocketCore.scala 984:27]
  wire  _fp_data_hazard_wb_T_9; // @[RocketCore.scala 984:50]
  wire  _fp_data_hazard_wb_T_7; // @[RocketCore.scala 984:27]
  wire  _fp_data_hazard_wb_T_10; // @[RocketCore.scala 984:50]
  wire  fp_data_hazard_wb; // @[RocketCore.scala 750:39]
  wire  _id_wb_hazard_T_1; // @[RocketCore.scala 751:71]
  wire  id_wb_hazard; // @[RocketCore.scala 751:35]
  wire  _ctrl_stalld_T_1; // @[RocketCore.scala 772:35]
  reg [31:0] _r; // @[RocketCore.scala 1001:25]
  reg [31:0] _RAND_90;
  wire [31:0] r; // @[RocketCore.scala 1002:40]
  wire [31:0] _id_sboard_hazard_T; // @[RocketCore.scala 998:35]
  wire  dmem_resp_valid; // @[RocketCore.scala 646:44]
  wire  dmem_resp_replay; // @[RocketCore.scala 647:42]
  wire  dmem_resp_xpu; // @[RocketCore.scala 643:23]
  wire  _T_117; // @[RocketCore.scala 662:26]
  wire  ll_wen_x1; // @[Decoupled.scala 40:37]
  wire  ll_wen; // @[RocketCore.scala 662:44]
  wire [4:0] dmem_resp_waddr; // @[RocketCore.scala 645:46]
  wire [4:0] ll_waddr; // @[RocketCore.scala 662:44]
  wire  _id_sboard_hazard_T_2; // @[RocketCore.scala 726:70]
  wire  _id_sboard_hazard_T_3; // @[RocketCore.scala 726:58]
  wire  _id_sboard_hazard_T_5; // @[RocketCore.scala 729:77]
  wire  _id_sboard_hazard_T_6; // @[RocketCore.scala 984:27]
  wire [31:0] _id_sboard_hazard_T_7; // @[RocketCore.scala 998:35]
  wire  _id_sboard_hazard_T_9; // @[RocketCore.scala 726:70]
  wire  _id_sboard_hazard_T_10; // @[RocketCore.scala 726:58]
  wire  _id_sboard_hazard_T_12; // @[RocketCore.scala 729:77]
  wire  _id_sboard_hazard_T_13; // @[RocketCore.scala 984:27]
  wire  _id_sboard_hazard_T_21; // @[RocketCore.scala 984:50]
  wire [31:0] _id_sboard_hazard_T_14; // @[RocketCore.scala 998:35]
  wire  _id_sboard_hazard_T_16; // @[RocketCore.scala 726:70]
  wire  _id_sboard_hazard_T_17; // @[RocketCore.scala 726:58]
  wire  _id_sboard_hazard_T_19; // @[RocketCore.scala 729:77]
  wire  _id_sboard_hazard_T_20; // @[RocketCore.scala 984:27]
  wire  id_sboard_hazard; // @[RocketCore.scala 984:50]
  wire  _ctrl_stalld_T_2; // @[RocketCore.scala 772:51]
  wire  _ctrl_stalld_T_3; // @[RocketCore.scala 773:40]
  wire  _ctrl_stalld_T_4; // @[RocketCore.scala 773:57]
  wire  _ctrl_stalld_T_5; // @[RocketCore.scala 773:23]
  wire  _ctrl_stalld_T_6; // @[RocketCore.scala 772:71]
  wire  _ctrl_stalld_T_7; // @[RocketCore.scala 774:15]
  wire  _ctrl_stalld_T_9; // @[RocketCore.scala 774:42]
  wire  _ctrl_stalld_T_10; // @[RocketCore.scala 773:74]
  reg [31:0] id_stall_fpu__r; // @[RocketCore.scala 1001:25]
  reg [31:0] _RAND_91;
  wire [31:0] _id_stall_fpu_T_18; // @[RocketCore.scala 998:35]
  wire  _id_stall_fpu_T_20; // @[RocketCore.scala 984:27]
  wire [31:0] _id_stall_fpu_T_21; // @[RocketCore.scala 998:35]
  wire  _id_stall_fpu_T_23; // @[RocketCore.scala 984:27]
  wire  _id_stall_fpu_T_30; // @[RocketCore.scala 984:50]
  wire [31:0] _id_stall_fpu_T_24; // @[RocketCore.scala 998:35]
  wire  _id_stall_fpu_T_26; // @[RocketCore.scala 984:27]
  wire  _id_stall_fpu_T_31; // @[RocketCore.scala 984:50]
  wire [31:0] _id_stall_fpu_T_27; // @[RocketCore.scala 998:35]
  wire  _id_stall_fpu_T_29; // @[RocketCore.scala 984:27]
  wire  id_stall_fpu; // @[RocketCore.scala 984:50]
  wire  _ctrl_stalld_T_11; // @[RocketCore.scala 775:16]
  wire  _ctrl_stalld_T_12; // @[RocketCore.scala 774:62]
  reg  blocked; // @[RocketCore.scala 764:22]
  reg [31:0] _RAND_92;
  wire  dcache_blocked; // @[RocketCore.scala 766:13]
  wire  _ctrl_stalld_T_13; // @[RocketCore.scala 776:17]
  wire  _ctrl_stalld_T_14; // @[RocketCore.scala 775:32]
  wire  wb_wxd; // @[RocketCore.scala 635:29]
  wire  _ctrl_stalld_T_18; // @[RocketCore.scala 778:62]
  wire  _ctrl_stalld_T_19; // @[RocketCore.scala 778:40]
  wire  _ctrl_stalld_T_21; // @[RocketCore.scala 778:75]
  wire  _ctrl_stalld_T_22; // @[RocketCore.scala 778:17]
  wire  _ctrl_stalld_T_23; // @[RocketCore.scala 777:34]
  wire  _ctrl_stalld_T_26; // @[RocketCore.scala 779:15]
  wire  _ctrl_stalld_T_27; // @[RocketCore.scala 780:17]
  wire  ctrl_stalld; // @[RocketCore.scala 781:22]
  wire  _ctrl_killd_T_3; // @[RocketCore.scala 784:89]
  wire  ctrl_killd; // @[RocketCore.scala 784:104]
  wire  _ex_reg_replay_T_1; // @[RocketCore.scala 424:29]
  wire  _T_29; // @[RocketCore.scala 434:42]
  wire  _T_30; // @[RocketCore.scala 434:25]
  wire  _GEN_1; // @[RocketCore.scala 434:49]
  wire  _GEN_2; // @[RocketCore.scala 435:26]
  wire [1:0] _T_31; // @[RocketCore.scala 441:22]
  wire  _T_32; // @[RocketCore.scala 441:29]
  wire  _GEN_5; // @[RocketCore.scala 441:34]
  wire [1:0] _T_33; // @[RocketCore.scala 446:40]
  wire  _T_34; // @[RocketCore.scala 446:47]
  wire  _T_35; // @[RocketCore.scala 446:28]
  wire  _GEN_9; // @[RocketCore.scala 436:20]
  wire  _ex_reg_flush_pipe_T; // @[RocketCore.scala 451:42]
  wire  _T_37; // @[package.scala 15:47]
  wire  _T_38; // @[package.scala 72:59]
  wire [1:0] _ex_reg_mem_size_T_1; // @[Cat.scala 30:58]
  wire  _do_bypass_T; // @[RocketCore.scala 464:48]
  wire  _do_bypass_T_1; // @[RocketCore.scala 464:48]
  wire  do_bypass; // @[RocketCore.scala 464:48]
  wire  _T_40; // @[RocketCore.scala 468:23]
  wire  _wb_valid_T_1; // @[RocketCore.scala 670:31]
  wire  wb_valid; // @[RocketCore.scala 670:45]
  wire  wb_wen; // @[RocketCore.scala 671:25]
  wire  rf_wen; // @[RocketCore.scala 672:23]
  wire [4:0] rf_waddr; // @[RocketCore.scala 673:21]
  wire  _T_118; // @[RocketCore.scala 1027:16]
  wire  _T_121; // @[RocketCore.scala 1030:20]
  wire  _rf_wdata_T; // @[RocketCore.scala 674:38]
  wire [63:0] ll_wdata;
  wire  _rf_wdata_T_2; // @[RocketCore.scala 676:34]
  wire [63:0] _rf_wdata_T_4; // @[RocketCore.scala 676:21]
  wire [63:0] _rf_wdata_T_5; // @[RocketCore.scala 675:21]
  wire [63:0] rf_wdata; // @[RocketCore.scala 674:21]
  wire [63:0] _GEN_226; // @[RocketCore.scala 1030:31]
  wire [63:0] _GEN_233; // @[RocketCore.scala 1027:29]
  wire [63:0] id_rs_0; // @[RocketCore.scala 679:17]
  wire  _do_bypass_T_2; // @[RocketCore.scala 464:48]
  wire  _do_bypass_T_3; // @[RocketCore.scala 464:48]
  wire  do_bypass_1; // @[RocketCore.scala 464:48]
  wire  _T_42; // @[RocketCore.scala 468:23]
  wire  _T_122; // @[RocketCore.scala 1030:20]
  wire [63:0] _GEN_227; // @[RocketCore.scala 1030:31]
  wire [63:0] _GEN_234; // @[RocketCore.scala 1027:29]
  wire [63:0] id_rs_1; // @[RocketCore.scala 679:17]
  wire [31:0] inst; // @[RocketCore.scala 474:21]
  wire  _id_load_use_T; // @[RocketCore.scala 746:32]
  wire  id_load_use; // @[RocketCore.scala 746:51]
  wire  _T_44; // @[RocketCore.scala 480:21]
  wire  _T_45; // @[RocketCore.scala 480:41]
  wire  _replay_ex_structural_T_1; // @[RocketCore.scala 492:42]
  wire  _replay_ex_structural_T_3; // @[RocketCore.scala 493:42]
  wire  replay_ex_structural; // @[RocketCore.scala 492:64]
  wire  replay_ex_load_use; // @[RocketCore.scala 494:43]
  wire  _replay_ex_T; // @[RocketCore.scala 495:75]
  wire  _replay_ex_T_1; // @[RocketCore.scala 495:50]
  wire  replay_ex; // @[RocketCore.scala 495:33]
  wire  _ctrl_killx_T; // @[RocketCore.scala 496:35]
  wire  ctrl_killx; // @[RocketCore.scala 496:48]
  wire  _ex_slow_bypass_T; // @[RocketCore.scala 498:40]
  wire  _ex_slow_bypass_T_1; // @[RocketCore.scala 498:69]
  wire  ex_slow_bypass; // @[RocketCore.scala 498:50]
  wire  _ex_sfence_T_1; // @[RocketCore.scala 499:67]
  wire  ex_sfence; // @[RocketCore.scala 499:48]
  wire  ex_xcpt; // @[RocketCore.scala 502:28]
  wire  _mem_pc_valid_T; // @[RocketCore.scala 508:36]
  wire  mem_pc_valid; // @[RocketCore.scala 508:54]
  wire  _mem_npc_misaligned_T_3; // @[RocketCore.scala 517:56]
  wire  mem_npc_misaligned; // @[RocketCore.scala 517:70]
  wire  _mem_int_wdata_T_1; // @[RocketCore.scala 518:59]
  wire  _mem_int_wdata_T_2; // @[RocketCore.scala 518:41]
  wire [63:0] mem_int_wdata; // @[RocketCore.scala 518:119]
  wire  _mem_cfi_T; // @[RocketCore.scala 519:33]
  wire  mem_cfi; // @[RocketCore.scala 519:50]
  wire  _mem_cfi_taken_T_1; // @[RocketCore.scala 520:57]
  wire  mem_cfi_taken; // @[RocketCore.scala 520:74]
  wire  _T_56; // @[RocketCore.scala 532:23]
  wire  _mem_reg_load_T; // @[Consts.scala 81:31]
  wire  _mem_reg_load_T_1; // @[Consts.scala 81:48]
  wire  _mem_reg_load_T_2; // @[Consts.scala 81:41]
  wire  _mem_reg_load_T_4; // @[Consts.scala 81:58]
  wire  _mem_reg_load_T_5; // @[package.scala 15:47]
  wire  _mem_reg_load_T_6; // @[package.scala 15:47]
  wire  _mem_reg_load_T_7; // @[package.scala 15:47]
  wire  _mem_reg_load_T_8; // @[package.scala 15:47]
  wire  _mem_reg_load_T_9; // @[package.scala 72:59]
  wire  _mem_reg_load_T_10; // @[package.scala 72:59]
  wire  _mem_reg_load_T_11; // @[package.scala 72:59]
  wire  _mem_reg_load_T_12; // @[package.scala 15:47]
  wire  _mem_reg_load_T_13; // @[package.scala 15:47]
  wire  _mem_reg_load_T_14; // @[package.scala 15:47]
  wire  _mem_reg_load_T_15; // @[package.scala 15:47]
  wire  _mem_reg_load_T_16; // @[package.scala 15:47]
  wire  _mem_reg_load_T_17; // @[package.scala 72:59]
  wire  _mem_reg_load_T_18; // @[package.scala 72:59]
  wire  _mem_reg_load_T_19; // @[package.scala 72:59]
  wire  _mem_reg_load_T_20; // @[package.scala 72:59]
  wire  _mem_reg_load_T_21; // @[Consts.scala 79:44]
  wire  _mem_reg_load_T_22; // @[Consts.scala 81:75]
  wire  _mem_reg_load_T_23; // @[RocketCore.scala 539:33]
  wire  _mem_reg_store_T; // @[Consts.scala 82:32]
  wire  _mem_reg_store_T_1; // @[Consts.scala 82:49]
  wire  _mem_reg_store_T_2; // @[Consts.scala 82:42]
  wire  _mem_reg_store_T_4; // @[Consts.scala 82:59]
  wire  _mem_reg_store_T_22; // @[Consts.scala 82:76]
  wire  _mem_reg_store_T_23; // @[RocketCore.scala 540:34]
  wire [63:0] _mem_reg_wdata_T; // @[RocketCore.scala 552:25]
  wire  _T_58; // @[RocketCore.scala 555:56]
  wire  _T_59; // @[RocketCore.scala 555:24]
  wire  _mem_reg_rs2_T; // @[AMOALU.scala 26:19]
  wire [7:0] mem_reg_rs2_hi; // @[AMOALU.scala 26:66]
  wire [63:0] _mem_reg_rs2_T_1; // @[Cat.scala 30:58]
  wire  _mem_reg_rs2_T_2; // @[AMOALU.scala 26:19]
  wire [15:0] mem_reg_rs2_hi_3; // @[AMOALU.scala 26:66]
  wire [63:0] _mem_reg_rs2_T_3; // @[Cat.scala 30:58]
  wire  _mem_reg_rs2_T_4; // @[AMOALU.scala 26:19]
  wire [31:0] mem_reg_rs2_hi_5; // @[AMOALU.scala 26:66]
  wire [63:0] _mem_reg_rs2_T_5; // @[Cat.scala 30:58]
  wire  _T_60; // @[RocketCore.scala 559:24]
  wire  _GEN_77; // @[RocketCore.scala 559:48]
  wire  _GEN_78; // @[RocketCore.scala 559:48]
  wire  _mem_breakpoint_T; // @[RocketCore.scala 566:38]
  wire  _mem_breakpoint_T_1; // @[RocketCore.scala 566:75]
  wire  mem_breakpoint; // @[RocketCore.scala 566:57]
  wire  _mem_debug_breakpoint_T; // @[RocketCore.scala 567:44]
  wire  _mem_debug_breakpoint_T_1; // @[RocketCore.scala 567:82]
  wire  mem_debug_breakpoint; // @[RocketCore.scala 567:64]
  wire  mem_ldst_xcpt; // @[RocketCore.scala 975:26]
  wire [3:0] mem_ldst_cause; // @[Mux.scala 47:69]
  wire  _T_61; // @[RocketCore.scala 573:29]
  wire  _T_62; // @[RocketCore.scala 574:20]
  wire  _T_63; // @[RocketCore.scala 575:20]
  wire  _T_64; // @[RocketCore.scala 975:26]
  wire  mem_xcpt; // @[RocketCore.scala 975:26]
  wire [3:0] _T_65; // @[Mux.scala 47:69]
  wire  dcache_kill_mem; // @[RocketCore.scala 584:55]
  wire  _fpu_kill_mem_T; // @[RocketCore.scala 585:36]
  wire  fpu_kill_mem; // @[RocketCore.scala 585:51]
  wire  _replay_mem_T; // @[RocketCore.scala 586:37]
  wire  replay_mem; // @[RocketCore.scala 586:55]
  wire  _killm_common_T; // @[RocketCore.scala 587:38]
  wire  _killm_common_T_1; // @[RocketCore.scala 587:52]
  wire  killm_common; // @[RocketCore.scala 587:68]
  reg  div_io_kill_REG; // @[RocketCore.scala 588:37]
  reg [31:0] _RAND_93;
  wire  _ctrl_killm_T; // @[RocketCore.scala 589:33]
  wire  ctrl_killm; // @[RocketCore.scala 589:45]
  wire  _wb_reg_wdata_T_1; // @[RocketCore.scala 600:25]
  wire  _wb_reg_wdata_T_2; // @[RocketCore.scala 600:40]
  wire [2:0] _T_100; // @[Mux.scala 47:69]
  wire [3:0] _T_101; // @[Mux.scala 47:69]
  wire [3:0] _T_102; // @[Mux.scala 47:69]
  wire [3:0] _T_103; // @[Mux.scala 47:69]
  wire [3:0] _T_104; // @[Mux.scala 47:69]
  wire [63:0] wb_cause; // @[Mux.scala 47:69]
  wire  _T_105; // @[RocketCore.scala 979:38]
  wire  _T_107; // @[RocketCore.scala 979:38]
  wire  _T_109; // @[RocketCore.scala 979:38]
  wire  _T_111; // @[RocketCore.scala 979:38]
  wire  _T_113; // @[RocketCore.scala 979:38]
  wire  _T_115; // @[RocketCore.scala 979:38]
  wire  _csr_io_inst_0_T_1; // @[RocketCore.scala 687:73]
  wire [15:0] csr_io_inst_0_hi; // @[RocketCore.scala 687:50]
  wire [15:0] csr_io_inst_0_lo; // @[RocketCore.scala 687:119]
  wire  _tval_valid_T; // @[package.scala 15:47]
  wire  _tval_valid_T_1; // @[package.scala 15:47]
  wire  _tval_valid_T_6; // @[package.scala 15:47]
  wire  _tval_valid_T_9; // @[package.scala 15:47]
  wire  _tval_valid_T_10; // @[package.scala 72:59]
  wire  _tval_valid_T_11; // @[package.scala 72:59]
  wire  _tval_valid_T_12; // @[package.scala 72:59]
  wire  _tval_valid_T_13; // @[package.scala 72:59]
  wire  _tval_valid_T_14; // @[package.scala 72:59]
  wire  _tval_valid_T_15; // @[package.scala 72:59]
  wire  _tval_valid_T_16; // @[package.scala 72:59]
  wire  _tval_valid_T_17; // @[package.scala 72:59]
  wire  _tval_valid_T_18; // @[package.scala 72:59]
  wire  tval_valid; // @[RocketCore.scala 696:28]
  wire [24:0] a_1; // @[RocketCore.scala 989:23]
  wire  _csr_io_tval_msb_T; // @[RocketCore.scala 990:21]
  wire  _csr_io_tval_msb_T_1; // @[RocketCore.scala 990:34]
  wire  _csr_io_tval_msb_T_2; // @[RocketCore.scala 990:29]
  wire  msb_1; // @[RocketCore.scala 990:18]
  wire [38:0] csr_io_tval_lo; // @[RocketCore.scala 991:16]
  wire [39:0] _csr_io_tval_T; // @[Cat.scala 30:58]
  wire [2:0] _csr_io_rw_cmd_T; // @[CSR.scala 132:15]
  wire [31:0] _T_129; // @[RocketCore.scala 1005:62]
  wire [31:0] _T_130; // @[RocketCore.scala 1005:49]
  wire [31:0] _T_132; // @[RocketCore.scala 997:62]
  wire  _T_134; // @[RocketCore.scala 730:28]
  wire [31:0] _T_135; // @[RocketCore.scala 1005:62]
  wire [31:0] _T_136; // @[RocketCore.scala 1005:49]
  wire [31:0] _T_137; // @[RocketCore.scala 996:60]
  wire  _T_138; // @[RocketCore.scala 1008:17]
  wire  _id_stall_fpu_T; // @[RocketCore.scala 755:35]
  wire  _id_stall_fpu_T_1; // @[RocketCore.scala 755:50]
  wire  _id_stall_fpu_T_2; // @[RocketCore.scala 755:72]
  wire [31:0] _id_stall_fpu_T_4; // @[RocketCore.scala 1005:49]
  wire [31:0] _id_stall_fpu_T_5; // @[RocketCore.scala 996:60]
  wire  _id_stall_fpu_T_7; // @[RocketCore.scala 756:38]
  wire [31:0] _id_stall_fpu_T_8; // @[RocketCore.scala 1005:62]
  wire [31:0] _id_stall_fpu_T_9; // @[RocketCore.scala 1005:49]
  wire [31:0] _id_stall_fpu_T_11; // @[RocketCore.scala 997:62]
  wire  _id_stall_fpu_T_12; // @[RocketCore.scala 1008:17]
  wire [31:0] _id_stall_fpu_T_13; // @[RocketCore.scala 1005:62]
  wire [31:0] _id_stall_fpu_T_14; // @[RocketCore.scala 1005:49]
  wire [31:0] _id_stall_fpu_T_16; // @[RocketCore.scala 997:62]
  wire  _id_stall_fpu_T_17; // @[RocketCore.scala 1008:17]
  wire  _dcache_blocked_blocked_T_3; // @[RocketCore.scala 765:60]
  wire  _dcache_blocked_blocked_T_4; // @[RocketCore.scala 765:95]
  wire  _dcache_blocked_blocked_T_5; // @[RocketCore.scala 765:116]
  wire  _io_imem_req_bits_pc_T; // @[RocketCore.scala 789:17]
  wire [39:0] _io_imem_req_bits_pc_T_1; // @[RocketCore.scala 790:8]
  wire  _io_imem_flush_icache_T; // @[RocketCore.scala 792:40]
  wire  _io_imem_might_request_imem_might_request_reg_T; // @[RocketCore.scala 794:43]
  wire  _io_imem_btb_update_valid_T_1; // @[RocketCore.scala 806:45]
  wire  _io_imem_btb_update_valid_T_2; // @[RocketCore.scala 806:60]
  wire  _io_imem_btb_update_valid_T_4; // @[RocketCore.scala 806:90]
  wire  _io_imem_btb_update_bits_cfiType_T; // @[RocketCore.scala 809:23]
  wire  _io_imem_btb_update_bits_cfiType_T_2; // @[RocketCore.scala 809:41]
  wire [4:0] _io_imem_btb_update_bits_cfiType_T_5; // @[RocketCore.scala 810:62]
  wire  _io_imem_btb_update_bits_cfiType_T_6; // @[RocketCore.scala 810:62]
  wire  _io_imem_btb_update_bits_cfiType_T_7; // @[RocketCore.scala 810:23]
  wire [1:0] _io_imem_btb_update_bits_cfiType_T_10; // @[RocketCore.scala 810:8]
  wire [1:0] _io_imem_btb_update_bits_br_pc_T; // @[RocketCore.scala 814:74]
  wire [39:0] _GEN_250; // @[RocketCore.scala 814:69]
  wire [39:0] _io_imem_btb_update_bits_br_pc_T_2; // @[RocketCore.scala 814:69]
  wire [38:0] _io_imem_btb_update_bits_pc_T_1; // @[RocketCore.scala 815:66]
  wire [5:0] ex_dcache_tag; // @[Cat.scala 30:58]
  wire [24:0] a_2; // @[RocketCore.scala 989:23]
  wire  _io_dmem_req_bits_addr_msb_T; // @[RocketCore.scala 990:21]
  wire  _io_dmem_req_bits_addr_msb_T_1; // @[RocketCore.scala 990:34]
  wire  _io_dmem_req_bits_addr_msb_T_2; // @[RocketCore.scala 990:29]
  wire  msb_2; // @[RocketCore.scala 990:18]
  wire [38:0] io_dmem_req_bits_addr_lo; // @[RocketCore.scala 991:16]
  wire  _io_dmem_s1_kill_T; // @[RocketCore.scala 848:35]
  wire  _unpause_T_1; // @[RocketCore.scala 861:62]
  wire  _unpause_T_2; // @[RocketCore.scala 861:68]
  wire  _unpause_T_3; // @[RocketCore.scala 861:92]
  wire  unpause; // @[RocketCore.scala 861:116]
  wire  coreMonitorBundle_valid; // @[RocketCore.scala 889:52]
  wire  coreMonitorBundle_wrenx; // @[RocketCore.scala 891:37]
  wire [5:0] _GEN_251; // @[RocketCore.scala 912:95]
  wire [5:0] _T_142; // @[RocketCore.scala 912:95]
  wire  _T_145; // @[RocketCore.scala 914:28]
  wire  _T_146; // @[RocketCore.scala 914:22]
  wire  _T_147; // @[RocketCore.scala 914:40]
  wire  _T_153; // @[RocketCore.scala 917:40]
  wire  _T_159; // @[RocketCore.scala 925:18]
  wire  _GEN_254; // @[RocketCore.scala 912:16]
  wire  _GEN_256; // @[RocketCore.scala 915:16]
  wire  _GEN_257; // @[RocketCore.scala 915:16]
  wire  _GEN_261; // @[RocketCore.scala 918:16]
  wire  _GEN_262; // @[RocketCore.scala 918:16]
  wire  _GEN_268; // @[RocketCore.scala 921:16]
  reg [19:0] Rocket_state; // @[Register tracking Rocket state]
  reg [31:0] _RAND_94;
  reg  Rocket_cov [0:1048575]; // @[Coverage map for Rocket]
  reg [31:0] _RAND_95;
  wire  Rocket_cov_read_data; // @[Coverage map for Rocket]
  wire [19:0] Rocket_cov_read_addr; // @[Coverage map for Rocket]
  wire  Rocket_cov_write_data; // @[Coverage map for Rocket]
  wire [19:0] Rocket_cov_write_addr; // @[Coverage map for Rocket]
  wire  Rocket_cov_write_mask; // @[Coverage map for Rocket]
  wire  Rocket_cov_write_en; // @[Coverage map for Rocket]
  reg [29:0] Rocket_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_96;
  wire  mux_cond_0;
  wire  mux_cond_1;
  wire  mux_cond_2;
  wire  mux_cond_3;
  wire  mux_cond_4;
  wire  mux_cond_5;
  wire [10:0] ex_ctrl_wfd_shl;
  wire [19:0] ex_ctrl_wfd_pad;
  wire [15:0] ex_ctrl_fp_shl;
  wire [19:0] ex_ctrl_fp_pad;
  wire [15:0] mem_ctrl_jalr_shl;
  wire [19:0] mem_ctrl_jalr_pad;
  wire [11:0] wb_ctrl_mem_shl;
  wire [19:0] wb_ctrl_mem_pad;
  wire [6:0] ex_ctrl_wxd_shl;
  wire [19:0] ex_ctrl_wxd_pad;
  wire [19:0] ex_ctrl_mem_shl;
  wire [19:0] ex_ctrl_mem_pad;
  wire [19:0] ex_ctrl_sel_alu1_shl;
  wire [19:0] ex_ctrl_sel_alu1_pad;
  wire [11:0] mem_reg_replay_shl;
  wire [19:0] mem_reg_replay_pad;
  wire [16:0] blocked_shl;
  wire [19:0] blocked_pad;
  wire [2:0] wb_ctrl_div_shl;
  wire [19:0] wb_ctrl_div_pad;
  wire [15:0] wb_reg_flush_pipe_shl;
  wire [19:0] wb_reg_flush_pipe_pad;
  wire [11:0] mem_ctrl_jal_shl;
  wire [19:0] mem_ctrl_jal_pad;
  wire [9:0] ex_ctrl_sel_imm_shl;
  wire [19:0] ex_ctrl_sel_imm_pad;
  wire [8:0] wb_ctrl_wfd_shl;
  wire [19:0] wb_ctrl_wfd_pad;
  wire [19:0] mem_reg_slow_bypass_shl;
  wire [19:0] mem_reg_slow_bypass_pad;
  wire [16:0] mem_reg_sfence_shl;
  wire [19:0] mem_reg_sfence_pad;
  wire [2:0] wb_reg_xcpt_shl;
  wire [19:0] wb_reg_xcpt_pad;
  wire [15:0] id_reg_pause_shl;
  wire [19:0] id_reg_pause_pad;
  wire [8:0] ex_reg_rvc_shl;
  wire [19:0] ex_reg_rvc_pad;
  wire [3:0] wb_reg_valid_shl;
  wire [19:0] wb_reg_valid_pad;
  wire [13:0] mem_br_taken_shl;
  wire [19:0] mem_br_taken_pad;
  wire [18:0] mem_reg_flush_pipe_shl;
  wire [19:0] mem_reg_flush_pipe_pad;
  wire [17:0] ex_ctrl_div_shl;
  wire [19:0] ex_ctrl_div_pad;
  wire [15:0] mem_ctrl_fp_shl;
  wire [19:0] mem_ctrl_fp_pad;
  wire [5:0] mem_reg_xcpt_shl;
  wire [19:0] mem_reg_xcpt_pad;
  wire [14:0] mem_ctrl_wxd_shl;
  wire [19:0] mem_ctrl_wxd_pad;
  wire [8:0] mem_ctrl_mem_shl;
  wire [19:0] mem_ctrl_mem_pad;
  wire [16:0] ex_reg_mem_size_shl;
  wire [19:0] ex_reg_mem_size_pad;
  wire [8:0] ex_ctrl_sel_alu2_shl;
  wire [19:0] ex_ctrl_sel_alu2_pad;
  wire [2:0] ex_ctrl_rxs2_shl;
  wire [19:0] ex_ctrl_rxs2_pad;
  wire [3:0] ex_ctrl_jalr_shl;
  wire [19:0] ex_ctrl_jalr_pad;
  wire [4:0] ex_reg_replay_shl;
  wire [19:0] ex_reg_replay_pad;
  wire [3:0] ex_reg_valid_shl;
  wire [19:0] ex_reg_valid_pad;
  wire [6:0] mem_reg_valid_shl;
  wire [19:0] mem_reg_valid_pad;
  wire  mem_reg_rvc_shl;
  wire [19:0] mem_reg_rvc_pad;
  wire  mem_ctrl_wfd_shl;
  wire [19:0] mem_ctrl_wfd_pad;
  wire [11:0] id_reg_fence_shl;
  wire [19:0] id_reg_fence_pad;
  wire [8:0] mem_reg_load_shl;
  wire [19:0] mem_reg_load_pad;
  wire [18:0] wb_ctrl_wxd_shl;
  wire [19:0] wb_ctrl_wxd_pad;
  wire [1:0] wb_reg_replay_shl;
  wire [19:0] wb_reg_replay_pad;
  wire [10:0] ex_reg_xcpt_interrupt_shl;
  wire [19:0] ex_reg_xcpt_interrupt_pad;
  wire [6:0] mem_ctrl_branch_shl;
  wire [19:0] mem_ctrl_branch_pad;
  wire [1:0] mem_reg_xcpt_interrupt_shl;
  wire [19:0] mem_reg_xcpt_interrupt_pad;
  wire [4:0] mem_reg_store_shl;
  wire [19:0] mem_reg_store_pad;
  wire [5:0] mem_ctrl_div_shl;
  wire [19:0] mem_ctrl_div_pad;
  wire [17:0] mux_cond_0_shl;
  wire [19:0] mux_cond_0_pad;
  wire [8:0] mux_cond_1_shl;
  wire [19:0] mux_cond_1_pad;
  wire [15:0] mux_cond_2_shl;
  wire [19:0] mux_cond_2_pad;
  wire [4:0] mux_cond_3_shl;
  wire [19:0] mux_cond_3_pad;
  wire [9:0] mux_cond_4_shl;
  wire [19:0] mux_cond_4_pad;
  wire [17:0] mux_cond_5_shl;
  wire [19:0] mux_cond_5_pad;
  wire [12:0] ex_reg_rs_lsb_0_shl;
  wire [19:0] ex_reg_rs_lsb_0_pad;
  wire [12:0] ex_reg_rs_lsb_1_shl;
  wire [19:0] ex_reg_rs_lsb_1_pad;
  wire [10:0] ex_reg_rs_bypass_0_shl;
  wire [19:0] ex_reg_rs_bypass_0_pad;
  wire [10:0] ex_reg_rs_bypass_1_shl;
  wire [19:0] ex_reg_rs_bypass_1_pad;
  wire [19:0] Rocket_xor32;
  wire [19:0] Rocket_xor15;
  wire [19:0] Rocket_xor34;
  wire [19:0] Rocket_xor16;
  wire [19:0] Rocket_xor7;
  wire [19:0] Rocket_xor36;
  wire [19:0] Rocket_xor17;
  wire [19:0] Rocket_xor37;
  wire [19:0] Rocket_xor38;
  wire [19:0] Rocket_xor18;
  wire [19:0] Rocket_xor8;
  wire [19:0] Rocket_xor3;
  wire [19:0] Rocket_xor40;
  wire [19:0] Rocket_xor19;
  wire [19:0] Rocket_xor41;
  wire [19:0] Rocket_xor42;
  wire [19:0] Rocket_xor20;
  wire [19:0] Rocket_xor9;
  wire [19:0] Rocket_xor44;
  wire [19:0] Rocket_xor21;
  wire [19:0] Rocket_xor45;
  wire [19:0] Rocket_xor46;
  wire [19:0] Rocket_xor22;
  wire [19:0] Rocket_xor10;
  wire [19:0] Rocket_xor4;
  wire [19:0] Rocket_xor1;
  wire [19:0] Rocket_xor48;
  wire [19:0] Rocket_xor23;
  wire [19:0] Rocket_xor49;
  wire [19:0] Rocket_xor50;
  wire [19:0] Rocket_xor24;
  wire [19:0] Rocket_xor11;
  wire [19:0] Rocket_xor52;
  wire [19:0] Rocket_xor25;
  wire [19:0] Rocket_xor53;
  wire [19:0] Rocket_xor54;
  wire [19:0] Rocket_xor26;
  wire [19:0] Rocket_xor12;
  wire [19:0] Rocket_xor5;
  wire [19:0] Rocket_xor56;
  wire [19:0] Rocket_xor27;
  wire [19:0] Rocket_xor57;
  wire [19:0] Rocket_xor58;
  wire [19:0] Rocket_xor28;
  wire [19:0] Rocket_xor13;
  wire [19:0] Rocket_xor60;
  wire [19:0] Rocket_xor29;
  wire [19:0] Rocket_xor61;
  wire [19:0] Rocket_xor62;
  wire [19:0] Rocket_xor30;
  wire [19:0] Rocket_xor14;
  wire [19:0] Rocket_xor6;
  wire [19:0] Rocket_xor2;
  wire [19:0] Rocket_xor0;
  wire [29:0] PlusArgTimeout_sum;
  wire [29:0] csr_sum;
  wire [29:0] bpu_sum;
  wire [29:0] ibuf_sum;
  wire [29:0] div_sum;
  wire [29:0] alu_sum;
  wire  alu_metaAssert_wire;
  wire  div_metaAssert_wire;
  wire  bpu_metaAssert_wire;
  wire  PlusArgTimeout_metaAssert_wire;
  wire  ibuf_metaAssert_wire;
  wire  csr_metaAssert_wire;
  wire  Rocket_or4;
  wire  Rocket_or1;
  wire  Rocket_or6;
  wire  Rocket_or2;
  wire  Rocket_or0;
  reg  Rocket_metaAssert;
  reg [31:0] _RAND_97;
  IBuf ibuf ( // @[RocketCore.scala 254:20]
    .clock(ibuf_clock),
    .reset(ibuf_reset),
    .io_imem_ready(ibuf_io_imem_ready),
    .io_imem_valid(ibuf_io_imem_valid),
    .io_imem_bits_btb_taken(ibuf_io_imem_bits_btb_taken),
    .io_imem_bits_btb_bridx(ibuf_io_imem_bits_btb_bridx),
    .io_imem_bits_btb_entry(ibuf_io_imem_bits_btb_entry),
    .io_imem_bits_btb_bht_history(ibuf_io_imem_bits_btb_bht_history),
    .io_imem_bits_pc(ibuf_io_imem_bits_pc),
    .io_imem_bits_data(ibuf_io_imem_bits_data),
    .io_imem_bits_xcpt_pf_inst(ibuf_io_imem_bits_xcpt_pf_inst),
    .io_imem_bits_xcpt_ae_inst(ibuf_io_imem_bits_xcpt_ae_inst),
    .io_imem_bits_replay(ibuf_io_imem_bits_replay),
    .io_kill(ibuf_io_kill),
    .io_pc(ibuf_io_pc),
    .io_btb_resp_entry(ibuf_io_btb_resp_entry),
    .io_btb_resp_bht_history(ibuf_io_btb_resp_bht_history),
    .io_inst_0_ready(ibuf_io_inst_0_ready),
    .io_inst_0_valid(ibuf_io_inst_0_valid),
    .io_inst_0_bits_xcpt0_pf_inst(ibuf_io_inst_0_bits_xcpt0_pf_inst),
    .io_inst_0_bits_xcpt0_ae_inst(ibuf_io_inst_0_bits_xcpt0_ae_inst),
    .io_inst_0_bits_xcpt1_pf_inst(ibuf_io_inst_0_bits_xcpt1_pf_inst),
    .io_inst_0_bits_xcpt1_ae_inst(ibuf_io_inst_0_bits_xcpt1_ae_inst),
    .io_inst_0_bits_replay(ibuf_io_inst_0_bits_replay),
    .io_inst_0_bits_rvc(ibuf_io_inst_0_bits_rvc),
    .io_inst_0_bits_inst_bits(ibuf_io_inst_0_bits_inst_bits),
    .io_inst_0_bits_inst_rd(ibuf_io_inst_0_bits_inst_rd),
    .io_inst_0_bits_inst_rs1(ibuf_io_inst_0_bits_inst_rs1),
    .io_inst_0_bits_inst_rs2(ibuf_io_inst_0_bits_inst_rs2),
    .io_inst_0_bits_inst_rs3(ibuf_io_inst_0_bits_inst_rs3),
    .io_inst_0_bits_raw(ibuf_io_inst_0_bits_raw),
    .io_covSum(ibuf_io_covSum),
    .metaAssert(ibuf_metaAssert),
    .metaReset(ibuf_metaReset)
  );
  CSRFile csr ( // @[RocketCore.scala 282:19]
    .clock(csr_clock),
    .reset(csr_reset),
    .io_ungated_clock(csr_io_ungated_clock),
    .io_interrupts_debug(csr_io_interrupts_debug),
    .io_interrupts_mtip(csr_io_interrupts_mtip),
    .io_interrupts_msip(csr_io_interrupts_msip),
    .io_interrupts_meip(csr_io_interrupts_meip),
    .io_interrupts_seip(csr_io_interrupts_seip),
    .io_hartid(csr_io_hartid),
    .io_rw_addr(csr_io_rw_addr),
    .io_rw_cmd(csr_io_rw_cmd),
    .io_rw_rdata(csr_io_rw_rdata),
    .io_rw_wdata(csr_io_rw_wdata),
    .io_decode_0_csr(csr_io_decode_0_csr),
    .io_decode_0_fp_illegal(csr_io_decode_0_fp_illegal),
    .io_decode_0_fp_csr(csr_io_decode_0_fp_csr),
    .io_decode_0_read_illegal(csr_io_decode_0_read_illegal),
    .io_decode_0_write_illegal(csr_io_decode_0_write_illegal),
    .io_decode_0_write_flush(csr_io_decode_0_write_flush),
    .io_decode_0_system_illegal(csr_io_decode_0_system_illegal),
    .io_csr_stall(csr_io_csr_stall),
    .io_eret(csr_io_eret),
    .io_singleStep(csr_io_singleStep),
    .io_status_debug(csr_io_status_debug),
    .io_status_cease(csr_io_status_cease),
    .io_status_wfi(csr_io_status_wfi),
    .io_status_isa(csr_io_status_isa),
    .io_status_dprv(csr_io_status_dprv),
    .io_status_prv(csr_io_status_prv),
    .io_status_sd(csr_io_status_sd),
    .io_status_zero2(csr_io_status_zero2),
    .io_status_sxl(csr_io_status_sxl),
    .io_status_uxl(csr_io_status_uxl),
    .io_status_sd_rv32(csr_io_status_sd_rv32),
    .io_status_zero1(csr_io_status_zero1),
    .io_status_tsr(csr_io_status_tsr),
    .io_status_tw(csr_io_status_tw),
    .io_status_tvm(csr_io_status_tvm),
    .io_status_mxr(csr_io_status_mxr),
    .io_status_sum(csr_io_status_sum),
    .io_status_mprv(csr_io_status_mprv),
    .io_status_xs(csr_io_status_xs),
    .io_status_fs(csr_io_status_fs),
    .io_status_mpp(csr_io_status_mpp),
    .io_status_vs(csr_io_status_vs),
    .io_status_spp(csr_io_status_spp),
    .io_status_mpie(csr_io_status_mpie),
    .io_status_hpie(csr_io_status_hpie),
    .io_status_spie(csr_io_status_spie),
    .io_status_upie(csr_io_status_upie),
    .io_status_mie(csr_io_status_mie),
    .io_status_hie(csr_io_status_hie),
    .io_status_sie(csr_io_status_sie),
    .io_status_uie(csr_io_status_uie),
    .io_ptbr_mode(csr_io_ptbr_mode),
    .io_ptbr_ppn(csr_io_ptbr_ppn),
    .io_evec(csr_io_evec),
    .io_exception(csr_io_exception),
    .io_retire(csr_io_retire),
    .io_cause(csr_io_cause),
    .io_pc(csr_io_pc),
    .io_tval(csr_io_tval),
    .io_time(csr_io_time),
    .io_fcsr_rm(csr_io_fcsr_rm),
    .io_fcsr_flags_valid(csr_io_fcsr_flags_valid),
    .io_fcsr_flags_bits(csr_io_fcsr_flags_bits),
    .io_interrupt(csr_io_interrupt),
    .io_interrupt_cause(csr_io_interrupt_cause),
    .io_bp_0_control_action(csr_io_bp_0_control_action),
    .io_bp_0_control_tmatch(csr_io_bp_0_control_tmatch),
    .io_bp_0_control_m(csr_io_bp_0_control_m),
    .io_bp_0_control_s(csr_io_bp_0_control_s),
    .io_bp_0_control_u(csr_io_bp_0_control_u),
    .io_bp_0_control_x(csr_io_bp_0_control_x),
    .io_bp_0_control_w(csr_io_bp_0_control_w),
    .io_bp_0_control_r(csr_io_bp_0_control_r),
    .io_bp_0_address(csr_io_bp_0_address),
    .io_pmp_0_cfg_l(csr_io_pmp_0_cfg_l),
    .io_pmp_0_cfg_a(csr_io_pmp_0_cfg_a),
    .io_pmp_0_cfg_x(csr_io_pmp_0_cfg_x),
    .io_pmp_0_cfg_w(csr_io_pmp_0_cfg_w),
    .io_pmp_0_cfg_r(csr_io_pmp_0_cfg_r),
    .io_pmp_0_addr(csr_io_pmp_0_addr),
    .io_pmp_0_mask(csr_io_pmp_0_mask),
    .io_pmp_1_cfg_l(csr_io_pmp_1_cfg_l),
    .io_pmp_1_cfg_a(csr_io_pmp_1_cfg_a),
    .io_pmp_1_cfg_x(csr_io_pmp_1_cfg_x),
    .io_pmp_1_cfg_w(csr_io_pmp_1_cfg_w),
    .io_pmp_1_cfg_r(csr_io_pmp_1_cfg_r),
    .io_pmp_1_addr(csr_io_pmp_1_addr),
    .io_pmp_1_mask(csr_io_pmp_1_mask),
    .io_pmp_2_cfg_l(csr_io_pmp_2_cfg_l),
    .io_pmp_2_cfg_a(csr_io_pmp_2_cfg_a),
    .io_pmp_2_cfg_x(csr_io_pmp_2_cfg_x),
    .io_pmp_2_cfg_w(csr_io_pmp_2_cfg_w),
    .io_pmp_2_cfg_r(csr_io_pmp_2_cfg_r),
    .io_pmp_2_addr(csr_io_pmp_2_addr),
    .io_pmp_2_mask(csr_io_pmp_2_mask),
    .io_pmp_3_cfg_l(csr_io_pmp_3_cfg_l),
    .io_pmp_3_cfg_a(csr_io_pmp_3_cfg_a),
    .io_pmp_3_cfg_x(csr_io_pmp_3_cfg_x),
    .io_pmp_3_cfg_w(csr_io_pmp_3_cfg_w),
    .io_pmp_3_cfg_r(csr_io_pmp_3_cfg_r),
    .io_pmp_3_addr(csr_io_pmp_3_addr),
    .io_pmp_3_mask(csr_io_pmp_3_mask),
    .io_pmp_4_cfg_l(csr_io_pmp_4_cfg_l),
    .io_pmp_4_cfg_a(csr_io_pmp_4_cfg_a),
    .io_pmp_4_cfg_x(csr_io_pmp_4_cfg_x),
    .io_pmp_4_cfg_w(csr_io_pmp_4_cfg_w),
    .io_pmp_4_cfg_r(csr_io_pmp_4_cfg_r),
    .io_pmp_4_addr(csr_io_pmp_4_addr),
    .io_pmp_4_mask(csr_io_pmp_4_mask),
    .io_pmp_5_cfg_l(csr_io_pmp_5_cfg_l),
    .io_pmp_5_cfg_a(csr_io_pmp_5_cfg_a),
    .io_pmp_5_cfg_x(csr_io_pmp_5_cfg_x),
    .io_pmp_5_cfg_w(csr_io_pmp_5_cfg_w),
    .io_pmp_5_cfg_r(csr_io_pmp_5_cfg_r),
    .io_pmp_5_addr(csr_io_pmp_5_addr),
    .io_pmp_5_mask(csr_io_pmp_5_mask),
    .io_pmp_6_cfg_l(csr_io_pmp_6_cfg_l),
    .io_pmp_6_cfg_a(csr_io_pmp_6_cfg_a),
    .io_pmp_6_cfg_x(csr_io_pmp_6_cfg_x),
    .io_pmp_6_cfg_w(csr_io_pmp_6_cfg_w),
    .io_pmp_6_cfg_r(csr_io_pmp_6_cfg_r),
    .io_pmp_6_addr(csr_io_pmp_6_addr),
    .io_pmp_6_mask(csr_io_pmp_6_mask),
    .io_pmp_7_cfg_l(csr_io_pmp_7_cfg_l),
    .io_pmp_7_cfg_a(csr_io_pmp_7_cfg_a),
    .io_pmp_7_cfg_x(csr_io_pmp_7_cfg_x),
    .io_pmp_7_cfg_w(csr_io_pmp_7_cfg_w),
    .io_pmp_7_cfg_r(csr_io_pmp_7_cfg_r),
    .io_pmp_7_addr(csr_io_pmp_7_addr),
    .io_pmp_7_mask(csr_io_pmp_7_mask),
    .io_inhibit_cycle(csr_io_inhibit_cycle),
    .io_inst_0(csr_io_inst_0),
    .io_trace_0_valid(csr_io_trace_0_valid),
    .io_trace_0_iaddr(csr_io_trace_0_iaddr),
    .io_trace_0_insn(csr_io_trace_0_insn),
    .io_trace_0_priv(csr_io_trace_0_priv),
    .io_trace_0_exception(csr_io_trace_0_exception),
    .io_trace_0_interrupt(csr_io_trace_0_interrupt),
    .io_trace_0_cause(csr_io_trace_0_cause),
    .io_trace_0_tval(csr_io_trace_0_tval),
    .io_customCSRs_0_value(csr_io_customCSRs_0_value),
    .io_covSum(csr_io_covSum),
    .metaAssert(csr_metaAssert),
    .metaReset(csr_metaReset)
  );
  BreakpointUnit bpu ( // @[RocketCore.scala 323:19]
    .io_status_debug(bpu_io_status_debug),
    .io_status_prv(bpu_io_status_prv),
    .io_bp_0_control_action(bpu_io_bp_0_control_action),
    .io_bp_0_control_tmatch(bpu_io_bp_0_control_tmatch),
    .io_bp_0_control_m(bpu_io_bp_0_control_m),
    .io_bp_0_control_s(bpu_io_bp_0_control_s),
    .io_bp_0_control_u(bpu_io_bp_0_control_u),
    .io_bp_0_control_x(bpu_io_bp_0_control_x),
    .io_bp_0_control_w(bpu_io_bp_0_control_w),
    .io_bp_0_control_r(bpu_io_bp_0_control_r),
    .io_bp_0_address(bpu_io_bp_0_address),
    .io_pc(bpu_io_pc),
    .io_ea(bpu_io_ea),
    .io_xcpt_if(bpu_io_xcpt_if),
    .io_xcpt_ld(bpu_io_xcpt_ld),
    .io_xcpt_st(bpu_io_xcpt_st),
    .io_debug_if(bpu_io_debug_if),
    .io_debug_ld(bpu_io_debug_ld),
    .io_debug_st(bpu_io_debug_st),
    .io_covSum(bpu_io_covSum),
    .metaAssert(bpu_metaAssert)
  );
  ALU alu ( // @[RocketCore.scala 385:19]
    .io_dw(alu_io_dw),
    .io_fn(alu_io_fn),
    .io_in2(alu_io_in2),
    .io_in1(alu_io_in1),
    .io_out(alu_io_out),
    .io_adder_out(alu_io_adder_out),
    .io_cmp_out(alu_io_cmp_out),
    .io_covSum(alu_io_covSum),
    .metaAssert(alu_metaAssert)
  );
  MulDiv div ( // @[RocketCore.scala 409:19]
    .clock(div_clock),
    .reset(div_reset),
    .io_req_ready(div_io_req_ready),
    .io_req_valid(div_io_req_valid),
    .io_req_bits_fn(div_io_req_bits_fn),
    .io_req_bits_dw(div_io_req_bits_dw),
    .io_req_bits_in1(div_io_req_bits_in1),
    .io_req_bits_in2(div_io_req_bits_in2),
    .io_req_bits_tag(div_io_req_bits_tag),
    .io_kill(div_io_kill),
    .io_resp_ready(div_io_resp_ready),
    .io_resp_valid(div_io_resp_valid),
    .io_resp_bits_data(div_io_resp_bits_data),
    .io_resp_bits_tag(div_io_resp_bits_tag),
    .io_covSum(div_io_covSum),
    .metaAssert(div_metaAssert),
    .metaReset(div_metaReset)
  );
  PlusArgTimeout PlusArgTimeout ( // @[PlusArg.scala 89:11]
    .clock(PlusArgTimeout_clock),
    .reset(PlusArgTimeout_reset),
    .io_count(PlusArgTimeout_io_count),
    .io_covSum(PlusArgTimeout_io_covSum),
    .metaAssert(PlusArgTimeout_metaAssert),
    .metaReset(PlusArgTimeout_metaReset)
  );
  assign rf_id_rs_MPORT_addr = ~id_raddr1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign rf_id_rs_MPORT_data = rf[rf_id_rs_MPORT_addr]; // @[RocketCore.scala 1015:15]
  `else
  assign rf_id_rs_MPORT_data = rf_id_rs_MPORT_addr >= 5'h1f ? _RAND_1[63:0] : rf[rf_id_rs_MPORT_addr]; // @[RocketCore.scala 1015:15]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign rf_id_rs_MPORT_1_addr = ~id_raddr2;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign rf_id_rs_MPORT_1_data = rf[rf_id_rs_MPORT_1_addr]; // @[RocketCore.scala 1015:15]
  `else
  assign rf_id_rs_MPORT_1_data = rf_id_rs_MPORT_1_addr >= 5'h1f ? _RAND_2[63:0] : rf[rf_id_rs_MPORT_1_addr]; // @[RocketCore.scala 1015:15]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign rf_MPORT_data = _rf_wdata_T ? io_dmem_resp_bits_data : _rf_wdata_T_5;
  assign rf_MPORT_addr = ~rf_waddr;
  assign rf_MPORT_mask = 1'h1;
  assign rf_MPORT_en = rf_wen & _T_118;
  assign replay_wb_common = io_dmem_s2_nack | wb_reg_replay; // @[RocketCore.scala 637:42]
  assign _T_83 = wb_reg_valid & wb_ctrl_mem; // @[RocketCore.scala 615:19]
  assign _T_84 = _T_83 & io_dmem_s2_xcpt_ma_st; // @[RocketCore.scala 615:34]
  assign _T_95 = wb_reg_xcpt | _T_84; // @[RocketCore.scala 975:26]
  assign _T_86 = _T_83 & io_dmem_s2_xcpt_ma_ld; // @[RocketCore.scala 616:34]
  assign _T_96 = _T_95 | _T_86; // @[RocketCore.scala 975:26]
  assign _T_88 = _T_83 & io_dmem_s2_xcpt_pf_st; // @[RocketCore.scala 617:34]
  assign _T_97 = _T_96 | _T_88; // @[RocketCore.scala 975:26]
  assign _T_90 = _T_83 & io_dmem_s2_xcpt_pf_ld; // @[RocketCore.scala 618:34]
  assign _T_98 = _T_97 | _T_90; // @[RocketCore.scala 975:26]
  assign _T_92 = _T_83 & io_dmem_s2_xcpt_ae_st; // @[RocketCore.scala 619:34]
  assign _T_99 = _T_98 | _T_92; // @[RocketCore.scala 975:26]
  assign _T_94 = _T_83 & io_dmem_s2_xcpt_ae_ld; // @[RocketCore.scala 620:34]
  assign wb_xcpt = _T_99 | _T_94; // @[RocketCore.scala 975:26]
  assign _take_pc_wb_T = replay_wb_common | wb_xcpt; // @[RocketCore.scala 640:27]
  assign _take_pc_wb_T_1 = _take_pc_wb_T | csr_io_eret; // @[RocketCore.scala 640:38]
  assign take_pc_wb = _take_pc_wb_T_1 | wb_reg_flush_pipe; // @[RocketCore.scala 640:53]
  assign _ex_pc_valid_T = ex_reg_valid | ex_reg_replay; // @[RocketCore.scala 490:34]
  assign ex_pc_valid = _ex_pc_valid_T | ex_reg_xcpt_interrupt; // @[RocketCore.scala 490:51]
  assign _mem_npc_T = mem_ctrl_jalr | mem_reg_sfence; // @[RocketCore.scala 513:36]
  assign a = mem_reg_wdata[63:39]; // @[RocketCore.scala 989:23]
  assign _mem_npc_msb_T = $signed(a) == 25'sh0; // @[RocketCore.scala 990:21]
  assign _mem_npc_msb_T_1 = $signed(a) == -25'sh1; // @[RocketCore.scala 990:34]
  assign _mem_npc_msb_T_2 = _mem_npc_msb_T | _mem_npc_msb_T_1; // @[RocketCore.scala 990:29]
  assign msb = _mem_npc_msb_T_2 ? mem_reg_wdata[39] : ~mem_reg_wdata[38]; // @[RocketCore.scala 990:18]
  assign mem_npc_lo = mem_reg_wdata[38:0]; // @[RocketCore.scala 991:16]
  assign _mem_npc_T_2 = {msb,mem_npc_lo}; // @[RocketCore.scala 513:106]
  assign _mem_br_target_T_1 = mem_ctrl_branch & mem_br_taken; // @[RocketCore.scala 510:25]
  assign mem_br_target_sign = mem_reg_inst[31]; // @[RocketCore.scala 1037:53]
  assign mem_br_target_hi_hi_hi = mem_reg_inst[31]; // @[Cat.scala 30:58]
  assign mem_br_target_hi_hi_lo = {11{mem_br_target_sign}}; // @[Cat.scala 30:58]
  assign mem_br_target_hi_lo_hi = {8{mem_br_target_sign}}; // @[Cat.scala 30:58]
  assign mem_br_target_hi_lo_lo = mem_reg_inst[7]; // @[Cat.scala 30:58]
  assign mem_br_target_lo_hi_hi = mem_reg_inst[30:25]; // @[RocketCore.scala 1043:66]
  assign mem_br_target_lo_hi_lo = mem_reg_inst[11:8]; // @[RocketCore.scala 1045:57]
  assign _mem_br_target_T_3 = {mem_br_target_hi_hi_hi,mem_br_target_hi_hi_lo,mem_br_target_hi_lo_hi,mem_br_target_hi_lo_lo,mem_br_target_lo_hi_hi,mem_br_target_lo_hi_lo,1'h0}; // @[RocketCore.scala 1051:53]
  assign mem_br_target_hi_lo_hi_1 = mem_reg_inst[19:12]; // @[Cat.scala 30:58]
  assign mem_br_target_hi_lo_lo_1 = mem_reg_inst[20]; // @[Cat.scala 30:58]
  assign _mem_br_target_T_5 = {mem_br_target_hi_hi_hi,mem_br_target_hi_hi_lo,mem_br_target_hi_lo_hi_1,mem_br_target_hi_lo_lo_1,mem_br_target_lo_hi_hi,mem_reg_inst[24:21],1'h0}; // @[RocketCore.scala 1051:53]
  assign _mem_br_target_T_6 = mem_reg_rvc ? $signed(4'sh2) : $signed(4'sh4); // @[RocketCore.scala 512:8]
  assign _mem_br_target_T_7 = mem_ctrl_jal ? $signed(_mem_br_target_T_5) : $signed({{28{_mem_br_target_T_6[3]}},_mem_br_target_T_6}); // @[RocketCore.scala 511:8]
  assign _mem_br_target_T_8 = _mem_br_target_T_1 ? $signed(_mem_br_target_T_3) : $signed(_mem_br_target_T_7); // @[RocketCore.scala 510:8]
  assign _GEN_248 = {{8{_mem_br_target_T_8[31]}},_mem_br_target_T_8}; // @[RocketCore.scala 509:41]
  assign mem_br_target = $signed(mem_reg_pc) + $signed(_GEN_248); // @[RocketCore.scala 509:41]
  assign _mem_npc_T_3 = _mem_npc_T ? $signed(_mem_npc_T_2) : $signed(mem_br_target); // @[RocketCore.scala 513:21]
  assign mem_npc = $signed(_mem_npc_T_3) & -40'sh2; // @[RocketCore.scala 513:141]
  assign _mem_wrong_npc_T = mem_npc != ex_reg_pc; // @[RocketCore.scala 515:30]
  assign _mem_wrong_npc_T_1 = ibuf_io_inst_0_valid | ibuf_io_imem_valid; // @[RocketCore.scala 516:31]
  assign _mem_wrong_npc_T_2 = mem_npc != ibuf_io_pc; // @[RocketCore.scala 516:62]
  assign _mem_wrong_npc_T_3 = _mem_wrong_npc_T_1 ? _mem_wrong_npc_T_2 : 1'h1; // @[RocketCore.scala 516:8]
  assign mem_wrong_npc = ex_pc_valid ? _mem_wrong_npc_T : _mem_wrong_npc_T_3; // @[RocketCore.scala 515:8]
  assign _take_pc_mem_T = mem_wrong_npc | mem_reg_sfence; // @[RocketCore.scala 523:54]
  assign take_pc_mem = mem_reg_valid & _take_pc_mem_T; // @[RocketCore.scala 523:32]
  assign take_pc_mem_wb = take_pc_wb | take_pc_mem; // @[RocketCore.scala 250:35]
  assign _id_ctrl_decoder_bit_T = ibuf_io_inst_0_bits_inst_bits & 32'hfe00707f; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_bit_T_1 = _id_ctrl_decoder_bit_T == 32'h2000033; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_3 = _id_ctrl_decoder_bit_T == 32'h2001033; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_5 = _id_ctrl_decoder_bit_T == 32'h2003033; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_7 = _id_ctrl_decoder_bit_T == 32'h2002033; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_9 = _id_ctrl_decoder_bit_T == 32'h2004033; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_11 = _id_ctrl_decoder_bit_T == 32'h2005033; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_13 = _id_ctrl_decoder_bit_T == 32'h2006033; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_15 = _id_ctrl_decoder_bit_T == 32'h2007033; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_17 = _id_ctrl_decoder_bit_T == 32'h200003b; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_19 = _id_ctrl_decoder_bit_T == 32'h200403b; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_21 = _id_ctrl_decoder_bit_T == 32'h200503b; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_23 = _id_ctrl_decoder_bit_T == 32'h200603b; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_25 = _id_ctrl_decoder_bit_T == 32'h200703b; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_26 = ibuf_io_inst_0_bits_inst_bits & 32'hf800707f; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_bit_T_27 = _id_ctrl_decoder_bit_T_26 == 32'h202f; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_29 = _id_ctrl_decoder_bit_T_26 == 32'h2000202f; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_31 = _id_ctrl_decoder_bit_T_26 == 32'h800202f; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_33 = _id_ctrl_decoder_bit_T_26 == 32'h6000202f; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_35 = _id_ctrl_decoder_bit_T_26 == 32'h4000202f; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_37 = _id_ctrl_decoder_bit_T_26 == 32'h8000202f; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_39 = _id_ctrl_decoder_bit_T_26 == 32'hc000202f; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_41 = _id_ctrl_decoder_bit_T_26 == 32'ha000202f; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_43 = _id_ctrl_decoder_bit_T_26 == 32'he000202f; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_44 = ibuf_io_inst_0_bits_inst_bits & 32'hf9f0707f; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_bit_T_45 = _id_ctrl_decoder_bit_T_44 == 32'h1000202f; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_47 = _id_ctrl_decoder_bit_T_26 == 32'h1800202f; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_49 = _id_ctrl_decoder_bit_T_26 == 32'h302f; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_51 = _id_ctrl_decoder_bit_T_26 == 32'h800302f; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_53 = _id_ctrl_decoder_bit_T_26 == 32'h2000302f; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_55 = _id_ctrl_decoder_bit_T_26 == 32'h6000302f; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_57 = _id_ctrl_decoder_bit_T_26 == 32'h4000302f; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_59 = _id_ctrl_decoder_bit_T_26 == 32'h8000302f; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_61 = _id_ctrl_decoder_bit_T_26 == 32'hc000302f; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_63 = _id_ctrl_decoder_bit_T_26 == 32'ha000302f; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_65 = _id_ctrl_decoder_bit_T_26 == 32'he000302f; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_67 = _id_ctrl_decoder_bit_T_44 == 32'h1000302f; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_69 = _id_ctrl_decoder_bit_T_26 == 32'h1800302f; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_71 = _id_ctrl_decoder_bit_T == 32'h20000053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_73 = _id_ctrl_decoder_bit_T == 32'h20002053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_75 = _id_ctrl_decoder_bit_T == 32'h20001053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_77 = _id_ctrl_decoder_bit_T == 32'h28000053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_79 = _id_ctrl_decoder_bit_T == 32'h28001053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_80 = ibuf_io_inst_0_bits_inst_bits & 32'hfe00007f; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_bit_T_81 = _id_ctrl_decoder_bit_T_80 == 32'h53; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_83 = _id_ctrl_decoder_bit_T_80 == 32'h8000053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_85 = _id_ctrl_decoder_bit_T_80 == 32'h10000053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_86 = ibuf_io_inst_0_bits_inst_bits & 32'h600007f; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_bit_T_87 = _id_ctrl_decoder_bit_T_86 == 32'h43; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_89 = _id_ctrl_decoder_bit_T_86 == 32'h47; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_91 = _id_ctrl_decoder_bit_T_86 == 32'h4f; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_93 = _id_ctrl_decoder_bit_T_86 == 32'h4b; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_94 = ibuf_io_inst_0_bits_inst_bits & 32'hfff0707f; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_bit_T_95 = _id_ctrl_decoder_bit_T_94 == 32'he0001053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_97 = _id_ctrl_decoder_bit_T_94 == 32'he0000053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_98 = ibuf_io_inst_0_bits_inst_bits & 32'hfff0007f; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_bit_T_99 = _id_ctrl_decoder_bit_T_98 == 32'hc0000053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_101 = _id_ctrl_decoder_bit_T_98 == 32'hc0100053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_103 = _id_ctrl_decoder_bit_T == 32'ha0002053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_105 = _id_ctrl_decoder_bit_T == 32'ha0001053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_107 = _id_ctrl_decoder_bit_T == 32'ha0000053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_109 = _id_ctrl_decoder_bit_T_94 == 32'hf0000053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_111 = _id_ctrl_decoder_bit_T_98 == 32'hd0000053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_113 = _id_ctrl_decoder_bit_T_98 == 32'hd0100053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_114 = ibuf_io_inst_0_bits_inst_bits & 32'h707f; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_bit_T_115 = _id_ctrl_decoder_bit_T_114 == 32'h2007; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_117 = _id_ctrl_decoder_bit_T_114 == 32'h2027; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_119 = _id_ctrl_decoder_bit_T_80 == 32'h18000053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_121 = _id_ctrl_decoder_bit_T_98 == 32'h58000053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_123 = _id_ctrl_decoder_bit_T_98 == 32'hc0200053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_125 = _id_ctrl_decoder_bit_T_98 == 32'hc0300053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_127 = _id_ctrl_decoder_bit_T_98 == 32'hd0200053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_129 = _id_ctrl_decoder_bit_T_98 == 32'hd0300053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_131 = _id_ctrl_decoder_bit_T_98 == 32'h40100053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_133 = _id_ctrl_decoder_bit_T_98 == 32'h42000053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_135 = _id_ctrl_decoder_bit_T == 32'h22000053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_137 = _id_ctrl_decoder_bit_T == 32'h22002053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_139 = _id_ctrl_decoder_bit_T == 32'h22001053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_141 = _id_ctrl_decoder_bit_T == 32'h2a000053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_143 = _id_ctrl_decoder_bit_T == 32'h2a001053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_145 = _id_ctrl_decoder_bit_T_80 == 32'h2000053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_147 = _id_ctrl_decoder_bit_T_80 == 32'ha000053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_149 = _id_ctrl_decoder_bit_T_80 == 32'h12000053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_151 = _id_ctrl_decoder_bit_T_86 == 32'h2000043; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_153 = _id_ctrl_decoder_bit_T_86 == 32'h2000047; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_155 = _id_ctrl_decoder_bit_T_86 == 32'h200004f; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_157 = _id_ctrl_decoder_bit_T_86 == 32'h200004b; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_159 = _id_ctrl_decoder_bit_T_94 == 32'he2001053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_161 = _id_ctrl_decoder_bit_T_98 == 32'hc2000053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_163 = _id_ctrl_decoder_bit_T_98 == 32'hc2100053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_165 = _id_ctrl_decoder_bit_T == 32'ha2002053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_167 = _id_ctrl_decoder_bit_T == 32'ha2001053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_169 = _id_ctrl_decoder_bit_T == 32'ha2000053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_171 = _id_ctrl_decoder_bit_T_98 == 32'hd2000053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_173 = _id_ctrl_decoder_bit_T_98 == 32'hd2100053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_175 = _id_ctrl_decoder_bit_T_114 == 32'h3007; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_177 = _id_ctrl_decoder_bit_T_114 == 32'h3027; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_179 = _id_ctrl_decoder_bit_T_80 == 32'h1a000053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_181 = _id_ctrl_decoder_bit_T_98 == 32'h5a000053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_183 = _id_ctrl_decoder_bit_T_94 == 32'he2000053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_185 = _id_ctrl_decoder_bit_T_98 == 32'hc2200053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_187 = _id_ctrl_decoder_bit_T_98 == 32'hc2300053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_189 = _id_ctrl_decoder_bit_T_94 == 32'hf2000053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_191 = _id_ctrl_decoder_bit_T_98 == 32'hd2200053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_193 = _id_ctrl_decoder_bit_T_98 == 32'hd2300053; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_195 = _id_ctrl_decoder_bit_T_114 == 32'h3003; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_197 = _id_ctrl_decoder_bit_T_114 == 32'h6003; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_199 = _id_ctrl_decoder_bit_T_114 == 32'h3023; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_200 = ibuf_io_inst_0_bits_inst_bits & 32'hfc00707f; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_bit_T_201 = _id_ctrl_decoder_bit_T_200 == 32'h1013; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_203 = _id_ctrl_decoder_bit_T_200 == 32'h5013; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_205 = _id_ctrl_decoder_bit_T_200 == 32'h40005013; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_207 = _id_ctrl_decoder_bit_T_114 == 32'h1b; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_209 = _id_ctrl_decoder_bit_T == 32'h101b; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_211 = _id_ctrl_decoder_bit_T == 32'h501b; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_213 = _id_ctrl_decoder_bit_T == 32'h4000501b; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_215 = _id_ctrl_decoder_bit_T == 32'h3b; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_217 = _id_ctrl_decoder_bit_T == 32'h4000003b; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_219 = _id_ctrl_decoder_bit_T == 32'h103b; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_221 = _id_ctrl_decoder_bit_T == 32'h503b; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_223 = _id_ctrl_decoder_bit_T == 32'h4000503b; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_224 = ibuf_io_inst_0_bits_inst_bits & 32'hfe007fff; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_bit_T_225 = _id_ctrl_decoder_bit_T_224 == 32'h12000073; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_226 = ibuf_io_inst_0_bits_inst_bits == 32'h10200073; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_227 = ibuf_io_inst_0_bits_inst_bits == 32'h7b200073; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_229 = _id_ctrl_decoder_bit_T_114 == 32'h100f; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_231 = _id_ctrl_decoder_bit_T_114 == 32'h1063; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_233 = _id_ctrl_decoder_bit_T_114 == 32'h63; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_235 = _id_ctrl_decoder_bit_T_114 == 32'h4063; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_237 = _id_ctrl_decoder_bit_T_114 == 32'h6063; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_239 = _id_ctrl_decoder_bit_T_114 == 32'h5063; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_241 = _id_ctrl_decoder_bit_T_114 == 32'h7063; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_242 = ibuf_io_inst_0_bits_inst_bits & 32'h7f; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_bit_T_243 = _id_ctrl_decoder_bit_T_242 == 32'h6f; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_245 = _id_ctrl_decoder_bit_T_114 == 32'h67; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_247 = _id_ctrl_decoder_bit_T_242 == 32'h17; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_249 = _id_ctrl_decoder_bit_T_114 == 32'h3; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_251 = _id_ctrl_decoder_bit_T_114 == 32'h1003; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_253 = _id_ctrl_decoder_bit_T_114 == 32'h2003; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_255 = _id_ctrl_decoder_bit_T_114 == 32'h4003; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_257 = _id_ctrl_decoder_bit_T_114 == 32'h5003; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_259 = _id_ctrl_decoder_bit_T_114 == 32'h23; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_261 = _id_ctrl_decoder_bit_T_114 == 32'h1023; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_263 = _id_ctrl_decoder_bit_T_114 == 32'h2023; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_265 = _id_ctrl_decoder_bit_T_242 == 32'h37; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_267 = _id_ctrl_decoder_bit_T_114 == 32'h13; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_269 = _id_ctrl_decoder_bit_T_114 == 32'h2013; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_271 = _id_ctrl_decoder_bit_T_114 == 32'h3013; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_273 = _id_ctrl_decoder_bit_T_114 == 32'h7013; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_275 = _id_ctrl_decoder_bit_T_114 == 32'h6013; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_277 = _id_ctrl_decoder_bit_T_114 == 32'h4013; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_279 = _id_ctrl_decoder_bit_T == 32'h33; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_281 = _id_ctrl_decoder_bit_T == 32'h40000033; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_283 = _id_ctrl_decoder_bit_T == 32'h2033; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_285 = _id_ctrl_decoder_bit_T == 32'h3033; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_287 = _id_ctrl_decoder_bit_T == 32'h7033; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_289 = _id_ctrl_decoder_bit_T == 32'h6033; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_291 = _id_ctrl_decoder_bit_T == 32'h4033; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_293 = _id_ctrl_decoder_bit_T == 32'h1033; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_295 = _id_ctrl_decoder_bit_T == 32'h5033; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_297 = _id_ctrl_decoder_bit_T == 32'h40005033; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_299 = _id_ctrl_decoder_bit_T_114 == 32'hf; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_300 = ibuf_io_inst_0_bits_inst_bits == 32'h73; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_301 = ibuf_io_inst_0_bits_inst_bits == 32'h100073; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_302 = ibuf_io_inst_0_bits_inst_bits == 32'h30200073; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_303 = ibuf_io_inst_0_bits_inst_bits == 32'h10500073; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_304 = ibuf_io_inst_0_bits_inst_bits == 32'h30500073; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_306 = _id_ctrl_decoder_bit_T_114 == 32'h1073; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_308 = _id_ctrl_decoder_bit_T_114 == 32'h2073; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_310 = _id_ctrl_decoder_bit_T_114 == 32'h3073; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_312 = _id_ctrl_decoder_bit_T_114 == 32'h5073; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_314 = _id_ctrl_decoder_bit_T_114 == 32'h6073; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_316 = _id_ctrl_decoder_bit_T_114 == 32'h7073; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_bit_T_318 = _id_ctrl_decoder_bit_T_1 | _id_ctrl_decoder_bit_T_3; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_319 = _id_ctrl_decoder_bit_T_318 | _id_ctrl_decoder_bit_T_5; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_320 = _id_ctrl_decoder_bit_T_319 | _id_ctrl_decoder_bit_T_7; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_321 = _id_ctrl_decoder_bit_T_320 | _id_ctrl_decoder_bit_T_9; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_322 = _id_ctrl_decoder_bit_T_321 | _id_ctrl_decoder_bit_T_11; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_323 = _id_ctrl_decoder_bit_T_322 | _id_ctrl_decoder_bit_T_13; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_324 = _id_ctrl_decoder_bit_T_323 | _id_ctrl_decoder_bit_T_15; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_325 = _id_ctrl_decoder_bit_T_324 | _id_ctrl_decoder_bit_T_17; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_326 = _id_ctrl_decoder_bit_T_325 | _id_ctrl_decoder_bit_T_19; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_327 = _id_ctrl_decoder_bit_T_326 | _id_ctrl_decoder_bit_T_21; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_328 = _id_ctrl_decoder_bit_T_327 | _id_ctrl_decoder_bit_T_23; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_329 = _id_ctrl_decoder_bit_T_328 | _id_ctrl_decoder_bit_T_25; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_330 = _id_ctrl_decoder_bit_T_329 | _id_ctrl_decoder_bit_T_27; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_331 = _id_ctrl_decoder_bit_T_330 | _id_ctrl_decoder_bit_T_29; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_332 = _id_ctrl_decoder_bit_T_331 | _id_ctrl_decoder_bit_T_31; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_333 = _id_ctrl_decoder_bit_T_332 | _id_ctrl_decoder_bit_T_33; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_334 = _id_ctrl_decoder_bit_T_333 | _id_ctrl_decoder_bit_T_35; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_335 = _id_ctrl_decoder_bit_T_334 | _id_ctrl_decoder_bit_T_37; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_336 = _id_ctrl_decoder_bit_T_335 | _id_ctrl_decoder_bit_T_39; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_337 = _id_ctrl_decoder_bit_T_336 | _id_ctrl_decoder_bit_T_41; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_338 = _id_ctrl_decoder_bit_T_337 | _id_ctrl_decoder_bit_T_43; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_339 = _id_ctrl_decoder_bit_T_338 | _id_ctrl_decoder_bit_T_45; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_340 = _id_ctrl_decoder_bit_T_339 | _id_ctrl_decoder_bit_T_47; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_341 = _id_ctrl_decoder_bit_T_340 | _id_ctrl_decoder_bit_T_49; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_342 = _id_ctrl_decoder_bit_T_341 | _id_ctrl_decoder_bit_T_51; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_343 = _id_ctrl_decoder_bit_T_342 | _id_ctrl_decoder_bit_T_53; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_344 = _id_ctrl_decoder_bit_T_343 | _id_ctrl_decoder_bit_T_55; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_345 = _id_ctrl_decoder_bit_T_344 | _id_ctrl_decoder_bit_T_57; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_346 = _id_ctrl_decoder_bit_T_345 | _id_ctrl_decoder_bit_T_59; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_347 = _id_ctrl_decoder_bit_T_346 | _id_ctrl_decoder_bit_T_61; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_348 = _id_ctrl_decoder_bit_T_347 | _id_ctrl_decoder_bit_T_63; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_349 = _id_ctrl_decoder_bit_T_348 | _id_ctrl_decoder_bit_T_65; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_350 = _id_ctrl_decoder_bit_T_349 | _id_ctrl_decoder_bit_T_67; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_351 = _id_ctrl_decoder_bit_T_350 | _id_ctrl_decoder_bit_T_69; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_352 = _id_ctrl_decoder_bit_T_351 | _id_ctrl_decoder_bit_T_71; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_353 = _id_ctrl_decoder_bit_T_352 | _id_ctrl_decoder_bit_T_73; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_354 = _id_ctrl_decoder_bit_T_353 | _id_ctrl_decoder_bit_T_75; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_355 = _id_ctrl_decoder_bit_T_354 | _id_ctrl_decoder_bit_T_77; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_356 = _id_ctrl_decoder_bit_T_355 | _id_ctrl_decoder_bit_T_79; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_357 = _id_ctrl_decoder_bit_T_356 | _id_ctrl_decoder_bit_T_81; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_358 = _id_ctrl_decoder_bit_T_357 | _id_ctrl_decoder_bit_T_83; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_359 = _id_ctrl_decoder_bit_T_358 | _id_ctrl_decoder_bit_T_85; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_360 = _id_ctrl_decoder_bit_T_359 | _id_ctrl_decoder_bit_T_87; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_361 = _id_ctrl_decoder_bit_T_360 | _id_ctrl_decoder_bit_T_89; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_362 = _id_ctrl_decoder_bit_T_361 | _id_ctrl_decoder_bit_T_91; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_363 = _id_ctrl_decoder_bit_T_362 | _id_ctrl_decoder_bit_T_93; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_364 = _id_ctrl_decoder_bit_T_363 | _id_ctrl_decoder_bit_T_95; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_365 = _id_ctrl_decoder_bit_T_364 | _id_ctrl_decoder_bit_T_97; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_366 = _id_ctrl_decoder_bit_T_365 | _id_ctrl_decoder_bit_T_99; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_367 = _id_ctrl_decoder_bit_T_366 | _id_ctrl_decoder_bit_T_101; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_368 = _id_ctrl_decoder_bit_T_367 | _id_ctrl_decoder_bit_T_103; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_369 = _id_ctrl_decoder_bit_T_368 | _id_ctrl_decoder_bit_T_105; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_370 = _id_ctrl_decoder_bit_T_369 | _id_ctrl_decoder_bit_T_107; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_371 = _id_ctrl_decoder_bit_T_370 | _id_ctrl_decoder_bit_T_109; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_372 = _id_ctrl_decoder_bit_T_371 | _id_ctrl_decoder_bit_T_111; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_373 = _id_ctrl_decoder_bit_T_372 | _id_ctrl_decoder_bit_T_113; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_374 = _id_ctrl_decoder_bit_T_373 | _id_ctrl_decoder_bit_T_115; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_375 = _id_ctrl_decoder_bit_T_374 | _id_ctrl_decoder_bit_T_117; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_376 = _id_ctrl_decoder_bit_T_375 | _id_ctrl_decoder_bit_T_119; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_377 = _id_ctrl_decoder_bit_T_376 | _id_ctrl_decoder_bit_T_121; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_378 = _id_ctrl_decoder_bit_T_377 | _id_ctrl_decoder_bit_T_123; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_379 = _id_ctrl_decoder_bit_T_378 | _id_ctrl_decoder_bit_T_125; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_380 = _id_ctrl_decoder_bit_T_379 | _id_ctrl_decoder_bit_T_127; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_381 = _id_ctrl_decoder_bit_T_380 | _id_ctrl_decoder_bit_T_129; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_382 = _id_ctrl_decoder_bit_T_381 | _id_ctrl_decoder_bit_T_131; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_383 = _id_ctrl_decoder_bit_T_382 | _id_ctrl_decoder_bit_T_133; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_384 = _id_ctrl_decoder_bit_T_383 | _id_ctrl_decoder_bit_T_135; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_385 = _id_ctrl_decoder_bit_T_384 | _id_ctrl_decoder_bit_T_137; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_386 = _id_ctrl_decoder_bit_T_385 | _id_ctrl_decoder_bit_T_139; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_387 = _id_ctrl_decoder_bit_T_386 | _id_ctrl_decoder_bit_T_141; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_388 = _id_ctrl_decoder_bit_T_387 | _id_ctrl_decoder_bit_T_143; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_389 = _id_ctrl_decoder_bit_T_388 | _id_ctrl_decoder_bit_T_145; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_390 = _id_ctrl_decoder_bit_T_389 | _id_ctrl_decoder_bit_T_147; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_391 = _id_ctrl_decoder_bit_T_390 | _id_ctrl_decoder_bit_T_149; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_392 = _id_ctrl_decoder_bit_T_391 | _id_ctrl_decoder_bit_T_151; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_393 = _id_ctrl_decoder_bit_T_392 | _id_ctrl_decoder_bit_T_153; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_394 = _id_ctrl_decoder_bit_T_393 | _id_ctrl_decoder_bit_T_155; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_395 = _id_ctrl_decoder_bit_T_394 | _id_ctrl_decoder_bit_T_157; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_396 = _id_ctrl_decoder_bit_T_395 | _id_ctrl_decoder_bit_T_159; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_397 = _id_ctrl_decoder_bit_T_396 | _id_ctrl_decoder_bit_T_161; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_398 = _id_ctrl_decoder_bit_T_397 | _id_ctrl_decoder_bit_T_163; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_399 = _id_ctrl_decoder_bit_T_398 | _id_ctrl_decoder_bit_T_165; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_400 = _id_ctrl_decoder_bit_T_399 | _id_ctrl_decoder_bit_T_167; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_401 = _id_ctrl_decoder_bit_T_400 | _id_ctrl_decoder_bit_T_169; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_402 = _id_ctrl_decoder_bit_T_401 | _id_ctrl_decoder_bit_T_171; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_403 = _id_ctrl_decoder_bit_T_402 | _id_ctrl_decoder_bit_T_173; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_404 = _id_ctrl_decoder_bit_T_403 | _id_ctrl_decoder_bit_T_175; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_405 = _id_ctrl_decoder_bit_T_404 | _id_ctrl_decoder_bit_T_177; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_406 = _id_ctrl_decoder_bit_T_405 | _id_ctrl_decoder_bit_T_179; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_407 = _id_ctrl_decoder_bit_T_406 | _id_ctrl_decoder_bit_T_181; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_408 = _id_ctrl_decoder_bit_T_407 | _id_ctrl_decoder_bit_T_183; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_409 = _id_ctrl_decoder_bit_T_408 | _id_ctrl_decoder_bit_T_185; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_410 = _id_ctrl_decoder_bit_T_409 | _id_ctrl_decoder_bit_T_187; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_411 = _id_ctrl_decoder_bit_T_410 | _id_ctrl_decoder_bit_T_189; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_412 = _id_ctrl_decoder_bit_T_411 | _id_ctrl_decoder_bit_T_191; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_413 = _id_ctrl_decoder_bit_T_412 | _id_ctrl_decoder_bit_T_193; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_414 = _id_ctrl_decoder_bit_T_413 | _id_ctrl_decoder_bit_T_195; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_415 = _id_ctrl_decoder_bit_T_414 | _id_ctrl_decoder_bit_T_197; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_416 = _id_ctrl_decoder_bit_T_415 | _id_ctrl_decoder_bit_T_199; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_417 = _id_ctrl_decoder_bit_T_416 | _id_ctrl_decoder_bit_T_201; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_418 = _id_ctrl_decoder_bit_T_417 | _id_ctrl_decoder_bit_T_203; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_419 = _id_ctrl_decoder_bit_T_418 | _id_ctrl_decoder_bit_T_205; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_420 = _id_ctrl_decoder_bit_T_419 | _id_ctrl_decoder_bit_T_207; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_421 = _id_ctrl_decoder_bit_T_420 | _id_ctrl_decoder_bit_T_209; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_422 = _id_ctrl_decoder_bit_T_421 | _id_ctrl_decoder_bit_T_211; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_423 = _id_ctrl_decoder_bit_T_422 | _id_ctrl_decoder_bit_T_213; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_424 = _id_ctrl_decoder_bit_T_423 | _id_ctrl_decoder_bit_T_215; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_425 = _id_ctrl_decoder_bit_T_424 | _id_ctrl_decoder_bit_T_217; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_426 = _id_ctrl_decoder_bit_T_425 | _id_ctrl_decoder_bit_T_219; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_427 = _id_ctrl_decoder_bit_T_426 | _id_ctrl_decoder_bit_T_221; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_428 = _id_ctrl_decoder_bit_T_427 | _id_ctrl_decoder_bit_T_223; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_429 = _id_ctrl_decoder_bit_T_428 | _id_ctrl_decoder_bit_T_225; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_430 = _id_ctrl_decoder_bit_T_429 | _id_ctrl_decoder_bit_T_226; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_431 = _id_ctrl_decoder_bit_T_430 | _id_ctrl_decoder_bit_T_227; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_432 = _id_ctrl_decoder_bit_T_431 | _id_ctrl_decoder_bit_T_229; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_433 = _id_ctrl_decoder_bit_T_432 | _id_ctrl_decoder_bit_T_231; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_434 = _id_ctrl_decoder_bit_T_433 | _id_ctrl_decoder_bit_T_233; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_435 = _id_ctrl_decoder_bit_T_434 | _id_ctrl_decoder_bit_T_235; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_436 = _id_ctrl_decoder_bit_T_435 | _id_ctrl_decoder_bit_T_237; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_437 = _id_ctrl_decoder_bit_T_436 | _id_ctrl_decoder_bit_T_239; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_438 = _id_ctrl_decoder_bit_T_437 | _id_ctrl_decoder_bit_T_241; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_439 = _id_ctrl_decoder_bit_T_438 | _id_ctrl_decoder_bit_T_243; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_440 = _id_ctrl_decoder_bit_T_439 | _id_ctrl_decoder_bit_T_245; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_441 = _id_ctrl_decoder_bit_T_440 | _id_ctrl_decoder_bit_T_247; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_442 = _id_ctrl_decoder_bit_T_441 | _id_ctrl_decoder_bit_T_249; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_443 = _id_ctrl_decoder_bit_T_442 | _id_ctrl_decoder_bit_T_251; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_444 = _id_ctrl_decoder_bit_T_443 | _id_ctrl_decoder_bit_T_253; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_445 = _id_ctrl_decoder_bit_T_444 | _id_ctrl_decoder_bit_T_255; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_446 = _id_ctrl_decoder_bit_T_445 | _id_ctrl_decoder_bit_T_257; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_447 = _id_ctrl_decoder_bit_T_446 | _id_ctrl_decoder_bit_T_259; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_448 = _id_ctrl_decoder_bit_T_447 | _id_ctrl_decoder_bit_T_261; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_449 = _id_ctrl_decoder_bit_T_448 | _id_ctrl_decoder_bit_T_263; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_450 = _id_ctrl_decoder_bit_T_449 | _id_ctrl_decoder_bit_T_265; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_451 = _id_ctrl_decoder_bit_T_450 | _id_ctrl_decoder_bit_T_267; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_452 = _id_ctrl_decoder_bit_T_451 | _id_ctrl_decoder_bit_T_269; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_453 = _id_ctrl_decoder_bit_T_452 | _id_ctrl_decoder_bit_T_271; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_454 = _id_ctrl_decoder_bit_T_453 | _id_ctrl_decoder_bit_T_273; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_455 = _id_ctrl_decoder_bit_T_454 | _id_ctrl_decoder_bit_T_275; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_456 = _id_ctrl_decoder_bit_T_455 | _id_ctrl_decoder_bit_T_277; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_457 = _id_ctrl_decoder_bit_T_456 | _id_ctrl_decoder_bit_T_279; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_458 = _id_ctrl_decoder_bit_T_457 | _id_ctrl_decoder_bit_T_281; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_459 = _id_ctrl_decoder_bit_T_458 | _id_ctrl_decoder_bit_T_283; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_460 = _id_ctrl_decoder_bit_T_459 | _id_ctrl_decoder_bit_T_285; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_461 = _id_ctrl_decoder_bit_T_460 | _id_ctrl_decoder_bit_T_287; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_462 = _id_ctrl_decoder_bit_T_461 | _id_ctrl_decoder_bit_T_289; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_463 = _id_ctrl_decoder_bit_T_462 | _id_ctrl_decoder_bit_T_291; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_464 = _id_ctrl_decoder_bit_T_463 | _id_ctrl_decoder_bit_T_293; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_465 = _id_ctrl_decoder_bit_T_464 | _id_ctrl_decoder_bit_T_295; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_466 = _id_ctrl_decoder_bit_T_465 | _id_ctrl_decoder_bit_T_297; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_467 = _id_ctrl_decoder_bit_T_466 | _id_ctrl_decoder_bit_T_299; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_468 = _id_ctrl_decoder_bit_T_467 | _id_ctrl_decoder_bit_T_300; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_469 = _id_ctrl_decoder_bit_T_468 | _id_ctrl_decoder_bit_T_301; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_470 = _id_ctrl_decoder_bit_T_469 | _id_ctrl_decoder_bit_T_302; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_471 = _id_ctrl_decoder_bit_T_470 | _id_ctrl_decoder_bit_T_303; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_472 = _id_ctrl_decoder_bit_T_471 | _id_ctrl_decoder_bit_T_304; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_473 = _id_ctrl_decoder_bit_T_472 | _id_ctrl_decoder_bit_T_306; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_474 = _id_ctrl_decoder_bit_T_473 | _id_ctrl_decoder_bit_T_308; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_475 = _id_ctrl_decoder_bit_T_474 | _id_ctrl_decoder_bit_T_310; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_476 = _id_ctrl_decoder_bit_T_475 | _id_ctrl_decoder_bit_T_312; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_477 = _id_ctrl_decoder_bit_T_476 | _id_ctrl_decoder_bit_T_314; // @[Decode.scala 15:30]
  assign id_ctrl_decoder_0 = _id_ctrl_decoder_bit_T_477 | _id_ctrl_decoder_bit_T_316; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_T = ibuf_io_inst_0_bits_inst_bits & 32'h5c; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_1 = _id_ctrl_decoder_T == 32'h4; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_2 = ibuf_io_inst_0_bits_inst_bits & 32'h60; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_3 = _id_ctrl_decoder_T_2 == 32'h40; // @[Decode.scala 14:121]
  assign id_ctrl_decoder_1 = _id_ctrl_decoder_T_1 | _id_ctrl_decoder_T_3; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_T_5 = ibuf_io_inst_0_bits_inst_bits & 32'h74; // @[Decode.scala 14:65]
  assign id_ctrl_decoder_3 = _id_ctrl_decoder_T_5 == 32'h60; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_7 = ibuf_io_inst_0_bits_inst_bits & 32'h68; // @[Decode.scala 14:65]
  assign id_ctrl_decoder_4 = _id_ctrl_decoder_T_7 == 32'h68; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_9 = ibuf_io_inst_0_bits_inst_bits & 32'h203c; // @[Decode.scala 14:65]
  assign id_ctrl_decoder_5 = _id_ctrl_decoder_T_9 == 32'h24; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_11 = ibuf_io_inst_0_bits_inst_bits & 32'h64; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_12 = _id_ctrl_decoder_T_11 == 32'h20; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_13 = ibuf_io_inst_0_bits_inst_bits & 32'h34; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_14 = _id_ctrl_decoder_T_13 == 32'h20; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_15 = ibuf_io_inst_0_bits_inst_bits & 32'h2048; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_16 = _id_ctrl_decoder_T_15 == 32'h2008; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_17 = ibuf_io_inst_0_bits_inst_bits & 32'h42003024; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_18 = _id_ctrl_decoder_T_17 == 32'h2000020; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_20 = _id_ctrl_decoder_T_12 | _id_ctrl_decoder_T_14; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_T_21 = _id_ctrl_decoder_T_20 | _id_ctrl_decoder_T_16; // @[Decode.scala 15:30]
  assign id_ctrl_decoder_6 = _id_ctrl_decoder_T_21 | _id_ctrl_decoder_T_18; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_T_22 = ibuf_io_inst_0_bits_inst_bits & 32'h44; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_23 = _id_ctrl_decoder_T_22 == 32'h0; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_24 = ibuf_io_inst_0_bits_inst_bits & 32'h4024; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_25 = _id_ctrl_decoder_T_24 == 32'h20; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_26 = ibuf_io_inst_0_bits_inst_bits & 32'h38; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_27 = _id_ctrl_decoder_T_26 == 32'h20; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_28 = ibuf_io_inst_0_bits_inst_bits & 32'h2050; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_29 = _id_ctrl_decoder_T_28 == 32'h2000; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_30 = ibuf_io_inst_0_bits_inst_bits & 32'h90000034; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_31 = _id_ctrl_decoder_T_30 == 32'h90000010; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_33 = _id_ctrl_decoder_T_23 | _id_ctrl_decoder_T_25; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_T_34 = _id_ctrl_decoder_T_33 | _id_ctrl_decoder_T_27; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_T_35 = _id_ctrl_decoder_T_34 | _id_ctrl_decoder_T_29; // @[Decode.scala 15:30]
  assign id_ctrl_decoder_7 = _id_ctrl_decoder_T_35 | _id_ctrl_decoder_T_31; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_T_36 = ibuf_io_inst_0_bits_inst_bits & 32'h58; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_37 = _id_ctrl_decoder_T_36 == 32'h0; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_38 = ibuf_io_inst_0_bits_inst_bits & 32'h20; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_39 = _id_ctrl_decoder_T_38 == 32'h0; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_40 = ibuf_io_inst_0_bits_inst_bits & 32'hc; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_41 = _id_ctrl_decoder_T_40 == 32'h4; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_42 = ibuf_io_inst_0_bits_inst_bits & 32'h48; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_43 = _id_ctrl_decoder_T_42 == 32'h48; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_44 = ibuf_io_inst_0_bits_inst_bits & 32'h4050; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_45 = _id_ctrl_decoder_T_44 == 32'h4050; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_47 = _id_ctrl_decoder_T_37 | _id_ctrl_decoder_T_39; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_T_48 = _id_ctrl_decoder_T_47 | _id_ctrl_decoder_T_41; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_T_49 = _id_ctrl_decoder_T_48 | _id_ctrl_decoder_T_43; // @[Decode.scala 15:30]
  assign id_ctrl_decoder_lo = _id_ctrl_decoder_T_49 | _id_ctrl_decoder_T_45; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_T_51 = _id_ctrl_decoder_T_42 == 32'h0; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_52 = ibuf_io_inst_0_bits_inst_bits & 32'h18; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_53 = _id_ctrl_decoder_T_52 == 32'h0; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_54 = ibuf_io_inst_0_bits_inst_bits & 32'h4008; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_55 = _id_ctrl_decoder_T_54 == 32'h4000; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_57 = _id_ctrl_decoder_T_51 | _id_ctrl_decoder_T_23; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_T_58 = _id_ctrl_decoder_T_57 | _id_ctrl_decoder_T_53; // @[Decode.scala 15:30]
  assign id_ctrl_decoder_hi = _id_ctrl_decoder_T_58 | _id_ctrl_decoder_T_55; // @[Decode.scala 15:30]
  assign id_ctrl_decoder_9 = {id_ctrl_decoder_hi,id_ctrl_decoder_lo}; // @[Cat.scala 30:58]
  assign _id_ctrl_decoder_T_59 = ibuf_io_inst_0_bits_inst_bits & 32'h4004; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_60 = _id_ctrl_decoder_T_59 == 32'h0; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_61 = ibuf_io_inst_0_bits_inst_bits & 32'h50; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_62 = _id_ctrl_decoder_T_61 == 32'h0; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_63 = ibuf_io_inst_0_bits_inst_bits & 32'h24; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_64 = _id_ctrl_decoder_T_63 == 32'h0; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_66 = _id_ctrl_decoder_T_60 | _id_ctrl_decoder_T_62; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_T_67 = _id_ctrl_decoder_T_66 | _id_ctrl_decoder_T_23; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_T_68 = _id_ctrl_decoder_T_67 | _id_ctrl_decoder_T_64; // @[Decode.scala 15:30]
  assign id_ctrl_decoder_lo_1 = _id_ctrl_decoder_T_68 | _id_ctrl_decoder_T_53; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_T_70 = _id_ctrl_decoder_T_13 == 32'h14; // @[Decode.scala 14:121]
  assign id_ctrl_decoder_hi_1 = _id_ctrl_decoder_T_70 | _id_ctrl_decoder_T_43; // @[Decode.scala 15:30]
  assign id_ctrl_decoder_10 = {id_ctrl_decoder_hi_1,id_ctrl_decoder_lo_1}; // @[Cat.scala 30:58]
  assign _id_ctrl_decoder_T_73 = _id_ctrl_decoder_T_52 == 32'h8; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_75 = _id_ctrl_decoder_T_22 == 32'h40; // @[Decode.scala 14:121]
  assign id_ctrl_decoder_lo_2 = _id_ctrl_decoder_T_73 | _id_ctrl_decoder_T_75; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_T_77 = ibuf_io_inst_0_bits_inst_bits & 32'h14; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_78 = _id_ctrl_decoder_T_77 == 32'h14; // @[Decode.scala 14:121]
  assign id_ctrl_decoder_hi_lo = _id_ctrl_decoder_T_73 | _id_ctrl_decoder_T_78; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_T_80 = ibuf_io_inst_0_bits_inst_bits & 32'h30; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_81 = _id_ctrl_decoder_T_80 == 32'h0; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_82 = ibuf_io_inst_0_bits_inst_bits & 32'h201c; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_83 = _id_ctrl_decoder_T_82 == 32'h4; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_85 = _id_ctrl_decoder_T_77 == 32'h10; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_87 = _id_ctrl_decoder_T_81 | _id_ctrl_decoder_T_83; // @[Decode.scala 15:30]
  assign id_ctrl_decoder_hi_hi = _id_ctrl_decoder_T_87 | _id_ctrl_decoder_T_85; // @[Decode.scala 15:30]
  assign id_ctrl_decoder_11 = {id_ctrl_decoder_hi_hi,id_ctrl_decoder_hi_lo,id_ctrl_decoder_lo_2}; // @[Cat.scala 30:58]
  assign _id_ctrl_decoder_T_88 = ibuf_io_inst_0_bits_inst_bits & 32'h10; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_89 = _id_ctrl_decoder_T_88 == 32'h0; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_90 = ibuf_io_inst_0_bits_inst_bits & 32'h8; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_91 = _id_ctrl_decoder_T_90 == 32'h0; // @[Decode.scala 14:121]
  assign id_ctrl_decoder_12 = _id_ctrl_decoder_T_89 | _id_ctrl_decoder_T_91; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_T_93 = ibuf_io_inst_0_bits_inst_bits & 32'h3054; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_94 = _id_ctrl_decoder_T_93 == 32'h1010; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_95 = ibuf_io_inst_0_bits_inst_bits & 32'h1058; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_96 = _id_ctrl_decoder_T_95 == 32'h1040; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_97 = ibuf_io_inst_0_bits_inst_bits & 32'h7044; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_98 = _id_ctrl_decoder_T_97 == 32'h7000; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_99 = ibuf_io_inst_0_bits_inst_bits & 32'h2001074; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_100 = _id_ctrl_decoder_T_99 == 32'h2001030; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_102 = _id_ctrl_decoder_T_94 | _id_ctrl_decoder_T_96; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_T_103 = _id_ctrl_decoder_T_102 | _id_ctrl_decoder_T_98; // @[Decode.scala 15:30]
  assign id_ctrl_decoder_lo_lo = _id_ctrl_decoder_T_103 | _id_ctrl_decoder_T_100; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_T_104 = ibuf_io_inst_0_bits_inst_bits & 32'h4054; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_105 = _id_ctrl_decoder_T_104 == 32'h40; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_106 = ibuf_io_inst_0_bits_inst_bits & 32'h2058; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_107 = _id_ctrl_decoder_T_106 == 32'h2040; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_109 = _id_ctrl_decoder_T_93 == 32'h3010; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_110 = ibuf_io_inst_0_bits_inst_bits & 32'h6054; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_111 = _id_ctrl_decoder_T_110 == 32'h6010; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_112 = ibuf_io_inst_0_bits_inst_bits & 32'h2002074; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_113 = _id_ctrl_decoder_T_112 == 32'h2002030; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_114 = ibuf_io_inst_0_bits_inst_bits & 32'h40003034; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_115 = _id_ctrl_decoder_T_114 == 32'h40000030; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_116 = ibuf_io_inst_0_bits_inst_bits & 32'h40001054; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_117 = _id_ctrl_decoder_T_116 == 32'h40001010; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_119 = _id_ctrl_decoder_T_105 | _id_ctrl_decoder_T_107; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_T_120 = _id_ctrl_decoder_T_119 | _id_ctrl_decoder_T_109; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_T_121 = _id_ctrl_decoder_T_120 | _id_ctrl_decoder_T_111; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_T_122 = _id_ctrl_decoder_T_121 | _id_ctrl_decoder_T_113; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_T_123 = _id_ctrl_decoder_T_122 | _id_ctrl_decoder_T_115; // @[Decode.scala 15:30]
  assign id_ctrl_decoder_lo_hi = _id_ctrl_decoder_T_123 | _id_ctrl_decoder_T_117; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_T_124 = ibuf_io_inst_0_bits_inst_bits & 32'h2002054; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_125 = _id_ctrl_decoder_T_124 == 32'h2010; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_126 = ibuf_io_inst_0_bits_inst_bits & 32'h2034; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_127 = _id_ctrl_decoder_T_126 == 32'h2010; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_128 = ibuf_io_inst_0_bits_inst_bits & 32'h40004054; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_129 = _id_ctrl_decoder_T_128 == 32'h4010; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_130 = ibuf_io_inst_0_bits_inst_bits & 32'h5054; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_131 = _id_ctrl_decoder_T_130 == 32'h4010; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_132 = ibuf_io_inst_0_bits_inst_bits & 32'h4058; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_133 = _id_ctrl_decoder_T_132 == 32'h4040; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_135 = _id_ctrl_decoder_T_125 | _id_ctrl_decoder_T_127; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_T_136 = _id_ctrl_decoder_T_135 | _id_ctrl_decoder_T_129; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_T_137 = _id_ctrl_decoder_T_136 | _id_ctrl_decoder_T_131; // @[Decode.scala 15:30]
  assign id_ctrl_decoder_hi_lo_1 = _id_ctrl_decoder_T_137 | _id_ctrl_decoder_T_133; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_T_138 = ibuf_io_inst_0_bits_inst_bits & 32'h2006054; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_139 = _id_ctrl_decoder_T_138 == 32'h2010; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_140 = ibuf_io_inst_0_bits_inst_bits & 32'h6034; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_141 = _id_ctrl_decoder_T_140 == 32'h2010; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_142 = ibuf_io_inst_0_bits_inst_bits & 32'h40003054; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_143 = _id_ctrl_decoder_T_142 == 32'h40001010; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_145 = _id_ctrl_decoder_T_139 | _id_ctrl_decoder_T_141; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_T_146 = _id_ctrl_decoder_T_145 | _id_ctrl_decoder_T_133; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_T_147 = _id_ctrl_decoder_T_146 | _id_ctrl_decoder_T_115; // @[Decode.scala 15:30]
  assign id_ctrl_decoder_hi_hi_1 = _id_ctrl_decoder_T_147 | _id_ctrl_decoder_T_143; // @[Decode.scala 15:30]
  assign id_ctrl_decoder_13 = {id_ctrl_decoder_hi_hi_1,id_ctrl_decoder_hi_lo_1,id_ctrl_decoder_lo_hi,id_ctrl_decoder_lo_lo}; // @[Cat.scala 30:58]
  assign _id_ctrl_decoder_bit_T_479 = _id_ctrl_decoder_bit_T_27 | _id_ctrl_decoder_bit_T_29; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_480 = _id_ctrl_decoder_bit_T_479 | _id_ctrl_decoder_bit_T_31; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_481 = _id_ctrl_decoder_bit_T_480 | _id_ctrl_decoder_bit_T_33; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_482 = _id_ctrl_decoder_bit_T_481 | _id_ctrl_decoder_bit_T_35; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_483 = _id_ctrl_decoder_bit_T_482 | _id_ctrl_decoder_bit_T_37; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_484 = _id_ctrl_decoder_bit_T_483 | _id_ctrl_decoder_bit_T_39; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_485 = _id_ctrl_decoder_bit_T_484 | _id_ctrl_decoder_bit_T_41; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_486 = _id_ctrl_decoder_bit_T_485 | _id_ctrl_decoder_bit_T_43; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_487 = _id_ctrl_decoder_bit_T_486 | _id_ctrl_decoder_bit_T_45; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_488 = _id_ctrl_decoder_bit_T_487 | _id_ctrl_decoder_bit_T_47; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_489 = _id_ctrl_decoder_bit_T_488 | _id_ctrl_decoder_bit_T_49; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_490 = _id_ctrl_decoder_bit_T_489 | _id_ctrl_decoder_bit_T_51; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_491 = _id_ctrl_decoder_bit_T_490 | _id_ctrl_decoder_bit_T_53; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_492 = _id_ctrl_decoder_bit_T_491 | _id_ctrl_decoder_bit_T_55; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_493 = _id_ctrl_decoder_bit_T_492 | _id_ctrl_decoder_bit_T_57; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_494 = _id_ctrl_decoder_bit_T_493 | _id_ctrl_decoder_bit_T_59; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_495 = _id_ctrl_decoder_bit_T_494 | _id_ctrl_decoder_bit_T_61; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_496 = _id_ctrl_decoder_bit_T_495 | _id_ctrl_decoder_bit_T_63; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_497 = _id_ctrl_decoder_bit_T_496 | _id_ctrl_decoder_bit_T_65; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_498 = _id_ctrl_decoder_bit_T_497 | _id_ctrl_decoder_bit_T_67; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_499 = _id_ctrl_decoder_bit_T_498 | _id_ctrl_decoder_bit_T_69; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_500 = _id_ctrl_decoder_bit_T_499 | _id_ctrl_decoder_bit_T_115; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_501 = _id_ctrl_decoder_bit_T_500 | _id_ctrl_decoder_bit_T_117; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_502 = _id_ctrl_decoder_bit_T_501 | _id_ctrl_decoder_bit_T_175; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_503 = _id_ctrl_decoder_bit_T_502 | _id_ctrl_decoder_bit_T_177; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_504 = _id_ctrl_decoder_bit_T_503 | _id_ctrl_decoder_bit_T_195; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_505 = _id_ctrl_decoder_bit_T_504 | _id_ctrl_decoder_bit_T_197; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_506 = _id_ctrl_decoder_bit_T_505 | _id_ctrl_decoder_bit_T_199; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_507 = _id_ctrl_decoder_bit_T_506 | _id_ctrl_decoder_bit_T_225; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_508 = _id_ctrl_decoder_bit_T_507 | _id_ctrl_decoder_bit_T_249; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_509 = _id_ctrl_decoder_bit_T_508 | _id_ctrl_decoder_bit_T_251; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_510 = _id_ctrl_decoder_bit_T_509 | _id_ctrl_decoder_bit_T_253; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_511 = _id_ctrl_decoder_bit_T_510 | _id_ctrl_decoder_bit_T_255; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_512 = _id_ctrl_decoder_bit_T_511 | _id_ctrl_decoder_bit_T_257; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_513 = _id_ctrl_decoder_bit_T_512 | _id_ctrl_decoder_bit_T_259; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_bit_T_514 = _id_ctrl_decoder_bit_T_513 | _id_ctrl_decoder_bit_T_261; // @[Decode.scala 15:30]
  assign id_ctrl_decoder_14 = _id_ctrl_decoder_bit_T_514 | _id_ctrl_decoder_bit_T_263; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_T_149 = _id_ctrl_decoder_T_7 == 32'h20; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_150 = ibuf_io_inst_0_bits_inst_bits & 32'h18000020; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_151 = _id_ctrl_decoder_T_150 == 32'h18000020; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_152 = ibuf_io_inst_0_bits_inst_bits & 32'h20000020; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_153 = _id_ctrl_decoder_T_152 == 32'h20000020; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_155 = _id_ctrl_decoder_T_149 | _id_ctrl_decoder_T_151; // @[Decode.scala 15:30]
  assign id_ctrl_decoder_lo_lo_1 = _id_ctrl_decoder_T_155 | _id_ctrl_decoder_T_153; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_T_156 = ibuf_io_inst_0_bits_inst_bits & 32'h10000008; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_157 = _id_ctrl_decoder_T_156 == 32'h10000008; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_158 = ibuf_io_inst_0_bits_inst_bits & 32'h40000008; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_159 = _id_ctrl_decoder_T_158 == 32'h40000008; // @[Decode.scala 14:121]
  assign id_ctrl_decoder_lo_hi_1 = _id_ctrl_decoder_T_157 | _id_ctrl_decoder_T_159; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_T_161 = ibuf_io_inst_0_bits_inst_bits & 32'h40; // @[Decode.scala 14:65]
  assign id_ctrl_decoder_hi_hi_hi = _id_ctrl_decoder_T_161 == 32'h40; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_163 = ibuf_io_inst_0_bits_inst_bits & 32'h8000008; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_164 = _id_ctrl_decoder_T_163 == 32'h8000008; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_165 = ibuf_io_inst_0_bits_inst_bits & 32'h80000008; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_166 = _id_ctrl_decoder_T_165 == 32'h80000008; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_168 = id_ctrl_decoder_hi_hi_hi | _id_ctrl_decoder_T_164; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_T_169 = _id_ctrl_decoder_T_168 | _id_ctrl_decoder_T_157; // @[Decode.scala 15:30]
  assign id_ctrl_decoder_hi_lo_2 = _id_ctrl_decoder_T_169 | _id_ctrl_decoder_T_166; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_T_170 = ibuf_io_inst_0_bits_inst_bits & 32'h18000008; // @[Decode.scala 14:65]
  assign id_ctrl_decoder_hi_hi_lo = _id_ctrl_decoder_T_170 == 32'h8; // @[Decode.scala 14:121]
  assign id_ctrl_decoder_15 = {id_ctrl_decoder_hi_hi_hi,id_ctrl_decoder_hi_hi_lo,id_ctrl_decoder_hi_lo_2,id_ctrl_decoder_lo_hi_1,id_ctrl_decoder_lo_lo_1}; // @[Cat.scala 30:58]
  assign _id_ctrl_decoder_T_172 = ibuf_io_inst_0_bits_inst_bits & 32'h80000060; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_173 = _id_ctrl_decoder_T_172 == 32'h40; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_174 = ibuf_io_inst_0_bits_inst_bits & 32'h10000060; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_176 = ibuf_io_inst_0_bits_inst_bits & 32'h70; // @[Decode.scala 14:65]
  assign id_ctrl_decoder_18 = _id_ctrl_decoder_T_176 == 32'h40; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_189 = ibuf_io_inst_0_bits_inst_bits & 32'h3c; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_190 = _id_ctrl_decoder_T_189 == 32'h4; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_192 = _id_ctrl_decoder_T_174 == 32'h10000040; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_194 = _id_ctrl_decoder_T_190 | _id_ctrl_decoder_T_173; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_T_195 = _id_ctrl_decoder_T_194 | id_ctrl_decoder_18; // @[Decode.scala 15:30]
  assign id_ctrl_decoder_19 = _id_ctrl_decoder_T_195 | _id_ctrl_decoder_T_192; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_T_196 = ibuf_io_inst_0_bits_inst_bits & 32'h2000074; // @[Decode.scala 14:65]
  assign id_ctrl_decoder_21 = _id_ctrl_decoder_T_196 == 32'h2000030; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_199 = _id_ctrl_decoder_T_11 == 32'h0; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_201 = _id_ctrl_decoder_T_61 == 32'h10; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_202 = ibuf_io_inst_0_bits_inst_bits & 32'h2024; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_203 = _id_ctrl_decoder_T_202 == 32'h24; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_204 = ibuf_io_inst_0_bits_inst_bits & 32'h28; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_205 = _id_ctrl_decoder_T_204 == 32'h28; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_206 = ibuf_io_inst_0_bits_inst_bits & 32'h1030; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_207 = _id_ctrl_decoder_T_206 == 32'h1030; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_208 = ibuf_io_inst_0_bits_inst_bits & 32'h2030; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_209 = _id_ctrl_decoder_T_208 == 32'h2030; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_210 = ibuf_io_inst_0_bits_inst_bits & 32'h90000010; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_211 = _id_ctrl_decoder_T_210 == 32'h80000010; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_213 = _id_ctrl_decoder_T_199 | _id_ctrl_decoder_T_201; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_T_214 = _id_ctrl_decoder_T_213 | _id_ctrl_decoder_T_203; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_T_215 = _id_ctrl_decoder_T_214 | _id_ctrl_decoder_T_205; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_T_216 = _id_ctrl_decoder_T_215 | _id_ctrl_decoder_T_207; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_T_217 = _id_ctrl_decoder_T_216 | _id_ctrl_decoder_T_209; // @[Decode.scala 15:30]
  assign id_ctrl_decoder_22 = _id_ctrl_decoder_T_217 | _id_ctrl_decoder_T_211; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_T_218 = ibuf_io_inst_0_bits_inst_bits & 32'h1070; // @[Decode.scala 14:65]
  assign id_ctrl_decoder_lo_5 = _id_ctrl_decoder_T_218 == 32'h1070; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_220 = ibuf_io_inst_0_bits_inst_bits & 32'h2070; // @[Decode.scala 14:65]
  assign id_ctrl_decoder_hi_lo_3 = _id_ctrl_decoder_T_220 == 32'h2070; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_222 = ibuf_io_inst_0_bits_inst_bits & 32'h10000070; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_223 = _id_ctrl_decoder_T_222 == 32'h70; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_224 = ibuf_io_inst_0_bits_inst_bits & 32'h12000034; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_225 = _id_ctrl_decoder_T_224 == 32'h10000030; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_226 = ibuf_io_inst_0_bits_inst_bits & 32'he0000050; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_227 = _id_ctrl_decoder_T_226 == 32'h60000050; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_229 = _id_ctrl_decoder_T_223 | id_ctrl_decoder_lo_5; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_T_230 = _id_ctrl_decoder_T_229 | id_ctrl_decoder_hi_lo_3; // @[Decode.scala 15:30]
  assign _id_ctrl_decoder_T_231 = _id_ctrl_decoder_T_230 | _id_ctrl_decoder_T_225; // @[Decode.scala 15:30]
  assign id_ctrl_decoder_hi_hi_3 = _id_ctrl_decoder_T_231 | _id_ctrl_decoder_T_227; // @[Decode.scala 15:30]
  assign id_ctrl_decoder_23 = {id_ctrl_decoder_hi_hi_3,id_ctrl_decoder_hi_lo_3,id_ctrl_decoder_lo_5}; // @[Cat.scala 30:58]
  assign _id_ctrl_decoder_T_232 = ibuf_io_inst_0_bits_inst_bits & 32'h3058; // @[Decode.scala 14:65]
  assign id_ctrl_decoder_24 = _id_ctrl_decoder_T_232 == 32'h1008; // @[Decode.scala 14:121]
  assign id_ctrl_decoder_25 = _id_ctrl_decoder_T_106 == 32'h8; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_236 = ibuf_io_inst_0_bits_inst_bits & 32'h6048; // @[Decode.scala 14:65]
  assign id_ctrl_decoder_26 = _id_ctrl_decoder_T_236 == 32'h2008; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_238 = ibuf_io_inst_0_bits_inst_bits & 32'h105c; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_239 = _id_ctrl_decoder_T_238 == 32'h1004; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_240 = ibuf_io_inst_0_bits_inst_bits & 32'h2000060; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_241 = _id_ctrl_decoder_T_240 == 32'h2000040; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_242 = ibuf_io_inst_0_bits_inst_bits & 32'hd0000070; // @[Decode.scala 14:65]
  assign _id_ctrl_decoder_T_243 = _id_ctrl_decoder_T_242 == 32'h40000050; // @[Decode.scala 14:121]
  assign _id_ctrl_decoder_T_245 = _id_ctrl_decoder_T_239 | _id_ctrl_decoder_T_241; // @[Decode.scala 15:30]
  assign id_ctrl_decoder_27 = _id_ctrl_decoder_T_245 | _id_ctrl_decoder_T_243; // @[Decode.scala 15:30]
  assign id_raddr3 = ibuf_io_inst_0_bits_inst_rs3; // @[RocketCore.scala 267:72]
  assign id_raddr2 = ibuf_io_inst_0_bits_inst_rs2; // @[RocketCore.scala 267:72]
  assign id_raddr1 = ibuf_io_inst_0_bits_inst_rs1; // @[RocketCore.scala 267:72]
  assign id_waddr = ibuf_io_inst_0_bits_inst_rd; // @[RocketCore.scala 267:72]
  assign _id_rs_T_4 = rf_id_rs_MPORT_data; // @[RocketCore.scala 1022:25]
  assign _id_rs_T_9 = rf_id_rs_MPORT_1_data; // @[RocketCore.scala 1022:25]
  assign _id_csr_en_T = id_ctrl_decoder_23 == 3'h6; // @[package.scala 15:47]
  assign _id_csr_en_T_1 = id_ctrl_decoder_23 == 3'h7; // @[package.scala 15:47]
  assign _id_csr_en_T_2 = id_ctrl_decoder_23 == 3'h5; // @[package.scala 15:47]
  assign _id_csr_en_T_3 = _id_csr_en_T | _id_csr_en_T_1; // @[package.scala 72:59]
  assign id_csr_en = _id_csr_en_T_3 | _id_csr_en_T_2; // @[package.scala 72:59]
  assign id_system_insn = id_ctrl_decoder_23 == 3'h4; // @[RocketCore.scala 284:36]
  assign _id_csr_ren_T_3 = ibuf_io_inst_0_bits_inst_rs1 == 5'h0; // @[RocketCore.scala 285:81]
  assign id_csr_ren = _id_csr_en_T_3 & _id_csr_ren_T_3; // @[RocketCore.scala 285:54]
  assign _id_sfence_T = id_ctrl_decoder_15 == 5'h14; // @[RocketCore.scala 287:50]
  assign id_sfence = id_ctrl_decoder_14 & _id_sfence_T; // @[RocketCore.scala 287:31]
  assign _id_csr_flush_T = id_sfence | id_system_insn; // @[RocketCore.scala 288:32]
  assign _id_csr_flush_T_2 = id_csr_en & ~id_csr_ren; // @[RocketCore.scala 288:64]
  assign _id_csr_flush_T_3 = _id_csr_flush_T_2 & csr_io_decode_0_write_flush; // @[RocketCore.scala 288:79]
  assign id_csr_flush = _id_csr_flush_T | _id_csr_flush_T_3; // @[RocketCore.scala 288:50]
  assign _id_illegal_insn_T_4 = id_ctrl_decoder_21 & ~csr_io_status_isa[12]; // @[RocketCore.scala 297:34]
  assign _id_illegal_insn_T_5 = ~id_ctrl_decoder_0 | _id_illegal_insn_T_4; // @[RocketCore.scala 296:40]
  assign _id_illegal_insn_T_8 = id_ctrl_decoder_26 & ~csr_io_status_isa[0]; // @[RocketCore.scala 298:17]
  assign _id_illegal_insn_T_9 = _id_illegal_insn_T_5 | _id_illegal_insn_T_8; // @[RocketCore.scala 297:65]
  assign _id_illegal_insn_T_10 = csr_io_decode_0_fp_illegal | io_fpu_illegal_rm; // @[RocketCore.scala 299:48]
  assign _id_illegal_insn_T_11 = id_ctrl_decoder_1 & _id_illegal_insn_T_10; // @[RocketCore.scala 299:16]
  assign _id_illegal_insn_T_12 = _id_illegal_insn_T_9 | _id_illegal_insn_T_11; // @[RocketCore.scala 298:48]
  assign _id_illegal_insn_T_15 = id_ctrl_decoder_27 & ~csr_io_status_isa[3]; // @[RocketCore.scala 300:16]
  assign _id_illegal_insn_T_16 = _id_illegal_insn_T_12 | _id_illegal_insn_T_15; // @[RocketCore.scala 299:70]
  assign _id_illegal_insn_T_19 = ibuf_io_inst_0_bits_rvc & ~csr_io_status_isa[2]; // @[RocketCore.scala 301:30]
  assign _id_illegal_insn_T_20 = _id_illegal_insn_T_16 | _id_illegal_insn_T_19; // @[RocketCore.scala 300:47]
  assign _id_illegal_insn_T_40 = ~id_csr_ren & csr_io_decode_0_write_illegal; // @[RocketCore.scala 307:64]
  assign _id_illegal_insn_T_41 = csr_io_decode_0_read_illegal | _id_illegal_insn_T_40; // @[RocketCore.scala 307:49]
  assign _id_illegal_insn_T_42 = id_csr_en & _id_illegal_insn_T_41; // @[RocketCore.scala 307:15]
  assign _id_illegal_insn_T_43 = _id_illegal_insn_T_20 | _id_illegal_insn_T_42; // @[RocketCore.scala 306:81]
  assign _id_illegal_insn_T_46 = _id_csr_flush_T & csr_io_decode_0_system_illegal; // @[RocketCore.scala 308:65]
  assign _id_illegal_insn_T_47 = ~ibuf_io_inst_0_bits_rvc & _id_illegal_insn_T_46; // @[RocketCore.scala 308:31]
  assign id_illegal_insn = _id_illegal_insn_T_43 | _id_illegal_insn_T_47; // @[RocketCore.scala 307:99]
  assign id_amo_aq = ibuf_io_inst_0_bits_inst_bits[26]; // @[RocketCore.scala 310:29]
  assign id_amo_rl = ibuf_io_inst_0_bits_inst_bits[25]; // @[RocketCore.scala 311:29]
  assign id_fence_succ = ibuf_io_inst_0_bits_inst_bits[23:20]; // @[RocketCore.scala 313:33]
  assign _id_fence_next_T = id_ctrl_decoder_26 & id_amo_aq; // @[RocketCore.scala 314:52]
  assign id_fence_next = id_ctrl_decoder_25 | _id_fence_next_T; // @[RocketCore.scala 314:37]
  assign id_mem_busy = ~io_dmem_ordered | io_dmem_req_valid; // @[RocketCore.scala 315:38]
  assign _GEN_0 = id_mem_busy ? id_reg_fence : 1'h0; // @[RocketCore.scala 316:23]
  assign _id_do_fence_x8_T_1 = id_ctrl_decoder_26 & id_amo_rl; // @[RocketCore.scala 321:33]
  assign _id_do_fence_x8_T_2 = _id_do_fence_x8_T_1 | id_ctrl_decoder_24; // @[RocketCore.scala 321:46]
  assign _id_do_fence_x8_T_4 = id_reg_fence & id_ctrl_decoder_14; // @[RocketCore.scala 321:81]
  assign _id_do_fence_x8_T_5 = _id_do_fence_x8_T_2 | _id_do_fence_x8_T_4; // @[RocketCore.scala 321:65]
  assign id_do_fence_x8 = id_mem_busy & _id_do_fence_x8_T_5; // @[RocketCore.scala 321:17]
  assign _T_1 = csr_io_interrupt | bpu_io_debug_if; // @[RocketCore.scala 975:26]
  assign _T_2 = _T_1 | bpu_io_xcpt_if; // @[RocketCore.scala 975:26]
  assign _T_3 = _T_2 | ibuf_io_inst_0_bits_xcpt0_pf_inst; // @[RocketCore.scala 975:26]
  assign _T_4 = _T_3 | ibuf_io_inst_0_bits_xcpt0_ae_inst; // @[RocketCore.scala 975:26]
  assign _T_5 = _T_4 | ibuf_io_inst_0_bits_xcpt1_pf_inst; // @[RocketCore.scala 975:26]
  assign _T_6 = _T_5 | ibuf_io_inst_0_bits_xcpt1_ae_inst; // @[RocketCore.scala 975:26]
  assign id_xcpt = _T_6 | id_illegal_insn; // @[RocketCore.scala 975:26]
  assign _T_7 = ibuf_io_inst_0_bits_xcpt1_ae_inst ? 2'h1 : 2'h2; // @[Mux.scala 47:69]
  assign _T_8 = ibuf_io_inst_0_bits_xcpt1_pf_inst ? 4'hc : {{2'd0}, _T_7}; // @[Mux.scala 47:69]
  assign _T_9 = ibuf_io_inst_0_bits_xcpt0_ae_inst ? 4'h1 : _T_8; // @[Mux.scala 47:69]
  assign _T_10 = ibuf_io_inst_0_bits_xcpt0_pf_inst ? 4'hc : _T_9; // @[Mux.scala 47:69]
  assign _T_11 = bpu_io_xcpt_if ? 4'h3 : _T_10; // @[Mux.scala 47:69]
  assign _T_12 = bpu_io_debug_if ? 4'he : _T_11; // @[Mux.scala 47:69]
  assign ex_waddr = ex_reg_inst[11:7]; // @[RocketCore.scala 359:29]
  assign mem_waddr = mem_reg_inst[11:7]; // @[RocketCore.scala 360:31]
  assign wb_waddr = wb_reg_inst[11:7]; // @[RocketCore.scala 361:29]
  assign _T_23 = ex_reg_valid & ex_ctrl_wxd; // @[RocketCore.scala 364:19]
  assign _T_24 = mem_reg_valid & mem_ctrl_wxd; // @[RocketCore.scala 365:20]
  assign _T_26 = _T_24 & ~mem_ctrl_mem; // @[RocketCore.scala 365:36]
  assign id_bypass_src_0_0 = 5'h0 == id_raddr1; // @[RocketCore.scala 367:82]
  assign _id_bypass_src_T_1 = ex_waddr == id_raddr1; // @[RocketCore.scala 367:82]
  assign id_bypass_src_0_1 = _T_23 & _id_bypass_src_T_1; // @[RocketCore.scala 367:74]
  assign _id_bypass_src_T_2 = mem_waddr == id_raddr1; // @[RocketCore.scala 367:82]
  assign id_bypass_src_0_2 = _T_26 & _id_bypass_src_T_2; // @[RocketCore.scala 367:74]
  assign id_bypass_src_0_3 = _T_24 & _id_bypass_src_T_2; // @[RocketCore.scala 367:74]
  assign id_bypass_src_1_0 = 5'h0 == id_raddr2; // @[RocketCore.scala 367:82]
  assign _id_bypass_src_T_5 = ex_waddr == id_raddr2; // @[RocketCore.scala 367:82]
  assign id_bypass_src_1_1 = _T_23 & _id_bypass_src_T_5; // @[RocketCore.scala 367:74]
  assign _id_bypass_src_T_6 = mem_waddr == id_raddr2; // @[RocketCore.scala 367:82]
  assign id_bypass_src_1_2 = _T_26 & _id_bypass_src_T_6; // @[RocketCore.scala 367:74]
  assign id_bypass_src_1_3 = _T_24 & _id_bypass_src_T_6; // @[RocketCore.scala 367:74]
  assign _ex_rs_T = ex_reg_rs_lsb_0 == 2'h1; // @[package.scala 32:86]
  assign _ex_rs_T_1 = _ex_rs_T ? mem_reg_wdata : 64'h0; // @[package.scala 32:76]
  assign _ex_rs_T_2 = ex_reg_rs_lsb_0 == 2'h2; // @[package.scala 32:86]
  assign _ex_rs_T_3 = _ex_rs_T_2 ? wb_reg_wdata : _ex_rs_T_1; // @[package.scala 32:76]
  assign _ex_rs_T_4 = ex_reg_rs_lsb_0 == 2'h3; // @[package.scala 32:86]
  assign _ex_rs_T_5 = _ex_rs_T_4 ? io_dmem_resp_bits_data_word_bypass : _ex_rs_T_3; // @[package.scala 32:76]
  assign _ex_rs_T_6 = {ex_reg_rs_msb_0,ex_reg_rs_lsb_0}; // @[Cat.scala 30:58]
  assign _ex_rs_T_7 = ex_reg_rs_lsb_1 == 2'h1; // @[package.scala 32:86]
  assign _ex_rs_T_8 = _ex_rs_T_7 ? mem_reg_wdata : 64'h0; // @[package.scala 32:76]
  assign _ex_rs_T_9 = ex_reg_rs_lsb_1 == 2'h2; // @[package.scala 32:86]
  assign _ex_rs_T_10 = _ex_rs_T_9 ? wb_reg_wdata : _ex_rs_T_8; // @[package.scala 32:76]
  assign _ex_rs_T_11 = ex_reg_rs_lsb_1 == 2'h3; // @[package.scala 32:86]
  assign _ex_rs_T_12 = _ex_rs_T_11 ? io_dmem_resp_bits_data_word_bypass : _ex_rs_T_10; // @[package.scala 32:76]
  assign _ex_rs_T_13 = {ex_reg_rs_msb_1,ex_reg_rs_lsb_1}; // @[Cat.scala 30:58]
  assign ex_rs_1 = ex_reg_rs_bypass_1 ? _ex_rs_T_12 : _ex_rs_T_13; // @[RocketCore.scala 375:14]
  assign _ex_imm_sign_T = ex_ctrl_sel_imm == 3'h5; // @[RocketCore.scala 1037:24]
  assign _ex_imm_sign_T_2 = ex_reg_inst[31]; // @[RocketCore.scala 1037:53]
  assign ex_imm_sign = _ex_imm_sign_T ? $signed(1'sh0) : $signed(_ex_imm_sign_T_2); // @[RocketCore.scala 1037:19]
  assign _ex_imm_b30_20_T = ex_ctrl_sel_imm == 3'h2; // @[RocketCore.scala 1038:26]
  assign _ex_imm_b30_20_T_2 = ex_reg_inst[30:20]; // @[RocketCore.scala 1038:49]
  assign _ex_imm_b19_12_T = ex_ctrl_sel_imm != 3'h2; // @[RocketCore.scala 1039:26]
  assign _ex_imm_b19_12_T_1 = ex_ctrl_sel_imm != 3'h3; // @[RocketCore.scala 1039:43]
  assign _ex_imm_b19_12_T_2 = _ex_imm_b19_12_T & _ex_imm_b19_12_T_1; // @[RocketCore.scala 1039:36]
  assign _ex_imm_b19_12_T_4 = ex_reg_inst[19:12]; // @[RocketCore.scala 1039:73]
  assign _ex_imm_b11_T_2 = _ex_imm_b30_20_T | _ex_imm_sign_T; // @[RocketCore.scala 1040:33]
  assign _ex_imm_b11_T_3 = ex_ctrl_sel_imm == 3'h3; // @[RocketCore.scala 1041:23]
  assign _ex_imm_b11_T_5 = ex_reg_inst[20]; // @[RocketCore.scala 1041:44]
  assign _ex_imm_b11_T_6 = ex_ctrl_sel_imm == 3'h1; // @[RocketCore.scala 1042:23]
  assign _ex_imm_b11_T_8 = ex_reg_inst[7]; // @[RocketCore.scala 1042:43]
  assign _ex_imm_b11_T_9 = _ex_imm_b11_T_6 ? $signed(_ex_imm_b11_T_8) : $signed(ex_imm_sign); // @[RocketCore.scala 1042:18]
  assign _ex_imm_b11_T_10 = _ex_imm_b11_T_3 ? $signed(_ex_imm_b11_T_5) : $signed(_ex_imm_b11_T_9); // @[RocketCore.scala 1041:18]
  assign ex_imm_lo_hi_hi = _ex_imm_b11_T_2 ? 6'h0 : ex_reg_inst[30:25]; // @[RocketCore.scala 1043:20]
  assign _ex_imm_b4_1_T_1 = ex_ctrl_sel_imm == 3'h0; // @[RocketCore.scala 1045:24]
  assign _ex_imm_b4_1_T_3 = _ex_imm_b4_1_T_1 | _ex_imm_b11_T_6; // @[RocketCore.scala 1045:34]
  assign _ex_imm_b4_1_T_8 = _ex_imm_sign_T ? ex_reg_inst[19:16] : ex_reg_inst[24:21]; // @[RocketCore.scala 1046:19]
  assign _ex_imm_b4_1_T_9 = _ex_imm_b4_1_T_3 ? ex_reg_inst[11:8] : _ex_imm_b4_1_T_8; // @[RocketCore.scala 1045:19]
  assign ex_imm_lo_hi_lo = _ex_imm_b30_20_T ? 4'h0 : _ex_imm_b4_1_T_9; // @[RocketCore.scala 1044:19]
  assign _ex_imm_b0_T_2 = ex_ctrl_sel_imm == 3'h4; // @[RocketCore.scala 1048:22]
  assign _ex_imm_b0_T_6 = _ex_imm_sign_T & ex_reg_inst[15]; // @[RocketCore.scala 1049:17]
  assign _ex_imm_b0_T_7 = _ex_imm_b0_T_2 ? ex_reg_inst[20] : _ex_imm_b0_T_6; // @[RocketCore.scala 1048:17]
  assign ex_imm_lo_lo = _ex_imm_b4_1_T_1 ? ex_reg_inst[7] : _ex_imm_b0_T_7; // @[RocketCore.scala 1047:17]
  assign ex_imm_hi_lo_lo = _ex_imm_b11_T_2 ? $signed(1'sh0) : $signed(_ex_imm_b11_T_10); // @[Cat.scala 30:58]
  assign ex_imm_hi_lo_hi = _ex_imm_b19_12_T_2 ? $signed({8{ex_imm_sign}}) : $signed(_ex_imm_b19_12_T_4); // @[Cat.scala 30:58]
  assign ex_imm_hi_hi_lo = _ex_imm_b30_20_T ? $signed(_ex_imm_b30_20_T_2) : $signed({11{ex_imm_sign}}); // @[Cat.scala 30:58]
  assign ex_imm_hi_hi_hi = _ex_imm_sign_T ? $signed(1'sh0) : $signed(_ex_imm_sign_T_2); // @[Cat.scala 30:58]
  assign ex_imm = {ex_imm_hi_hi_hi,ex_imm_hi_hi_lo,ex_imm_hi_lo_hi,ex_imm_hi_lo_lo,ex_imm_lo_hi_hi,ex_imm_lo_hi_lo,ex_imm_lo_lo}; // @[RocketCore.scala 1051:53]
  assign _ex_op1_T = ex_reg_rs_bypass_0 ? _ex_rs_T_5 : _ex_rs_T_6; // @[RocketCore.scala 378:24]
  assign _ex_op1_T_2 = 2'h1 == ex_ctrl_sel_alu1; // @[Mux.scala 80:60]
  assign _ex_op1_T_3 = _ex_op1_T_2 ? $signed(_ex_op1_T) : $signed(64'sh0); // @[Mux.scala 80:57]
  assign _ex_op1_T_4 = 2'h2 == ex_ctrl_sel_alu1; // @[Mux.scala 80:60]
  assign _ex_op2_T = ex_reg_rs_bypass_1 ? _ex_rs_T_12 : _ex_rs_T_13; // @[RocketCore.scala 381:24]
  assign _ex_op2_T_1 = ex_reg_rvc ? $signed(4'sh2) : $signed(4'sh4); // @[RocketCore.scala 383:19]
  assign _ex_op2_T_2 = 2'h2 == ex_ctrl_sel_alu2; // @[Mux.scala 80:60]
  assign _ex_op2_T_3 = _ex_op2_T_2 ? $signed(_ex_op2_T) : $signed(64'sh0); // @[Mux.scala 80:57]
  assign _ex_op2_T_4 = 2'h3 == ex_ctrl_sel_alu2; // @[Mux.scala 80:60]
  assign _ex_op2_T_5 = _ex_op2_T_4 ? $signed({{32{ex_imm[31]}},ex_imm}) : $signed(_ex_op2_T_3); // @[Mux.scala 80:57]
  assign _ex_op2_T_6 = 2'h1 == ex_ctrl_sel_alu2; // @[Mux.scala 80:60]
  assign _ctrl_killd_T_1 = ~ibuf_io_inst_0_valid | ibuf_io_inst_0_bits_replay; // @[RocketCore.scala 784:40]
  assign _ctrl_killd_T_2 = _ctrl_killd_T_1 | take_pc_mem_wb; // @[RocketCore.scala 784:71]
  assign _T_123 = id_raddr1 != 5'h0; // @[RocketCore.scala 714:55]
  assign _T_124 = id_ctrl_decoder_7 & _T_123; // @[RocketCore.scala 714:42]
  assign _data_hazard_ex_T = id_raddr1 == ex_waddr; // @[RocketCore.scala 734:70]
  assign _data_hazard_ex_T_1 = _T_124 & _data_hazard_ex_T; // @[RocketCore.scala 984:27]
  assign _T_125 = id_raddr2 != 5'h0; // @[RocketCore.scala 715:55]
  assign _T_126 = id_ctrl_decoder_6 & _T_125; // @[RocketCore.scala 715:42]
  assign _data_hazard_ex_T_2 = id_raddr2 == ex_waddr; // @[RocketCore.scala 734:70]
  assign _data_hazard_ex_T_3 = _T_126 & _data_hazard_ex_T_2; // @[RocketCore.scala 984:27]
  assign _data_hazard_ex_T_6 = _data_hazard_ex_T_1 | _data_hazard_ex_T_3; // @[RocketCore.scala 984:50]
  assign _T_127 = id_waddr != 5'h0; // @[RocketCore.scala 716:55]
  assign _T_128 = id_ctrl_decoder_22 & _T_127; // @[RocketCore.scala 716:42]
  assign _data_hazard_ex_T_4 = id_waddr == ex_waddr; // @[RocketCore.scala 734:70]
  assign _data_hazard_ex_T_5 = _T_128 & _data_hazard_ex_T_4; // @[RocketCore.scala 984:27]
  assign _data_hazard_ex_T_7 = _data_hazard_ex_T_6 | _data_hazard_ex_T_5; // @[RocketCore.scala 984:50]
  assign data_hazard_ex = ex_ctrl_wxd & _data_hazard_ex_T_7; // @[RocketCore.scala 734:36]
  assign _ex_cannot_bypass_T = ex_ctrl_csr != 3'h0; // @[RocketCore.scala 733:38]
  assign _ex_cannot_bypass_T_1 = _ex_cannot_bypass_T | ex_ctrl_jalr; // @[RocketCore.scala 733:48]
  assign _ex_cannot_bypass_T_2 = _ex_cannot_bypass_T_1 | ex_ctrl_mem; // @[RocketCore.scala 733:64]
  assign _ex_cannot_bypass_T_4 = _ex_cannot_bypass_T_2 | ex_ctrl_div; // @[RocketCore.scala 733:94]
  assign ex_cannot_bypass = _ex_cannot_bypass_T_4 | ex_ctrl_fp; // @[RocketCore.scala 733:109]
  assign _id_ex_hazard_T = data_hazard_ex & ex_cannot_bypass; // @[RocketCore.scala 736:54]
  assign _fp_data_hazard_ex_T_1 = io_fpu_dec_ren1 & _data_hazard_ex_T; // @[RocketCore.scala 984:27]
  assign _fp_data_hazard_ex_T_3 = io_fpu_dec_ren2 & _data_hazard_ex_T_2; // @[RocketCore.scala 984:27]
  assign _fp_data_hazard_ex_T_8 = _fp_data_hazard_ex_T_1 | _fp_data_hazard_ex_T_3; // @[RocketCore.scala 984:50]
  assign _fp_data_hazard_ex_T_4 = id_raddr3 == ex_waddr; // @[RocketCore.scala 735:76]
  assign _fp_data_hazard_ex_T_5 = io_fpu_dec_ren3 & _fp_data_hazard_ex_T_4; // @[RocketCore.scala 984:27]
  assign _fp_data_hazard_ex_T_9 = _fp_data_hazard_ex_T_8 | _fp_data_hazard_ex_T_5; // @[RocketCore.scala 984:50]
  assign _fp_data_hazard_ex_T_7 = io_fpu_dec_wen & _data_hazard_ex_T_4; // @[RocketCore.scala 984:27]
  assign _fp_data_hazard_ex_T_10 = _fp_data_hazard_ex_T_9 | _fp_data_hazard_ex_T_7; // @[RocketCore.scala 984:50]
  assign fp_data_hazard_ex = ex_ctrl_wfd & _fp_data_hazard_ex_T_10; // @[RocketCore.scala 735:39]
  assign _id_ex_hazard_T_1 = _id_ex_hazard_T | fp_data_hazard_ex; // @[RocketCore.scala 736:74]
  assign id_ex_hazard = ex_reg_valid & _id_ex_hazard_T_1; // @[RocketCore.scala 736:35]
  assign _data_hazard_mem_T = id_raddr1 == mem_waddr; // @[RocketCore.scala 743:72]
  assign _data_hazard_mem_T_1 = _T_124 & _data_hazard_mem_T; // @[RocketCore.scala 984:27]
  assign _data_hazard_mem_T_2 = id_raddr2 == mem_waddr; // @[RocketCore.scala 743:72]
  assign _data_hazard_mem_T_3 = _T_126 & _data_hazard_mem_T_2; // @[RocketCore.scala 984:27]
  assign _data_hazard_mem_T_6 = _data_hazard_mem_T_1 | _data_hazard_mem_T_3; // @[RocketCore.scala 984:50]
  assign _data_hazard_mem_T_4 = id_waddr == mem_waddr; // @[RocketCore.scala 743:72]
  assign _data_hazard_mem_T_5 = _T_128 & _data_hazard_mem_T_4; // @[RocketCore.scala 984:27]
  assign _data_hazard_mem_T_7 = _data_hazard_mem_T_6 | _data_hazard_mem_T_5; // @[RocketCore.scala 984:50]
  assign data_hazard_mem = mem_ctrl_wxd & _data_hazard_mem_T_7; // @[RocketCore.scala 743:38]
  assign _mem_cannot_bypass_T = mem_ctrl_csr != 3'h0; // @[RocketCore.scala 742:40]
  assign _mem_cannot_bypass_T_1 = mem_ctrl_mem & mem_reg_slow_bypass; // @[RocketCore.scala 742:66]
  assign _mem_cannot_bypass_T_2 = _mem_cannot_bypass_T | _mem_cannot_bypass_T_1; // @[RocketCore.scala 742:50]
  assign _mem_cannot_bypass_T_4 = _mem_cannot_bypass_T_2 | mem_ctrl_div; // @[RocketCore.scala 742:100]
  assign mem_cannot_bypass = _mem_cannot_bypass_T_4 | mem_ctrl_fp; // @[RocketCore.scala 742:116]
  assign _id_mem_hazard_T = data_hazard_mem & mem_cannot_bypass; // @[RocketCore.scala 745:57]
  assign _fp_data_hazard_mem_T_1 = io_fpu_dec_ren1 & _data_hazard_mem_T; // @[RocketCore.scala 984:27]
  assign _fp_data_hazard_mem_T_3 = io_fpu_dec_ren2 & _data_hazard_mem_T_2; // @[RocketCore.scala 984:27]
  assign _fp_data_hazard_mem_T_8 = _fp_data_hazard_mem_T_1 | _fp_data_hazard_mem_T_3; // @[RocketCore.scala 984:50]
  assign _fp_data_hazard_mem_T_4 = id_raddr3 == mem_waddr; // @[RocketCore.scala 744:78]
  assign _fp_data_hazard_mem_T_5 = io_fpu_dec_ren3 & _fp_data_hazard_mem_T_4; // @[RocketCore.scala 984:27]
  assign _fp_data_hazard_mem_T_9 = _fp_data_hazard_mem_T_8 | _fp_data_hazard_mem_T_5; // @[RocketCore.scala 984:50]
  assign _fp_data_hazard_mem_T_7 = io_fpu_dec_wen & _data_hazard_mem_T_4; // @[RocketCore.scala 984:27]
  assign _fp_data_hazard_mem_T_10 = _fp_data_hazard_mem_T_9 | _fp_data_hazard_mem_T_7; // @[RocketCore.scala 984:50]
  assign fp_data_hazard_mem = mem_ctrl_wfd & _fp_data_hazard_mem_T_10; // @[RocketCore.scala 744:41]
  assign _id_mem_hazard_T_1 = _id_mem_hazard_T | fp_data_hazard_mem; // @[RocketCore.scala 745:78]
  assign id_mem_hazard = mem_reg_valid & _id_mem_hazard_T_1; // @[RocketCore.scala 745:37]
  assign _ctrl_stalld_T = id_ex_hazard | id_mem_hazard; // @[RocketCore.scala 772:18]
  assign _data_hazard_wb_T = id_raddr1 == wb_waddr; // @[RocketCore.scala 749:70]
  assign _data_hazard_wb_T_1 = _T_124 & _data_hazard_wb_T; // @[RocketCore.scala 984:27]
  assign _data_hazard_wb_T_2 = id_raddr2 == wb_waddr; // @[RocketCore.scala 749:70]
  assign _data_hazard_wb_T_3 = _T_126 & _data_hazard_wb_T_2; // @[RocketCore.scala 984:27]
  assign _data_hazard_wb_T_6 = _data_hazard_wb_T_1 | _data_hazard_wb_T_3; // @[RocketCore.scala 984:50]
  assign _data_hazard_wb_T_4 = id_waddr == wb_waddr; // @[RocketCore.scala 749:70]
  assign _data_hazard_wb_T_5 = _T_128 & _data_hazard_wb_T_4; // @[RocketCore.scala 984:27]
  assign _data_hazard_wb_T_7 = _data_hazard_wb_T_6 | _data_hazard_wb_T_5; // @[RocketCore.scala 984:50]
  assign data_hazard_wb = wb_ctrl_wxd & _data_hazard_wb_T_7; // @[RocketCore.scala 749:36]
  assign wb_dcache_miss = wb_ctrl_mem & ~io_dmem_resp_valid; // @[RocketCore.scala 491:36]
  assign wb_set_sboard = wb_ctrl_div | wb_dcache_miss; // @[RocketCore.scala 636:35]
  assign _id_wb_hazard_T = data_hazard_wb & wb_set_sboard; // @[RocketCore.scala 751:54]
  assign _fp_data_hazard_wb_T_1 = io_fpu_dec_ren1 & _data_hazard_wb_T; // @[RocketCore.scala 984:27]
  assign _fp_data_hazard_wb_T_3 = io_fpu_dec_ren2 & _data_hazard_wb_T_2; // @[RocketCore.scala 984:27]
  assign _fp_data_hazard_wb_T_8 = _fp_data_hazard_wb_T_1 | _fp_data_hazard_wb_T_3; // @[RocketCore.scala 984:50]
  assign _fp_data_hazard_wb_T_4 = id_raddr3 == wb_waddr; // @[RocketCore.scala 750:76]
  assign _fp_data_hazard_wb_T_5 = io_fpu_dec_ren3 & _fp_data_hazard_wb_T_4; // @[RocketCore.scala 984:27]
  assign _fp_data_hazard_wb_T_9 = _fp_data_hazard_wb_T_8 | _fp_data_hazard_wb_T_5; // @[RocketCore.scala 984:50]
  assign _fp_data_hazard_wb_T_7 = io_fpu_dec_wen & _data_hazard_wb_T_4; // @[RocketCore.scala 984:27]
  assign _fp_data_hazard_wb_T_10 = _fp_data_hazard_wb_T_9 | _fp_data_hazard_wb_T_7; // @[RocketCore.scala 984:50]
  assign fp_data_hazard_wb = wb_ctrl_wfd & _fp_data_hazard_wb_T_10; // @[RocketCore.scala 750:39]
  assign _id_wb_hazard_T_1 = _id_wb_hazard_T | fp_data_hazard_wb; // @[RocketCore.scala 751:71]
  assign id_wb_hazard = wb_reg_valid & _id_wb_hazard_T_1; // @[RocketCore.scala 751:35]
  assign _ctrl_stalld_T_1 = _ctrl_stalld_T | id_wb_hazard; // @[RocketCore.scala 772:35]
  assign r = {_r[31:1], 1'h0}; // @[RocketCore.scala 1002:40]
  assign _id_sboard_hazard_T = r >> id_raddr1; // @[RocketCore.scala 998:35]
  assign dmem_resp_valid = io_dmem_resp_valid & io_dmem_resp_bits_has_data; // @[RocketCore.scala 646:44]
  assign dmem_resp_replay = dmem_resp_valid & io_dmem_resp_bits_replay; // @[RocketCore.scala 647:42]
  assign dmem_resp_xpu = ~io_dmem_resp_bits_tag[0]; // @[RocketCore.scala 643:23]
  assign _T_117 = dmem_resp_replay & dmem_resp_xpu; // @[RocketCore.scala 662:26]
  assign ll_wen_x1 = div_io_resp_ready & div_io_resp_valid; // @[Decoupled.scala 40:37]
  assign ll_wen = _T_117 | ll_wen_x1; // @[RocketCore.scala 662:44]
  assign dmem_resp_waddr = io_dmem_resp_bits_tag[5:1]; // @[RocketCore.scala 645:46]
  assign ll_waddr = _T_117 ? dmem_resp_waddr : div_io_resp_bits_tag; // @[RocketCore.scala 662:44]
  assign _id_sboard_hazard_T_2 = ll_waddr == id_raddr1; // @[RocketCore.scala 726:70]
  assign _id_sboard_hazard_T_3 = ll_wen & _id_sboard_hazard_T_2; // @[RocketCore.scala 726:58]
  assign _id_sboard_hazard_T_5 = _id_sboard_hazard_T[0] & ~_id_sboard_hazard_T_3; // @[RocketCore.scala 729:77]
  assign _id_sboard_hazard_T_6 = _T_124 & _id_sboard_hazard_T_5; // @[RocketCore.scala 984:27]
  assign _id_sboard_hazard_T_7 = r >> id_raddr2; // @[RocketCore.scala 998:35]
  assign _id_sboard_hazard_T_9 = ll_waddr == id_raddr2; // @[RocketCore.scala 726:70]
  assign _id_sboard_hazard_T_10 = ll_wen & _id_sboard_hazard_T_9; // @[RocketCore.scala 726:58]
  assign _id_sboard_hazard_T_12 = _id_sboard_hazard_T_7[0] & ~_id_sboard_hazard_T_10; // @[RocketCore.scala 729:77]
  assign _id_sboard_hazard_T_13 = _T_126 & _id_sboard_hazard_T_12; // @[RocketCore.scala 984:27]
  assign _id_sboard_hazard_T_21 = _id_sboard_hazard_T_6 | _id_sboard_hazard_T_13; // @[RocketCore.scala 984:50]
  assign _id_sboard_hazard_T_14 = r >> id_waddr; // @[RocketCore.scala 998:35]
  assign _id_sboard_hazard_T_16 = ll_waddr == id_waddr; // @[RocketCore.scala 726:70]
  assign _id_sboard_hazard_T_17 = ll_wen & _id_sboard_hazard_T_16; // @[RocketCore.scala 726:58]
  assign _id_sboard_hazard_T_19 = _id_sboard_hazard_T_14[0] & ~_id_sboard_hazard_T_17; // @[RocketCore.scala 729:77]
  assign _id_sboard_hazard_T_20 = _T_128 & _id_sboard_hazard_T_19; // @[RocketCore.scala 984:27]
  assign id_sboard_hazard = _id_sboard_hazard_T_21 | _id_sboard_hazard_T_20; // @[RocketCore.scala 984:50]
  assign _ctrl_stalld_T_2 = _ctrl_stalld_T_1 | id_sboard_hazard; // @[RocketCore.scala 772:51]
  assign _ctrl_stalld_T_3 = ex_reg_valid | mem_reg_valid; // @[RocketCore.scala 773:40]
  assign _ctrl_stalld_T_4 = _ctrl_stalld_T_3 | wb_reg_valid; // @[RocketCore.scala 773:57]
  assign _ctrl_stalld_T_5 = csr_io_singleStep & _ctrl_stalld_T_4; // @[RocketCore.scala 773:23]
  assign _ctrl_stalld_T_6 = _ctrl_stalld_T_2 | _ctrl_stalld_T_5; // @[RocketCore.scala 772:71]
  assign _ctrl_stalld_T_7 = id_csr_en & csr_io_decode_0_fp_csr; // @[RocketCore.scala 774:15]
  assign _ctrl_stalld_T_9 = _ctrl_stalld_T_7 & ~io_fpu_fcsr_rdy; // @[RocketCore.scala 774:42]
  assign _ctrl_stalld_T_10 = _ctrl_stalld_T_6 | _ctrl_stalld_T_9; // @[RocketCore.scala 773:74]
  assign _id_stall_fpu_T_18 = id_stall_fpu__r >> id_raddr1; // @[RocketCore.scala 998:35]
  assign _id_stall_fpu_T_20 = io_fpu_dec_ren1 & _id_stall_fpu_T_18[0]; // @[RocketCore.scala 984:27]
  assign _id_stall_fpu_T_21 = id_stall_fpu__r >> id_raddr2; // @[RocketCore.scala 998:35]
  assign _id_stall_fpu_T_23 = io_fpu_dec_ren2 & _id_stall_fpu_T_21[0]; // @[RocketCore.scala 984:27]
  assign _id_stall_fpu_T_30 = _id_stall_fpu_T_20 | _id_stall_fpu_T_23; // @[RocketCore.scala 984:50]
  assign _id_stall_fpu_T_24 = id_stall_fpu__r >> id_raddr3; // @[RocketCore.scala 998:35]
  assign _id_stall_fpu_T_26 = io_fpu_dec_ren3 & _id_stall_fpu_T_24[0]; // @[RocketCore.scala 984:27]
  assign _id_stall_fpu_T_31 = _id_stall_fpu_T_30 | _id_stall_fpu_T_26; // @[RocketCore.scala 984:50]
  assign _id_stall_fpu_T_27 = id_stall_fpu__r >> id_waddr; // @[RocketCore.scala 998:35]
  assign _id_stall_fpu_T_29 = io_fpu_dec_wen & _id_stall_fpu_T_27[0]; // @[RocketCore.scala 984:27]
  assign id_stall_fpu = _id_stall_fpu_T_31 | _id_stall_fpu_T_29; // @[RocketCore.scala 984:50]
  assign _ctrl_stalld_T_11 = id_ctrl_decoder_1 & id_stall_fpu; // @[RocketCore.scala 775:16]
  assign _ctrl_stalld_T_12 = _ctrl_stalld_T_10 | _ctrl_stalld_T_11; // @[RocketCore.scala 774:62]
  assign dcache_blocked = blocked & ~io_dmem_perf_grant; // @[RocketCore.scala 766:13]
  assign _ctrl_stalld_T_13 = id_ctrl_decoder_14 & dcache_blocked; // @[RocketCore.scala 776:17]
  assign _ctrl_stalld_T_14 = _ctrl_stalld_T_12 | _ctrl_stalld_T_13; // @[RocketCore.scala 775:32]
  assign wb_wxd = wb_reg_valid & wb_ctrl_wxd; // @[RocketCore.scala 635:29]
  assign _ctrl_stalld_T_18 = div_io_resp_valid & ~wb_wxd; // @[RocketCore.scala 778:62]
  assign _ctrl_stalld_T_19 = div_io_req_ready | _ctrl_stalld_T_18; // @[RocketCore.scala 778:40]
  assign _ctrl_stalld_T_21 = ~_ctrl_stalld_T_19 | div_io_req_valid; // @[RocketCore.scala 778:75]
  assign _ctrl_stalld_T_22 = id_ctrl_decoder_21 & _ctrl_stalld_T_21; // @[RocketCore.scala 778:17]
  assign _ctrl_stalld_T_23 = _ctrl_stalld_T_14 | _ctrl_stalld_T_22; // @[RocketCore.scala 777:34]
  assign _ctrl_stalld_T_26 = _ctrl_stalld_T_23 | id_do_fence_x8; // @[RocketCore.scala 779:15]
  assign _ctrl_stalld_T_27 = _ctrl_stalld_T_26 | csr_io_csr_stall; // @[RocketCore.scala 780:17]
  assign ctrl_stalld = _ctrl_stalld_T_27 | id_reg_pause; // @[RocketCore.scala 781:22]
  assign _ctrl_killd_T_3 = _ctrl_killd_T_2 | ctrl_stalld; // @[RocketCore.scala 784:89]
  assign ctrl_killd = _ctrl_killd_T_3 | csr_io_interrupt; // @[RocketCore.scala 784:104]
  assign _ex_reg_replay_T_1 = ~take_pc_mem_wb & ibuf_io_inst_0_valid; // @[RocketCore.scala 424:29]
  assign _T_29 = id_fence_succ == 4'h0; // @[RocketCore.scala 434:42]
  assign _T_30 = id_ctrl_decoder_25 & _T_29; // @[RocketCore.scala 434:25]
  assign _GEN_1 = _T_30 | id_reg_pause; // @[RocketCore.scala 434:49]
  assign _GEN_2 = id_fence_next | _GEN_0; // @[RocketCore.scala 435:26]
  assign _T_31 = {ibuf_io_inst_0_bits_xcpt1_pf_inst,ibuf_io_inst_0_bits_xcpt1_ae_inst}; // @[RocketCore.scala 441:22]
  assign _T_32 = |_T_31; // @[RocketCore.scala 441:29]
  assign _GEN_5 = _T_32 | ibuf_io_inst_0_bits_rvc; // @[RocketCore.scala 441:34]
  assign _T_33 = {ibuf_io_inst_0_bits_xcpt0_pf_inst,ibuf_io_inst_0_bits_xcpt0_ae_inst}; // @[RocketCore.scala 446:40]
  assign _T_34 = |_T_33; // @[RocketCore.scala 446:47]
  assign _T_35 = bpu_io_xcpt_if | _T_34; // @[RocketCore.scala 446:28]
  assign _GEN_9 = id_xcpt | id_ctrl_decoder_12; // @[RocketCore.scala 436:20]
  assign _ex_reg_flush_pipe_T = id_ctrl_decoder_24 | id_csr_flush; // @[RocketCore.scala 451:42]
  assign _T_37 = id_ctrl_decoder_15 == 5'h5; // @[package.scala 15:47]
  assign _T_38 = _id_sfence_T | _T_37; // @[package.scala 72:59]
  assign _ex_reg_mem_size_T_1 = {_T_125,_T_123}; // @[Cat.scala 30:58]
  assign _do_bypass_T = id_bypass_src_0_0 | id_bypass_src_0_1; // @[RocketCore.scala 464:48]
  assign _do_bypass_T_1 = _do_bypass_T | id_bypass_src_0_2; // @[RocketCore.scala 464:48]
  assign do_bypass = _do_bypass_T_1 | id_bypass_src_0_3; // @[RocketCore.scala 464:48]
  assign _T_40 = id_ctrl_decoder_7 & ~do_bypass; // @[RocketCore.scala 468:23]
  assign _wb_valid_T_1 = wb_reg_valid & ~replay_wb_common; // @[RocketCore.scala 670:31]
  assign wb_valid = _wb_valid_T_1 & ~wb_xcpt; // @[RocketCore.scala 670:45]
  assign wb_wen = wb_valid & wb_ctrl_wxd; // @[RocketCore.scala 671:25]
  assign rf_wen = wb_wen | ll_wen; // @[RocketCore.scala 672:23]
  assign rf_waddr = ll_wen ? ll_waddr : wb_waddr; // @[RocketCore.scala 673:21]
  assign _T_118 = rf_waddr != 5'h0; // @[RocketCore.scala 1027:16]
  assign _T_121 = rf_waddr == id_raddr1; // @[RocketCore.scala 1030:20]
  assign _rf_wdata_T = dmem_resp_valid & dmem_resp_xpu; // @[RocketCore.scala 674:38]
  assign ll_wdata = div_io_resp_bits_data;
  assign _rf_wdata_T_2 = wb_ctrl_csr != 3'h0; // @[RocketCore.scala 676:34]
  assign _rf_wdata_T_4 = _rf_wdata_T_2 ? csr_io_rw_rdata : wb_reg_wdata; // @[RocketCore.scala 676:21]
  assign _rf_wdata_T_5 = ll_wen ? ll_wdata : _rf_wdata_T_4; // @[RocketCore.scala 675:21]
  assign rf_wdata = _rf_wdata_T ? io_dmem_resp_bits_data : _rf_wdata_T_5; // @[RocketCore.scala 674:21]
  assign _GEN_226 = _T_121 ? rf_wdata : _id_rs_T_4; // @[RocketCore.scala 1030:31]
  assign _GEN_233 = _T_118 ? _GEN_226 : _id_rs_T_4; // @[RocketCore.scala 1027:29]
  assign id_rs_0 = rf_wen ? _GEN_233 : _id_rs_T_4; // @[RocketCore.scala 679:17]
  assign _do_bypass_T_2 = id_bypass_src_1_0 | id_bypass_src_1_1; // @[RocketCore.scala 464:48]
  assign _do_bypass_T_3 = _do_bypass_T_2 | id_bypass_src_1_2; // @[RocketCore.scala 464:48]
  assign do_bypass_1 = _do_bypass_T_3 | id_bypass_src_1_3; // @[RocketCore.scala 464:48]
  assign _T_42 = id_ctrl_decoder_6 & ~do_bypass_1; // @[RocketCore.scala 468:23]
  assign _T_122 = rf_waddr == id_raddr2; // @[RocketCore.scala 1030:20]
  assign _GEN_227 = _T_122 ? rf_wdata : _id_rs_T_9; // @[RocketCore.scala 1030:31]
  assign _GEN_234 = _T_118 ? _GEN_227 : _id_rs_T_9; // @[RocketCore.scala 1027:29]
  assign id_rs_1 = rf_wen ? _GEN_234 : _id_rs_T_9; // @[RocketCore.scala 679:17]
  assign inst = ibuf_io_inst_0_bits_rvc ? {{16'd0}, ibuf_io_inst_0_bits_raw[15:0]} : ibuf_io_inst_0_bits_raw; // @[RocketCore.scala 474:21]
  assign _id_load_use_T = mem_reg_valid & data_hazard_mem; // @[RocketCore.scala 746:32]
  assign id_load_use = _id_load_use_T & mem_ctrl_mem; // @[RocketCore.scala 746:51]
  assign _T_44 = ~ctrl_killd | csr_io_interrupt; // @[RocketCore.scala 480:21]
  assign _T_45 = _T_44 | ibuf_io_inst_0_bits_replay; // @[RocketCore.scala 480:41]
  assign _replay_ex_structural_T_1 = ex_ctrl_mem & ~io_dmem_req_ready; // @[RocketCore.scala 492:42]
  assign _replay_ex_structural_T_3 = ex_ctrl_div & ~div_io_req_ready; // @[RocketCore.scala 493:42]
  assign replay_ex_structural = _replay_ex_structural_T_1 | _replay_ex_structural_T_3; // @[RocketCore.scala 492:64]
  assign replay_ex_load_use = wb_dcache_miss & ex_reg_load_use; // @[RocketCore.scala 494:43]
  assign _replay_ex_T = replay_ex_structural | replay_ex_load_use; // @[RocketCore.scala 495:75]
  assign _replay_ex_T_1 = ex_reg_valid & _replay_ex_T; // @[RocketCore.scala 495:50]
  assign replay_ex = ex_reg_replay | _replay_ex_T_1; // @[RocketCore.scala 495:33]
  assign _ctrl_killx_T = take_pc_mem_wb | replay_ex; // @[RocketCore.scala 496:35]
  assign ctrl_killx = _ctrl_killx_T | ~ex_reg_valid; // @[RocketCore.scala 496:48]
  assign _ex_slow_bypass_T = ex_ctrl_mem_cmd == 5'h7; // @[RocketCore.scala 498:40]
  assign _ex_slow_bypass_T_1 = ex_reg_mem_size < 2'h2; // @[RocketCore.scala 498:69]
  assign ex_slow_bypass = _ex_slow_bypass_T | _ex_slow_bypass_T_1; // @[RocketCore.scala 498:50]
  assign _ex_sfence_T_1 = ex_ctrl_mem_cmd == 5'h14; // @[RocketCore.scala 499:67]
  assign ex_sfence = ex_ctrl_mem & _ex_sfence_T_1; // @[RocketCore.scala 499:48]
  assign ex_xcpt = ex_reg_xcpt_interrupt | ex_reg_xcpt; // @[RocketCore.scala 502:28]
  assign _mem_pc_valid_T = mem_reg_valid | mem_reg_replay; // @[RocketCore.scala 508:36]
  assign mem_pc_valid = _mem_pc_valid_T | mem_reg_xcpt_interrupt; // @[RocketCore.scala 508:54]
  assign _mem_npc_misaligned_T_3 = ~csr_io_status_isa[2] & mem_npc[1]; // @[RocketCore.scala 517:56]
  assign mem_npc_misaligned = _mem_npc_misaligned_T_3 & ~mem_reg_sfence; // @[RocketCore.scala 517:70]
  assign _mem_int_wdata_T_1 = mem_ctrl_jalr ^ mem_npc_misaligned; // @[RocketCore.scala 518:59]
  assign _mem_int_wdata_T_2 = ~mem_reg_xcpt & _mem_int_wdata_T_1; // @[RocketCore.scala 518:41]
  assign mem_int_wdata = _mem_int_wdata_T_2 ? $signed({{24{mem_br_target[39]}},mem_br_target}) : $signed(mem_reg_wdata); // @[RocketCore.scala 518:119]
  assign _mem_cfi_T = mem_ctrl_branch | mem_ctrl_jalr; // @[RocketCore.scala 519:33]
  assign mem_cfi = _mem_cfi_T | mem_ctrl_jal; // @[RocketCore.scala 519:50]
  assign _mem_cfi_taken_T_1 = _mem_br_target_T_1 | mem_ctrl_jalr; // @[RocketCore.scala 520:57]
  assign mem_cfi_taken = _mem_cfi_taken_T_1 | mem_ctrl_jal; // @[RocketCore.scala 520:74]
  assign _T_56 = mem_reg_valid & mem_reg_flush_pipe; // @[RocketCore.scala 532:23]
  assign _mem_reg_load_T = ex_ctrl_mem_cmd == 5'h0; // @[Consts.scala 81:31]
  assign _mem_reg_load_T_1 = ex_ctrl_mem_cmd == 5'h6; // @[Consts.scala 81:48]
  assign _mem_reg_load_T_2 = _mem_reg_load_T | _mem_reg_load_T_1; // @[Consts.scala 81:41]
  assign _mem_reg_load_T_4 = _mem_reg_load_T_2 | _ex_slow_bypass_T; // @[Consts.scala 81:58]
  assign _mem_reg_load_T_5 = ex_ctrl_mem_cmd == 5'h4; // @[package.scala 15:47]
  assign _mem_reg_load_T_6 = ex_ctrl_mem_cmd == 5'h9; // @[package.scala 15:47]
  assign _mem_reg_load_T_7 = ex_ctrl_mem_cmd == 5'ha; // @[package.scala 15:47]
  assign _mem_reg_load_T_8 = ex_ctrl_mem_cmd == 5'hb; // @[package.scala 15:47]
  assign _mem_reg_load_T_9 = _mem_reg_load_T_5 | _mem_reg_load_T_6; // @[package.scala 72:59]
  assign _mem_reg_load_T_10 = _mem_reg_load_T_9 | _mem_reg_load_T_7; // @[package.scala 72:59]
  assign _mem_reg_load_T_11 = _mem_reg_load_T_10 | _mem_reg_load_T_8; // @[package.scala 72:59]
  assign _mem_reg_load_T_12 = ex_ctrl_mem_cmd == 5'h8; // @[package.scala 15:47]
  assign _mem_reg_load_T_13 = ex_ctrl_mem_cmd == 5'hc; // @[package.scala 15:47]
  assign _mem_reg_load_T_14 = ex_ctrl_mem_cmd == 5'hd; // @[package.scala 15:47]
  assign _mem_reg_load_T_15 = ex_ctrl_mem_cmd == 5'he; // @[package.scala 15:47]
  assign _mem_reg_load_T_16 = ex_ctrl_mem_cmd == 5'hf; // @[package.scala 15:47]
  assign _mem_reg_load_T_17 = _mem_reg_load_T_12 | _mem_reg_load_T_13; // @[package.scala 72:59]
  assign _mem_reg_load_T_18 = _mem_reg_load_T_17 | _mem_reg_load_T_14; // @[package.scala 72:59]
  assign _mem_reg_load_T_19 = _mem_reg_load_T_18 | _mem_reg_load_T_15; // @[package.scala 72:59]
  assign _mem_reg_load_T_20 = _mem_reg_load_T_19 | _mem_reg_load_T_16; // @[package.scala 72:59]
  assign _mem_reg_load_T_21 = _mem_reg_load_T_11 | _mem_reg_load_T_20; // @[Consts.scala 79:44]
  assign _mem_reg_load_T_22 = _mem_reg_load_T_4 | _mem_reg_load_T_21; // @[Consts.scala 81:75]
  assign _mem_reg_load_T_23 = ex_ctrl_mem & _mem_reg_load_T_22; // @[RocketCore.scala 539:33]
  assign _mem_reg_store_T = ex_ctrl_mem_cmd == 5'h1; // @[Consts.scala 82:32]
  assign _mem_reg_store_T_1 = ex_ctrl_mem_cmd == 5'h11; // @[Consts.scala 82:49]
  assign _mem_reg_store_T_2 = _mem_reg_store_T | _mem_reg_store_T_1; // @[Consts.scala 82:42]
  assign _mem_reg_store_T_4 = _mem_reg_store_T_2 | _ex_slow_bypass_T; // @[Consts.scala 82:59]
  assign _mem_reg_store_T_22 = _mem_reg_store_T_4 | _mem_reg_load_T_21; // @[Consts.scala 82:76]
  assign _mem_reg_store_T_23 = ex_ctrl_mem & _mem_reg_store_T_22; // @[RocketCore.scala 540:34]
  assign _mem_reg_wdata_T = alu_io_out; // @[RocketCore.scala 552:25]
  assign _T_58 = ex_ctrl_mem | ex_sfence; // @[RocketCore.scala 555:56]
  assign _T_59 = ex_ctrl_rxs2 & _T_58; // @[RocketCore.scala 555:24]
  assign _mem_reg_rs2_T = ex_reg_mem_size == 2'h0; // @[AMOALU.scala 26:19]
  assign mem_reg_rs2_hi = ex_rs_1[7:0]; // @[AMOALU.scala 26:66]
  assign _mem_reg_rs2_T_1 = {mem_reg_rs2_hi,mem_reg_rs2_hi,mem_reg_rs2_hi,mem_reg_rs2_hi,mem_reg_rs2_hi,mem_reg_rs2_hi,mem_reg_rs2_hi,mem_reg_rs2_hi}; // @[Cat.scala 30:58]
  assign _mem_reg_rs2_T_2 = ex_reg_mem_size == 2'h1; // @[AMOALU.scala 26:19]
  assign mem_reg_rs2_hi_3 = ex_rs_1[15:0]; // @[AMOALU.scala 26:66]
  assign _mem_reg_rs2_T_3 = {mem_reg_rs2_hi_3,mem_reg_rs2_hi_3,mem_reg_rs2_hi_3,mem_reg_rs2_hi_3}; // @[Cat.scala 30:58]
  assign _mem_reg_rs2_T_4 = ex_reg_mem_size == 2'h2; // @[AMOALU.scala 26:19]
  assign mem_reg_rs2_hi_5 = ex_rs_1[31:0]; // @[AMOALU.scala 26:66]
  assign _mem_reg_rs2_T_5 = {mem_reg_rs2_hi_5,mem_reg_rs2_hi_5}; // @[Cat.scala 30:58]
  assign _T_60 = ex_ctrl_jalr & csr_io_status_debug; // @[RocketCore.scala 559:24]
  assign _GEN_77 = _T_60 | ex_ctrl_fence_i; // @[RocketCore.scala 559:48]
  assign _GEN_78 = _T_60 | ex_reg_flush_pipe; // @[RocketCore.scala 559:48]
  assign _mem_breakpoint_T = mem_reg_load & bpu_io_xcpt_ld; // @[RocketCore.scala 566:38]
  assign _mem_breakpoint_T_1 = mem_reg_store & bpu_io_xcpt_st; // @[RocketCore.scala 566:75]
  assign mem_breakpoint = _mem_breakpoint_T | _mem_breakpoint_T_1; // @[RocketCore.scala 566:57]
  assign _mem_debug_breakpoint_T = mem_reg_load & bpu_io_debug_ld; // @[RocketCore.scala 567:44]
  assign _mem_debug_breakpoint_T_1 = mem_reg_store & bpu_io_debug_st; // @[RocketCore.scala 567:82]
  assign mem_debug_breakpoint = _mem_debug_breakpoint_T | _mem_debug_breakpoint_T_1; // @[RocketCore.scala 567:64]
  assign mem_ldst_xcpt = mem_debug_breakpoint | mem_breakpoint; // @[RocketCore.scala 975:26]
  assign mem_ldst_cause = mem_debug_breakpoint ? 4'he : 4'h3; // @[Mux.scala 47:69]
  assign _T_61 = mem_reg_xcpt_interrupt | mem_reg_xcpt; // @[RocketCore.scala 573:29]
  assign _T_62 = mem_reg_valid & mem_npc_misaligned; // @[RocketCore.scala 574:20]
  assign _T_63 = mem_reg_valid & mem_ldst_xcpt; // @[RocketCore.scala 575:20]
  assign _T_64 = _T_61 | _T_62; // @[RocketCore.scala 975:26]
  assign mem_xcpt = _T_64 | _T_63; // @[RocketCore.scala 975:26]
  assign _T_65 = _T_62 ? 4'h0 : mem_ldst_cause; // @[Mux.scala 47:69]
  assign dcache_kill_mem = _T_24 & io_dmem_replay_next; // @[RocketCore.scala 584:55]
  assign _fpu_kill_mem_T = mem_reg_valid & mem_ctrl_fp; // @[RocketCore.scala 585:36]
  assign fpu_kill_mem = _fpu_kill_mem_T & io_fpu_nack_mem; // @[RocketCore.scala 585:51]
  assign _replay_mem_T = dcache_kill_mem | mem_reg_replay; // @[RocketCore.scala 586:37]
  assign replay_mem = _replay_mem_T | fpu_kill_mem; // @[RocketCore.scala 586:55]
  assign _killm_common_T = dcache_kill_mem | take_pc_wb; // @[RocketCore.scala 587:38]
  assign _killm_common_T_1 = _killm_common_T | mem_reg_xcpt; // @[RocketCore.scala 587:52]
  assign killm_common = _killm_common_T_1 | ~mem_reg_valid; // @[RocketCore.scala 587:68]
  assign _ctrl_killm_T = killm_common | mem_xcpt; // @[RocketCore.scala 589:33]
  assign ctrl_killm = _ctrl_killm_T | fpu_kill_mem; // @[RocketCore.scala 589:45]
  assign _wb_reg_wdata_T_1 = ~mem_reg_xcpt & mem_ctrl_fp; // @[RocketCore.scala 600:25]
  assign _wb_reg_wdata_T_2 = _wb_reg_wdata_T_1 & mem_ctrl_wxd; // @[RocketCore.scala 600:40]
  assign _T_100 = _T_92 ? 3'h7 : 3'h5; // @[Mux.scala 47:69]
  assign _T_101 = _T_90 ? 4'hd : {{1'd0}, _T_100}; // @[Mux.scala 47:69]
  assign _T_102 = _T_88 ? 4'hf : _T_101; // @[Mux.scala 47:69]
  assign _T_103 = _T_86 ? 4'h4 : _T_102; // @[Mux.scala 47:69]
  assign _T_104 = _T_84 ? 4'h6 : _T_103; // @[Mux.scala 47:69]
  assign wb_cause = wb_reg_xcpt ? wb_reg_cause : {{60'd0}, _T_104}; // @[Mux.scala 47:69]
  assign _T_105 = wb_cause == 64'h6; // @[RocketCore.scala 979:38]
  assign _T_107 = wb_cause == 64'h4; // @[RocketCore.scala 979:38]
  assign _T_109 = wb_cause == 64'h7; // @[RocketCore.scala 979:38]
  assign _T_111 = wb_cause == 64'h5; // @[RocketCore.scala 979:38]
  assign _T_113 = wb_cause == 64'hf; // @[RocketCore.scala 979:38]
  assign _T_115 = wb_cause == 64'hd; // @[RocketCore.scala 979:38]
  assign _csr_io_inst_0_T_1 = &wb_reg_raw_inst[1:0]; // @[RocketCore.scala 687:73]
  assign csr_io_inst_0_hi = _csr_io_inst_0_T_1 ? wb_reg_inst[31:16] : 16'h0; // @[RocketCore.scala 687:50]
  assign csr_io_inst_0_lo = wb_reg_raw_inst[15:0]; // @[RocketCore.scala 687:119]
  assign _tval_valid_T = wb_cause == 64'h2; // @[package.scala 15:47]
  assign _tval_valid_T_1 = wb_cause == 64'h3; // @[package.scala 15:47]
  assign _tval_valid_T_6 = wb_cause == 64'h1; // @[package.scala 15:47]
  assign _tval_valid_T_9 = wb_cause == 64'hc; // @[package.scala 15:47]
  assign _tval_valid_T_10 = _tval_valid_T | _tval_valid_T_1; // @[package.scala 72:59]
  assign _tval_valid_T_11 = _tval_valid_T_10 | _T_107; // @[package.scala 72:59]
  assign _tval_valid_T_12 = _tval_valid_T_11 | _T_105; // @[package.scala 72:59]
  assign _tval_valid_T_13 = _tval_valid_T_12 | _T_111; // @[package.scala 72:59]
  assign _tval_valid_T_14 = _tval_valid_T_13 | _T_109; // @[package.scala 72:59]
  assign _tval_valid_T_15 = _tval_valid_T_14 | _tval_valid_T_6; // @[package.scala 72:59]
  assign _tval_valid_T_16 = _tval_valid_T_15 | _T_115; // @[package.scala 72:59]
  assign _tval_valid_T_17 = _tval_valid_T_16 | _T_113; // @[package.scala 72:59]
  assign _tval_valid_T_18 = _tval_valid_T_17 | _tval_valid_T_9; // @[package.scala 72:59]
  assign tval_valid = wb_xcpt & _tval_valid_T_18; // @[RocketCore.scala 696:28]
  assign a_1 = wb_reg_wdata[63:39]; // @[RocketCore.scala 989:23]
  assign _csr_io_tval_msb_T = $signed(a_1) == 25'sh0; // @[RocketCore.scala 990:21]
  assign _csr_io_tval_msb_T_1 = $signed(a_1) == -25'sh1; // @[RocketCore.scala 990:34]
  assign _csr_io_tval_msb_T_2 = _csr_io_tval_msb_T | _csr_io_tval_msb_T_1; // @[RocketCore.scala 990:29]
  assign msb_1 = _csr_io_tval_msb_T_2 ? wb_reg_wdata[39] : ~wb_reg_wdata[38]; // @[RocketCore.scala 990:18]
  assign csr_io_tval_lo = wb_reg_wdata[38:0]; // @[RocketCore.scala 991:16]
  assign _csr_io_tval_T = {msb_1,csr_io_tval_lo}; // @[Cat.scala 30:58]
  assign _csr_io_rw_cmd_T = wb_reg_valid ? 3'h0 : 3'h4; // @[CSR.scala 132:15]
  assign _T_129 = 32'h1 << ll_waddr; // @[RocketCore.scala 1005:62]
  assign _T_130 = ll_wen ? _T_129 : 32'h0; // @[RocketCore.scala 1005:49]
  assign _T_132 = r & ~_T_130; // @[RocketCore.scala 997:62]
  assign _T_134 = wb_set_sboard & wb_wen; // @[RocketCore.scala 730:28]
  assign _T_135 = 32'h1 << wb_waddr; // @[RocketCore.scala 1005:62]
  assign _T_136 = _T_134 ? _T_135 : 32'h0; // @[RocketCore.scala 1005:49]
  assign _T_137 = _T_132 | _T_136; // @[RocketCore.scala 996:60]
  assign _T_138 = ll_wen | _T_134; // @[RocketCore.scala 1008:17]
  assign _id_stall_fpu_T = wb_dcache_miss & wb_ctrl_wfd; // @[RocketCore.scala 755:35]
  assign _id_stall_fpu_T_1 = _id_stall_fpu_T | io_fpu_sboard_set; // @[RocketCore.scala 755:50]
  assign _id_stall_fpu_T_2 = _id_stall_fpu_T_1 & wb_valid; // @[RocketCore.scala 755:72]
  assign _id_stall_fpu_T_4 = _id_stall_fpu_T_2 ? _T_135 : 32'h0; // @[RocketCore.scala 1005:49]
  assign _id_stall_fpu_T_5 = id_stall_fpu__r | _id_stall_fpu_T_4; // @[RocketCore.scala 996:60]
  assign _id_stall_fpu_T_7 = dmem_resp_replay & io_dmem_resp_bits_tag[0]; // @[RocketCore.scala 756:38]
  assign _id_stall_fpu_T_8 = 32'h1 << dmem_resp_waddr; // @[RocketCore.scala 1005:62]
  assign _id_stall_fpu_T_9 = _id_stall_fpu_T_7 ? _id_stall_fpu_T_8 : 32'h0; // @[RocketCore.scala 1005:49]
  assign _id_stall_fpu_T_11 = _id_stall_fpu_T_5 & ~_id_stall_fpu_T_9; // @[RocketCore.scala 997:62]
  assign _id_stall_fpu_T_12 = _id_stall_fpu_T_2 | _id_stall_fpu_T_7; // @[RocketCore.scala 1008:17]
  assign _id_stall_fpu_T_13 = 32'h1 << io_fpu_sboard_clra; // @[RocketCore.scala 1005:62]
  assign _id_stall_fpu_T_14 = io_fpu_sboard_clr ? _id_stall_fpu_T_13 : 32'h0; // @[RocketCore.scala 1005:49]
  assign _id_stall_fpu_T_16 = _id_stall_fpu_T_11 & ~_id_stall_fpu_T_14; // @[RocketCore.scala 997:62]
  assign _id_stall_fpu_T_17 = _id_stall_fpu_T_12 | io_fpu_sboard_clr; // @[RocketCore.scala 1008:17]
  assign _dcache_blocked_blocked_T_3 = ~io_dmem_req_ready & ~io_dmem_perf_grant; // @[RocketCore.scala 765:60]
  assign _dcache_blocked_blocked_T_4 = blocked | io_dmem_req_valid; // @[RocketCore.scala 765:95]
  assign _dcache_blocked_blocked_T_5 = _dcache_blocked_blocked_T_4 | io_dmem_s2_nack; // @[RocketCore.scala 765:116]
  assign _io_imem_req_bits_pc_T = wb_xcpt | csr_io_eret; // @[RocketCore.scala 789:17]
  assign _io_imem_req_bits_pc_T_1 = replay_wb_common ? wb_reg_pc : mem_npc; // @[RocketCore.scala 790:8]
  assign _io_imem_flush_icache_T = wb_reg_valid & wb_ctrl_fence_i; // @[RocketCore.scala 792:40]
  assign _io_imem_might_request_imem_might_request_reg_T = ex_pc_valid | mem_pc_valid; // @[RocketCore.scala 794:43]
  assign _io_imem_btb_update_valid_T_1 = mem_reg_valid & ~take_pc_wb; // @[RocketCore.scala 806:45]
  assign _io_imem_btb_update_valid_T_2 = _io_imem_btb_update_valid_T_1 & mem_wrong_npc; // @[RocketCore.scala 806:60]
  assign _io_imem_btb_update_valid_T_4 = ~mem_cfi | mem_cfi_taken; // @[RocketCore.scala 806:90]
  assign _io_imem_btb_update_bits_cfiType_T = mem_ctrl_jal | mem_ctrl_jalr; // @[RocketCore.scala 809:23]
  assign _io_imem_btb_update_bits_cfiType_T_2 = _io_imem_btb_update_bits_cfiType_T & mem_waddr[0]; // @[RocketCore.scala 809:41]
  assign _io_imem_btb_update_bits_cfiType_T_5 = mem_reg_inst[19:15] & 5'h1b; // @[RocketCore.scala 810:62]
  assign _io_imem_btb_update_bits_cfiType_T_6 = 5'h1 == _io_imem_btb_update_bits_cfiType_T_5; // @[RocketCore.scala 810:62]
  assign _io_imem_btb_update_bits_cfiType_T_7 = mem_ctrl_jalr & _io_imem_btb_update_bits_cfiType_T_6; // @[RocketCore.scala 810:23]
  assign _io_imem_btb_update_bits_cfiType_T_10 = _io_imem_btb_update_bits_cfiType_T_7 ? 2'h3 : {{1'd0}, _io_imem_btb_update_bits_cfiType_T}; // @[RocketCore.scala 810:8]
  assign _io_imem_btb_update_bits_br_pc_T = mem_reg_rvc ? 2'h0 : 2'h2; // @[RocketCore.scala 814:74]
  assign _GEN_250 = {{38'd0}, _io_imem_btb_update_bits_br_pc_T}; // @[RocketCore.scala 814:69]
  assign _io_imem_btb_update_bits_br_pc_T_2 = mem_reg_pc + _GEN_250; // @[RocketCore.scala 814:69]
  assign _io_imem_btb_update_bits_pc_T_1 = ~io_imem_btb_update_bits_br_pc | 39'h3; // @[RocketCore.scala 815:66]
  assign ex_dcache_tag = {ex_waddr,ex_ctrl_fp}; // @[Cat.scala 30:58]
  assign a_2 = _ex_op1_T[63:39]; // @[RocketCore.scala 989:23]
  assign _io_dmem_req_bits_addr_msb_T = $signed(a_2) == 25'sh0; // @[RocketCore.scala 990:21]
  assign _io_dmem_req_bits_addr_msb_T_1 = $signed(a_2) == -25'sh1; // @[RocketCore.scala 990:34]
  assign _io_dmem_req_bits_addr_msb_T_2 = _io_dmem_req_bits_addr_msb_T | _io_dmem_req_bits_addr_msb_T_1; // @[RocketCore.scala 990:29]
  assign msb_2 = _io_dmem_req_bits_addr_msb_T_2 ? alu_io_adder_out[39] : ~alu_io_adder_out[38]; // @[RocketCore.scala 990:18]
  assign io_dmem_req_bits_addr_lo = alu_io_adder_out[38:0]; // @[RocketCore.scala 991:16]
  assign _io_dmem_s1_kill_T = killm_common | mem_ldst_xcpt; // @[RocketCore.scala 848:35]
  assign _unpause_T_1 = csr_io_time[4:0] == 5'h0; // @[RocketCore.scala 861:62]
  assign _unpause_T_2 = _unpause_T_1 | csr_io_inhibit_cycle; // @[RocketCore.scala 861:68]
  assign _unpause_T_3 = _unpause_T_2 | io_dmem_perf_release; // @[RocketCore.scala 861:92]
  assign unpause = _unpause_T_3 | take_pc_mem_wb; // @[RocketCore.scala 861:116]
  reg reg_coreMonitorBundle_valid; //SC
  assign reg_coreMonitorBundle_valid = coreMonitorBundle_valid;  
  assign coreMonitorBundle_valid = csr_io_trace_0_valid & ~csr_io_trace_0_exception; // @[RocketCore.scala 889:52]
  assign coreMonitorBundle_wrenx = wb_wen & ~wb_set_sboard; // @[RocketCore.scala 891:37]
  assign _GEN_251 = {{1'd0}, wb_waddr}; // @[RocketCore.scala 912:95]
  assign _T_142 = _GEN_251 + 6'h20; // @[RocketCore.scala 912:95]
  assign _T_145 = wb_waddr != 5'h0; // @[RocketCore.scala 914:28]
  assign _T_146 = wb_ctrl_wxd & _T_145; // @[RocketCore.scala 914:22]
  assign _T_147 = _T_146 & coreMonitorBundle_wrenx; // @[RocketCore.scala 914:40]
  assign _T_153 = _T_146 & ~coreMonitorBundle_wrenx; // @[RocketCore.scala 917:40]
  assign _T_159 = ll_wen & _T_118; // @[RocketCore.scala 925:18]
  assign io_imem_might_request = imem_might_request_reg; // @[RocketCore.scala 793:25]
  assign io_imem_req_valid = take_pc_wb | take_pc_mem; // @[RocketCore.scala 786:21]
  assign io_imem_req_bits_pc = _io_imem_req_bits_pc_T ? csr_io_evec : _io_imem_req_bits_pc_T_1; // @[RocketCore.scala 788:23]
  assign io_imem_req_bits_speculative = ~take_pc_wb; // @[RocketCore.scala 787:32]
  assign io_imem_sfence_valid = wb_reg_valid & wb_reg_sfence; // @[RocketCore.scala 797:24]
  assign io_imem_sfence_bits_rs1 = wb_reg_mem_size[0]; // @[RocketCore.scala 798:27]
  assign io_imem_sfence_bits_rs2 = wb_reg_mem_size[1]; // @[RocketCore.scala 799:27]
  assign io_imem_sfence_bits_addr = wb_reg_wdata[38:0]; // @[RocketCore.scala 800:28]
  assign io_imem_resp_ready = ibuf_io_imem_ready; // @[RocketCore.scala 258:16]
  assign io_imem_btb_update_valid = _io_imem_btb_update_valid_T_2 & _io_imem_btb_update_valid_T_4; // @[RocketCore.scala 806:28]
  assign io_imem_btb_update_bits_prediction_entry = mem_reg_btb_resp_entry; // @[RocketCore.scala 816:38]
  assign io_imem_btb_update_bits_pc = ~_io_imem_btb_update_bits_pc_T_1; // @[RocketCore.scala 815:30]
  assign io_imem_btb_update_bits_isValid = _mem_cfi_T | mem_ctrl_jal; // @[RocketCore.scala 807:35]
  assign io_imem_btb_update_bits_br_pc = _io_imem_btb_update_bits_br_pc_T_2[38:0]; // @[RocketCore.scala 814:33]
  assign io_imem_btb_update_bits_cfiType = _io_imem_btb_update_bits_cfiType_T_2 ? 2'h2 : _io_imem_btb_update_bits_cfiType_T_10; // @[RocketCore.scala 808:35]
  assign io_imem_bht_update_valid = mem_reg_valid & ~take_pc_wb; // @[RocketCore.scala 818:28]
  assign io_imem_bht_update_bits_prediction_history = mem_reg_btb_resp_bht_history; // @[RocketCore.scala 823:38]
  assign io_imem_bht_update_bits_pc = io_imem_btb_update_bits_pc; // @[RocketCore.scala 819:30]
  assign io_imem_bht_update_bits_branch = mem_ctrl_branch; // @[RocketCore.scala 822:34]
  assign io_imem_bht_update_bits_taken = mem_br_taken; // @[RocketCore.scala 820:33]
  assign io_imem_bht_update_bits_mispredict = ex_pc_valid ? _mem_wrong_npc_T : _mem_wrong_npc_T_3; // @[RocketCore.scala 821:38]
  assign io_imem_flush_icache = _io_imem_flush_icache_T & ~io_dmem_s2_nack; // @[RocketCore.scala 792:24]
  assign io_dmem_req_valid = ex_reg_valid & ex_ctrl_mem; // @[RocketCore.scala 836:25]
  assign io_dmem_req_bits_addr = {msb_2,io_dmem_req_bits_addr_lo}; // @[RocketCore.scala 844:25]
  assign io_dmem_req_bits_tag = {{1'd0}, ex_dcache_tag}; // @[RocketCore.scala 839:25]
  assign io_dmem_req_bits_cmd = ex_ctrl_mem_cmd; // @[RocketCore.scala 840:25]
  assign io_dmem_req_bits_size = ex_reg_mem_size; // @[RocketCore.scala 841:25]
  assign io_dmem_req_bits_signed = ~ex_reg_inst[14]; // @[RocketCore.scala 842:27]
  assign io_dmem_s1_kill = _io_dmem_s1_kill_T | fpu_kill_mem; // @[RocketCore.scala 848:19]
  assign io_dmem_s1_data_data = mem_ctrl_fp ? io_fpu_store_data : mem_reg_rs2; // @[RocketCore.scala 847:24]
  assign io_ptw_ptbr_mode = csr_io_ptbr_mode; // @[RocketCore.scala 701:15]
  assign io_ptw_ptbr_ppn = csr_io_ptbr_ppn; // @[RocketCore.scala 701:15]
  assign io_ptw_sfence_valid = io_imem_sfence_valid; // @[RocketCore.scala 802:17]
  assign io_ptw_sfence_bits_rs1 = io_imem_sfence_bits_rs1; // @[RocketCore.scala 802:17]
  assign io_ptw_status_debug = csr_io_status_debug; // @[RocketCore.scala 703:17]
  assign io_ptw_status_dprv = csr_io_status_dprv; // @[RocketCore.scala 703:17]
  assign io_ptw_status_prv = csr_io_status_prv; // @[RocketCore.scala 703:17]
  assign io_ptw_status_mxr = csr_io_status_mxr; // @[RocketCore.scala 703:17]
  assign io_ptw_status_sum = csr_io_status_sum; // @[RocketCore.scala 703:17]
  assign io_ptw_pmp_0_cfg_l = csr_io_pmp_0_cfg_l; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_0_cfg_a = csr_io_pmp_0_cfg_a; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_0_cfg_x = csr_io_pmp_0_cfg_x; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_0_cfg_w = csr_io_pmp_0_cfg_w; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_0_cfg_r = csr_io_pmp_0_cfg_r; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_0_addr = csr_io_pmp_0_addr; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_0_mask = csr_io_pmp_0_mask; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_1_cfg_l = csr_io_pmp_1_cfg_l; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_1_cfg_a = csr_io_pmp_1_cfg_a; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_1_cfg_x = csr_io_pmp_1_cfg_x; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_1_cfg_w = csr_io_pmp_1_cfg_w; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_1_cfg_r = csr_io_pmp_1_cfg_r; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_1_addr = csr_io_pmp_1_addr; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_1_mask = csr_io_pmp_1_mask; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_2_cfg_l = csr_io_pmp_2_cfg_l; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_2_cfg_a = csr_io_pmp_2_cfg_a; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_2_cfg_x = csr_io_pmp_2_cfg_x; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_2_cfg_w = csr_io_pmp_2_cfg_w; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_2_cfg_r = csr_io_pmp_2_cfg_r; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_2_addr = csr_io_pmp_2_addr; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_2_mask = csr_io_pmp_2_mask; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_3_cfg_l = csr_io_pmp_3_cfg_l; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_3_cfg_a = csr_io_pmp_3_cfg_a; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_3_cfg_x = csr_io_pmp_3_cfg_x; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_3_cfg_w = csr_io_pmp_3_cfg_w; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_3_cfg_r = csr_io_pmp_3_cfg_r; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_3_addr = csr_io_pmp_3_addr; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_3_mask = csr_io_pmp_3_mask; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_4_cfg_l = csr_io_pmp_4_cfg_l; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_4_cfg_a = csr_io_pmp_4_cfg_a; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_4_cfg_x = csr_io_pmp_4_cfg_x; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_4_cfg_w = csr_io_pmp_4_cfg_w; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_4_cfg_r = csr_io_pmp_4_cfg_r; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_4_addr = csr_io_pmp_4_addr; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_4_mask = csr_io_pmp_4_mask; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_5_cfg_l = csr_io_pmp_5_cfg_l; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_5_cfg_a = csr_io_pmp_5_cfg_a; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_5_cfg_x = csr_io_pmp_5_cfg_x; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_5_cfg_w = csr_io_pmp_5_cfg_w; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_5_cfg_r = csr_io_pmp_5_cfg_r; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_5_addr = csr_io_pmp_5_addr; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_5_mask = csr_io_pmp_5_mask; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_6_cfg_l = csr_io_pmp_6_cfg_l; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_6_cfg_a = csr_io_pmp_6_cfg_a; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_6_cfg_x = csr_io_pmp_6_cfg_x; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_6_cfg_w = csr_io_pmp_6_cfg_w; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_6_cfg_r = csr_io_pmp_6_cfg_r; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_6_addr = csr_io_pmp_6_addr; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_6_mask = csr_io_pmp_6_mask; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_7_cfg_l = csr_io_pmp_7_cfg_l; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_7_cfg_a = csr_io_pmp_7_cfg_a; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_7_cfg_x = csr_io_pmp_7_cfg_x; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_7_cfg_w = csr_io_pmp_7_cfg_w; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_7_cfg_r = csr_io_pmp_7_cfg_r; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_7_addr = csr_io_pmp_7_addr; // @[RocketCore.scala 704:14]
  assign io_ptw_pmp_7_mask = csr_io_pmp_7_mask; // @[RocketCore.scala 704:14]
  assign io_ptw_customCSRs_csrs_0_value = csr_io_customCSRs_0_value; // @[RocketCore.scala 702:79]
  assign io_fpu_inst = ibuf_io_inst_0_bits_inst_bits; // @[RocketCore.scala 828:15]
  assign io_fpu_fromint_data = ex_reg_rs_bypass_0 ? _ex_rs_T_5 : _ex_rs_T_6; // @[RocketCore.scala 829:23]
  assign io_fpu_fcsr_rm = csr_io_fcsr_rm; // @[RocketCore.scala 690:18]
  assign io_fpu_dmem_resp_val = dmem_resp_valid & io_dmem_resp_bits_tag[0]; // @[RocketCore.scala 830:24]
  assign io_fpu_dmem_resp_type = {{1'd0}, io_dmem_resp_bits_size}; // @[RocketCore.scala 832:25]
  assign io_fpu_dmem_resp_tag = io_dmem_resp_bits_tag[5:1]; // @[RocketCore.scala 833:24]
  assign io_fpu_dmem_resp_data = io_dmem_resp_bits_data_word_bypass; // @[RocketCore.scala 831:25]
  assign io_fpu_valid = ~ctrl_killd & id_ctrl_decoder_1; // @[RocketCore.scala 825:16]
  assign io_fpu_killx = _ctrl_killx_T | ~ex_reg_valid; // @[RocketCore.scala 826:16]
  assign io_fpu_killm = _killm_common_T_1 | ~mem_reg_valid; // @[RocketCore.scala 827:16]
  assign io_trace_0_valid = csr_io_trace_0_valid; // @[RocketCore.scala 708:12]
  assign io_trace_0_iaddr = csr_io_trace_0_iaddr; // @[RocketCore.scala 708:12]
  assign io_trace_0_insn = csr_io_trace_0_insn; // @[RocketCore.scala 708:12]
  assign io_trace_0_priv = csr_io_trace_0_priv; // @[RocketCore.scala 708:12]
  assign io_trace_0_exception = csr_io_trace_0_exception; // @[RocketCore.scala 708:12]
  assign io_trace_0_interrupt = csr_io_trace_0_interrupt; // @[RocketCore.scala 708:12]
  assign io_trace_0_cause = csr_io_trace_0_cause; // @[RocketCore.scala 708:12]
  assign io_trace_0_tval = csr_io_trace_0_tval; // @[RocketCore.scala 708:12]
  assign io_wfi = csr_io_status_wfi; // @[RocketCore.scala 864:10]
  assign ibuf_clock = clock;
  assign ibuf_reset = reset;
  assign ibuf_io_imem_valid = io_imem_resp_valid; // @[RocketCore.scala 258:16]
  assign ibuf_io_imem_bits_btb_taken = io_imem_resp_bits_btb_taken; // @[RocketCore.scala 258:16]
  assign ibuf_io_imem_bits_btb_bridx = io_imem_resp_bits_btb_bridx; // @[RocketCore.scala 258:16]
  assign ibuf_io_imem_bits_btb_entry = io_imem_resp_bits_btb_entry; // @[RocketCore.scala 258:16]
  assign ibuf_io_imem_bits_btb_bht_history = io_imem_resp_bits_btb_bht_history; // @[RocketCore.scala 258:16]
  assign ibuf_io_imem_bits_pc = io_imem_resp_bits_pc; // @[RocketCore.scala 258:16]
  assign ibuf_io_imem_bits_data = io_imem_resp_bits_data; // @[RocketCore.scala 258:16]
  assign ibuf_io_imem_bits_xcpt_pf_inst = io_imem_resp_bits_xcpt_pf_inst; // @[RocketCore.scala 258:16]
  assign ibuf_io_imem_bits_xcpt_ae_inst = io_imem_resp_bits_xcpt_ae_inst; // @[RocketCore.scala 258:16]
  assign ibuf_io_imem_bits_replay = io_imem_resp_bits_replay; // @[RocketCore.scala 258:16]
  assign ibuf_io_kill = take_pc_wb | take_pc_mem; // @[RocketCore.scala 259:16]
  assign ibuf_io_inst_0_ready = ~ctrl_stalld; // @[RocketCore.scala 804:25]
  assign csr_clock = clock;
  assign csr_reset = reset;
  assign csr_io_ungated_clock = clock; // @[RocketCore.scala 682:24]
  assign csr_io_interrupts_debug = io_interrupts_debug; // @[RocketCore.scala 688:21]
  assign csr_io_interrupts_mtip = io_interrupts_mtip; // @[RocketCore.scala 688:21]
  assign csr_io_interrupts_msip = io_interrupts_msip; // @[RocketCore.scala 688:21]
  assign csr_io_interrupts_meip = io_interrupts_meip; // @[RocketCore.scala 688:21]
  assign csr_io_interrupts_seip = io_interrupts_seip; // @[RocketCore.scala 688:21]
  assign csr_io_hartid = io_hartid; // @[RocketCore.scala 689:17]
  assign csr_io_rw_addr = wb_reg_inst[31:20]; // @[RocketCore.scala 705:18]
  assign csr_io_rw_cmd = wb_ctrl_csr & ~_csr_io_rw_cmd_T; // @[RocketCore.scala 706:17]
  assign csr_io_rw_wdata = wb_reg_wdata; // @[RocketCore.scala 707:19]
  assign csr_io_decode_0_csr = ibuf_io_inst_0_bits_raw[31:20]; // @[RocketCore.scala 683:24]
  assign csr_io_exception = _T_99 | _T_94; // @[RocketCore.scala 684:20]
  assign csr_io_retire = _wb_valid_T_1 & ~wb_xcpt; // @[RocketCore.scala 686:17]
  assign csr_io_cause = wb_reg_xcpt ? wb_reg_cause : {{60'd0}, _T_104}; // @[RocketCore.scala 685:16]
  assign csr_io_pc = wb_reg_pc; // @[RocketCore.scala 695:13]
  assign csr_io_tval = tval_valid ? _csr_io_tval_T : 40'h0; // @[RocketCore.scala 700:15]
  assign csr_io_fcsr_flags_valid = io_fpu_fcsr_flags_valid; // @[RocketCore.scala 691:21]
  assign csr_io_fcsr_flags_bits = io_fpu_fcsr_flags_bits; // @[RocketCore.scala 691:21]
  assign csr_io_inst_0 = {csr_io_inst_0_hi,csr_io_inst_0_lo}; // @[RocketCore.scala 687:18]
  assign bpu_io_status_debug = csr_io_status_debug; // @[RocketCore.scala 324:17]
  assign bpu_io_status_prv = csr_io_status_prv; // @[RocketCore.scala 324:17]
  assign bpu_io_bp_0_control_action = csr_io_bp_0_control_action; // @[RocketCore.scala 325:13]
  assign bpu_io_bp_0_control_tmatch = csr_io_bp_0_control_tmatch; // @[RocketCore.scala 325:13]
  assign bpu_io_bp_0_control_m = csr_io_bp_0_control_m; // @[RocketCore.scala 325:13]
  assign bpu_io_bp_0_control_s = csr_io_bp_0_control_s; // @[RocketCore.scala 325:13]
  assign bpu_io_bp_0_control_u = csr_io_bp_0_control_u; // @[RocketCore.scala 325:13]
  assign bpu_io_bp_0_control_x = csr_io_bp_0_control_x; // @[RocketCore.scala 325:13]
  assign bpu_io_bp_0_control_w = csr_io_bp_0_control_w; // @[RocketCore.scala 325:13]
  assign bpu_io_bp_0_control_r = csr_io_bp_0_control_r; // @[RocketCore.scala 325:13]
  assign bpu_io_bp_0_address = csr_io_bp_0_address; // @[RocketCore.scala 325:13]
  assign bpu_io_pc = ibuf_io_pc[38:0]; // @[RocketCore.scala 326:13]
  assign bpu_io_ea = mem_reg_wdata[38:0]; // @[RocketCore.scala 327:13]
  assign alu_io_dw = ex_ctrl_alu_dw; // @[RocketCore.scala 386:13]
  assign alu_io_fn = ex_ctrl_alu_fn; // @[RocketCore.scala 387:13]
  assign alu_io_in2 = _ex_op2_T_6 ? $signed({{60{_ex_op2_T_1[3]}},_ex_op2_T_1}) : $signed(_ex_op2_T_5); // @[RocketCore.scala 388:14]
  assign alu_io_in1 = _ex_op1_T_4 ? $signed({{24{ex_reg_pc[39]}},ex_reg_pc}) : $signed(_ex_op1_T_3); // @[RocketCore.scala 389:14]
  assign div_clock = clock;
  assign div_reset = reset;
  assign div_io_req_valid = ex_reg_valid & ex_ctrl_div; // @[RocketCore.scala 410:20]
  assign div_io_req_bits_fn = ex_ctrl_alu_fn; // @[RocketCore.scala 412:22]
  assign div_io_req_bits_dw = ex_ctrl_alu_dw; // @[RocketCore.scala 411:22]
  assign div_io_req_bits_in1 = ex_reg_rs_bypass_0 ? _ex_rs_T_5 : _ex_rs_T_6; // @[RocketCore.scala 413:23]
  assign div_io_req_bits_in2 = ex_reg_rs_bypass_1 ? _ex_rs_T_12 : _ex_rs_T_13; // @[RocketCore.scala 414:23]
  assign div_io_req_bits_tag = ex_reg_inst[11:7]; // @[RocketCore.scala 415:23]
  assign div_io_kill = killm_common & div_io_kill_REG; // @[RocketCore.scala 588:15]
  assign div_io_resp_ready = _T_117 ? 1'h0 : ~wb_wxd; // @[RocketCore.scala 649:21 RocketCore.scala 663:23]
  assign PlusArgTimeout_clock = clock;
  assign PlusArgTimeout_reset = reset;
  assign PlusArgTimeout_io_count = csr_io_time[31:0]; // @[PlusArg.scala 89:82]
  assign _GEN_254 = coreMonitorBundle_valid & wb_ctrl_wfd; // @[RocketCore.scala 912:16]
  assign _GEN_256 = coreMonitorBundle_valid & ~wb_ctrl_wfd; // @[RocketCore.scala 915:16]
  assign _GEN_257 = _GEN_256 & _T_147; // @[RocketCore.scala 915:16]
  assign _GEN_261 = _GEN_256 & ~_T_147; // @[RocketCore.scala 918:16]
  assign _GEN_262 = _GEN_261 & _T_153; // @[RocketCore.scala 918:16]
  assign _GEN_268 = _GEN_261 & ~_T_153; // @[RocketCore.scala 921:16]
  assign Rocket_cov_read_addr = Rocket_state;
  assign Rocket_cov_read_data = Rocket_cov[Rocket_cov_read_addr]; // @[Coverage map for Rocket]
  assign Rocket_cov_write_data = 1'h1;
  assign Rocket_cov_write_addr = Rocket_state;
  assign Rocket_cov_write_mask = 1'h1;
  assign Rocket_cov_write_en = 1'h1;
  assign mux_cond_0 = _T_122;
  assign mux_cond_1 = _csr_io_tval_msb_T_2;
  assign mux_cond_2 = _mem_npc_msb_T_2;
  assign mux_cond_3 = _csr_io_inst_0_T_1;
  assign mux_cond_4 = _T_118;
  assign mux_cond_5 = _T_121;
  assign ex_ctrl_wfd_shl = {ex_ctrl_wfd, 10'h0};
  assign ex_ctrl_wfd_pad = {9'h0,ex_ctrl_wfd_shl};
  assign ex_ctrl_fp_shl = {ex_ctrl_fp, 15'h0};
  assign ex_ctrl_fp_pad = {4'h0,ex_ctrl_fp_shl};
  assign mem_ctrl_jalr_shl = {mem_ctrl_jalr, 15'h0};
  assign mem_ctrl_jalr_pad = {4'h0,mem_ctrl_jalr_shl};
  assign wb_ctrl_mem_shl = {wb_ctrl_mem, 11'h0};
  assign wb_ctrl_mem_pad = {8'h0,wb_ctrl_mem_shl};
  assign ex_ctrl_wxd_shl = {ex_ctrl_wxd, 6'h0};
  assign ex_ctrl_wxd_pad = {13'h0,ex_ctrl_wxd_shl};
  assign ex_ctrl_mem_shl = {ex_ctrl_mem, 19'h0};
  assign ex_ctrl_mem_pad = ex_ctrl_mem_shl;
  assign ex_ctrl_sel_alu1_shl = {ex_ctrl_sel_alu1, 18'h0};
  assign ex_ctrl_sel_alu1_pad = ex_ctrl_sel_alu1_shl;
  assign mem_reg_replay_shl = {mem_reg_replay, 11'h0};
  assign mem_reg_replay_pad = {8'h0,mem_reg_replay_shl};
  assign blocked_shl = {blocked, 16'h0};
  assign blocked_pad = {3'h0,blocked_shl};
  assign wb_ctrl_div_shl = {wb_ctrl_div, 2'h0};
  assign wb_ctrl_div_pad = {17'h0,wb_ctrl_div_shl};
  assign wb_reg_flush_pipe_shl = {wb_reg_flush_pipe, 15'h0};
  assign wb_reg_flush_pipe_pad = {4'h0,wb_reg_flush_pipe_shl};
  assign mem_ctrl_jal_shl = {mem_ctrl_jal, 11'h0};
  assign mem_ctrl_jal_pad = {8'h0,mem_ctrl_jal_shl};
  assign ex_ctrl_sel_imm_shl = {ex_ctrl_sel_imm, 7'h0};
  assign ex_ctrl_sel_imm_pad = {10'h0,ex_ctrl_sel_imm_shl};
  assign wb_ctrl_wfd_shl = {wb_ctrl_wfd, 8'h0};
  assign wb_ctrl_wfd_pad = {11'h0,wb_ctrl_wfd_shl};
  assign mem_reg_slow_bypass_shl = {mem_reg_slow_bypass, 19'h0};
  assign mem_reg_slow_bypass_pad = mem_reg_slow_bypass_shl;
  assign mem_reg_sfence_shl = {mem_reg_sfence, 16'h0};
  assign mem_reg_sfence_pad = {3'h0,mem_reg_sfence_shl};
  assign wb_reg_xcpt_shl = {wb_reg_xcpt, 2'h0};
  assign wb_reg_xcpt_pad = {17'h0,wb_reg_xcpt_shl};
  assign id_reg_pause_shl = {id_reg_pause, 15'h0};
  assign id_reg_pause_pad = {4'h0,id_reg_pause_shl};
  assign ex_reg_rvc_shl = {ex_reg_rvc, 8'h0};
  assign ex_reg_rvc_pad = {11'h0,ex_reg_rvc_shl};
  assign wb_reg_valid_shl = {wb_reg_valid, 3'h0};
  assign wb_reg_valid_pad = {16'h0,wb_reg_valid_shl};
  assign mem_br_taken_shl = {mem_br_taken, 13'h0};
  assign mem_br_taken_pad = {6'h0,mem_br_taken_shl};
  assign mem_reg_flush_pipe_shl = {mem_reg_flush_pipe, 18'h0};
  assign mem_reg_flush_pipe_pad = {1'h0,mem_reg_flush_pipe_shl};
  assign ex_ctrl_div_shl = {ex_ctrl_div, 17'h0};
  assign ex_ctrl_div_pad = {2'h0,ex_ctrl_div_shl};
  assign mem_ctrl_fp_shl = {mem_ctrl_fp, 15'h0};
  assign mem_ctrl_fp_pad = {4'h0,mem_ctrl_fp_shl};
  assign mem_reg_xcpt_shl = {mem_reg_xcpt, 5'h0};
  assign mem_reg_xcpt_pad = {14'h0,mem_reg_xcpt_shl};
  assign mem_ctrl_wxd_shl = {mem_ctrl_wxd, 14'h0};
  assign mem_ctrl_wxd_pad = {5'h0,mem_ctrl_wxd_shl};
  assign mem_ctrl_mem_shl = {mem_ctrl_mem, 8'h0};
  assign mem_ctrl_mem_pad = {11'h0,mem_ctrl_mem_shl};
  assign ex_reg_mem_size_shl = {ex_reg_mem_size, 15'h0};
  assign ex_reg_mem_size_pad = {3'h0,ex_reg_mem_size_shl};
  assign ex_ctrl_sel_alu2_shl = {ex_ctrl_sel_alu2, 7'h0};
  assign ex_ctrl_sel_alu2_pad = {11'h0,ex_ctrl_sel_alu2_shl};
  assign ex_ctrl_rxs2_shl = {ex_ctrl_rxs2, 2'h0};
  assign ex_ctrl_rxs2_pad = {17'h0,ex_ctrl_rxs2_shl};
  assign ex_ctrl_jalr_shl = {ex_ctrl_jalr, 3'h0};
  assign ex_ctrl_jalr_pad = {16'h0,ex_ctrl_jalr_shl};
  assign ex_reg_replay_shl = {ex_reg_replay, 4'h0};
  assign ex_reg_replay_pad = {15'h0,ex_reg_replay_shl};
  assign ex_reg_valid_shl = {ex_reg_valid, 3'h0};
  assign ex_reg_valid_pad = {16'h0,ex_reg_valid_shl};
  assign mem_reg_valid_shl = {mem_reg_valid, 6'h0};
  assign mem_reg_valid_pad = {13'h0,mem_reg_valid_shl};
  assign mem_reg_rvc_shl = mem_reg_rvc;
  assign mem_reg_rvc_pad = {19'h0,mem_reg_rvc_shl};
  assign mem_ctrl_wfd_shl = mem_ctrl_wfd;
  assign mem_ctrl_wfd_pad = {19'h0,mem_ctrl_wfd_shl};
  assign id_reg_fence_shl = {id_reg_fence, 11'h0};
  assign id_reg_fence_pad = {8'h0,id_reg_fence_shl};
  assign mem_reg_load_shl = {mem_reg_load, 8'h0};
  assign mem_reg_load_pad = {11'h0,mem_reg_load_shl};
  assign wb_ctrl_wxd_shl = {wb_ctrl_wxd, 18'h0};
  assign wb_ctrl_wxd_pad = {1'h0,wb_ctrl_wxd_shl};
  assign wb_reg_replay_shl = {wb_reg_replay, 1'h0};
  assign wb_reg_replay_pad = {18'h0,wb_reg_replay_shl};
  assign ex_reg_xcpt_interrupt_shl = {ex_reg_xcpt_interrupt, 10'h0};
  assign ex_reg_xcpt_interrupt_pad = {9'h0,ex_reg_xcpt_interrupt_shl};
  assign mem_ctrl_branch_shl = {mem_ctrl_branch, 6'h0};
  assign mem_ctrl_branch_pad = {13'h0,mem_ctrl_branch_shl};
  assign mem_reg_xcpt_interrupt_shl = {mem_reg_xcpt_interrupt, 1'h0};
  assign mem_reg_xcpt_interrupt_pad = {18'h0,mem_reg_xcpt_interrupt_shl};
  assign mem_reg_store_shl = {mem_reg_store, 4'h0};
  assign mem_reg_store_pad = {15'h0,mem_reg_store_shl};
  assign mem_ctrl_div_shl = {mem_ctrl_div, 5'h0};
  assign mem_ctrl_div_pad = {14'h0,mem_ctrl_div_shl};
  assign mux_cond_0_shl = {mux_cond_0, 17'h0};
  assign mux_cond_0_pad = {2'h0,mux_cond_0_shl};
  assign mux_cond_1_shl = {mux_cond_1, 8'h0};
  assign mux_cond_1_pad = {11'h0,mux_cond_1_shl};
  assign mux_cond_2_shl = {mux_cond_2, 15'h0};
  assign mux_cond_2_pad = {4'h0,mux_cond_2_shl};
  assign mux_cond_3_shl = {mux_cond_3, 4'h0};
  assign mux_cond_3_pad = {15'h0,mux_cond_3_shl};
  assign mux_cond_4_shl = {mux_cond_4, 9'h0};
  assign mux_cond_4_pad = {10'h0,mux_cond_4_shl};
  assign mux_cond_5_shl = {mux_cond_5, 17'h0};
  assign mux_cond_5_pad = {2'h0,mux_cond_5_shl};
  assign ex_reg_rs_lsb_0_shl = {ex_reg_rs_lsb_0, 11'h0};
  assign ex_reg_rs_lsb_0_pad = {7'h0,ex_reg_rs_lsb_0_shl};
  assign ex_reg_rs_lsb_1_shl = {ex_reg_rs_lsb_1, 11'h0};
  assign ex_reg_rs_lsb_1_pad = {7'h0,ex_reg_rs_lsb_1_shl};
  assign ex_reg_rs_bypass_0_shl = {ex_reg_rs_bypass_0, 10'h0};
  assign ex_reg_rs_bypass_0_pad = {9'h0,ex_reg_rs_bypass_0_shl};
  assign ex_reg_rs_bypass_1_shl = {ex_reg_rs_bypass_1, 10'h0};
  assign ex_reg_rs_bypass_1_pad = {9'h0,ex_reg_rs_bypass_1_shl};
  assign Rocket_xor32 = ex_ctrl_fp_pad ^ mem_ctrl_jalr_pad;
  assign Rocket_xor15 = ex_ctrl_wfd_pad ^ Rocket_xor32;
  assign Rocket_xor34 = ex_ctrl_wxd_pad ^ ex_ctrl_mem_pad;
  assign Rocket_xor16 = wb_ctrl_mem_pad ^ Rocket_xor34;
  assign Rocket_xor7 = Rocket_xor15 ^ Rocket_xor16;
  assign Rocket_xor36 = mem_reg_replay_pad ^ blocked_pad;
  assign Rocket_xor17 = ex_ctrl_sel_alu1_pad ^ Rocket_xor36;
  assign Rocket_xor37 = wb_ctrl_div_pad ^ wb_reg_flush_pipe_pad;
  assign Rocket_xor38 = mem_ctrl_jal_pad ^ ex_ctrl_sel_imm_pad;
  assign Rocket_xor18 = Rocket_xor37 ^ Rocket_xor38;
  assign Rocket_xor8 = Rocket_xor17 ^ Rocket_xor18;
  assign Rocket_xor3 = Rocket_xor7 ^ Rocket_xor8;
  assign Rocket_xor40 = mem_reg_slow_bypass_pad ^ mem_reg_sfence_pad;
  assign Rocket_xor19 = wb_ctrl_wfd_pad ^ Rocket_xor40;
  assign Rocket_xor41 = wb_reg_xcpt_pad ^ id_reg_pause_pad;
  assign Rocket_xor42 = ex_reg_rvc_pad ^ wb_reg_valid_pad;
  assign Rocket_xor20 = Rocket_xor41 ^ Rocket_xor42;
  assign Rocket_xor9 = Rocket_xor19 ^ Rocket_xor20;
  assign Rocket_xor44 = mem_reg_flush_pipe_pad ^ ex_ctrl_div_pad;
  assign Rocket_xor21 = mem_br_taken_pad ^ Rocket_xor44;
  assign Rocket_xor45 = mem_ctrl_fp_pad ^ mem_reg_xcpt_pad;
  assign Rocket_xor46 = mem_ctrl_wxd_pad ^ mem_ctrl_mem_pad;
  assign Rocket_xor22 = Rocket_xor45 ^ Rocket_xor46;
  assign Rocket_xor10 = Rocket_xor21 ^ Rocket_xor22;
  assign Rocket_xor4 = Rocket_xor9 ^ Rocket_xor10;
  assign Rocket_xor1 = Rocket_xor3 ^ Rocket_xor4;
  assign Rocket_xor48 = ex_ctrl_sel_alu2_pad ^ ex_ctrl_rxs2_pad;
  assign Rocket_xor23 = ex_reg_mem_size_pad ^ Rocket_xor48;
  assign Rocket_xor49 = ex_ctrl_jalr_pad ^ ex_reg_replay_pad;
  assign Rocket_xor50 = ex_reg_valid_pad ^ mem_reg_valid_pad;
  assign Rocket_xor24 = Rocket_xor49 ^ Rocket_xor50;
  assign Rocket_xor11 = Rocket_xor23 ^ Rocket_xor24;
  assign Rocket_xor52 = mem_ctrl_wfd_pad ^ id_reg_fence_pad;
  assign Rocket_xor25 = mem_reg_rvc_pad ^ Rocket_xor52;
  assign Rocket_xor53 = mem_reg_load_pad ^ wb_ctrl_wxd_pad;
  assign Rocket_xor54 = wb_reg_replay_pad ^ ex_reg_xcpt_interrupt_pad;
  assign Rocket_xor26 = Rocket_xor53 ^ Rocket_xor54;
  assign Rocket_xor12 = Rocket_xor25 ^ Rocket_xor26;
  assign Rocket_xor5 = Rocket_xor11 ^ Rocket_xor12;
  assign Rocket_xor56 = mem_reg_xcpt_interrupt_pad ^ mem_reg_store_pad;
  assign Rocket_xor27 = mem_ctrl_branch_pad ^ Rocket_xor56;
  assign Rocket_xor57 = mem_ctrl_div_pad ^ mux_cond_0_pad;
  assign Rocket_xor58 = mux_cond_1_pad ^ mux_cond_2_pad;
  assign Rocket_xor28 = Rocket_xor57 ^ Rocket_xor58;
  assign Rocket_xor13 = Rocket_xor27 ^ Rocket_xor28;
  assign Rocket_xor60 = mux_cond_4_pad ^ mux_cond_5_pad;
  assign Rocket_xor29 = mux_cond_3_pad ^ Rocket_xor60;
  assign Rocket_xor61 = ex_reg_rs_lsb_0_pad ^ ex_reg_rs_lsb_1_pad;
  assign Rocket_xor62 = ex_reg_rs_bypass_0_pad ^ ex_reg_rs_bypass_1_pad;
  assign Rocket_xor30 = Rocket_xor61 ^ Rocket_xor62;
  assign Rocket_xor14 = Rocket_xor29 ^ Rocket_xor30;
  assign Rocket_xor6 = Rocket_xor13 ^ Rocket_xor14;
  assign Rocket_xor2 = Rocket_xor5 ^ Rocket_xor6;
  assign Rocket_xor0 = Rocket_xor1 ^ Rocket_xor2;
  assign PlusArgTimeout_sum = Rocket_covSum + PlusArgTimeout_io_covSum;
  assign csr_sum = PlusArgTimeout_sum + csr_io_covSum;
  assign bpu_sum = csr_sum + bpu_io_covSum;
  assign ibuf_sum = bpu_sum + ibuf_io_covSum;
  assign div_sum = ibuf_sum + div_io_covSum;
  assign alu_sum = div_sum + alu_io_covSum;
  assign io_covSum = alu_sum;
  assign alu_metaAssert_wire = alu_metaAssert;
  assign bpu_metaAssert_wire = bpu_metaAssert;
  assign PlusArgTimeout_metaAssert_wire = PlusArgTimeout_metaAssert;
  assign csr_metaAssert_wire = csr_metaAssert;
  assign ibuf_metaAssert_wire = ibuf_metaAssert;
  assign div_metaAssert_wire = div_metaAssert;
  assign Rocket_or4 = alu_metaAssert_wire | PlusArgTimeout_metaAssert_wire;
  assign Rocket_or1 = ibuf_metaAssert_wire | Rocket_or4;
  assign Rocket_or6 = div_metaAssert_wire | csr_metaAssert_wire;
  assign Rocket_or2 = bpu_metaAssert_wire | Rocket_or6;
  assign Rocket_or0 = Rocket_or1 | Rocket_or2;
  assign metaAssert = Rocket_metaAssert;
  assign PlusArgTimeout_metaReset = metaReset | PlusArgTimeout_halt;
  assign csr_metaReset = metaReset | csr_halt;
  assign ibuf_metaReset = metaReset | ibuf_halt;
  assign div_metaReset = metaReset | div_halt;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 31; initvar = initvar+1)
    rf[initvar] = _RAND_0[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {2{`RANDOM}};
  _RAND_2 = {2{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  id_reg_pause = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  imem_might_request_reg = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  ex_ctrl_fp = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  ex_ctrl_branch = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  ex_ctrl_jal = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  ex_ctrl_jalr = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  ex_ctrl_rxs2 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  ex_ctrl_sel_alu2 = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  ex_ctrl_sel_alu1 = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  ex_ctrl_sel_imm = _RAND_12[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  ex_ctrl_alu_dw = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  ex_ctrl_alu_fn = _RAND_14[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  ex_ctrl_mem = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  ex_ctrl_mem_cmd = _RAND_16[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  ex_ctrl_wfd = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  ex_ctrl_div = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  ex_ctrl_wxd = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  ex_ctrl_csr = _RAND_20[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  ex_ctrl_fence_i = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  mem_ctrl_fp = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  mem_ctrl_branch = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  mem_ctrl_jal = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  mem_ctrl_jalr = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  mem_ctrl_mem = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  mem_ctrl_wfd = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  mem_ctrl_div = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  mem_ctrl_wxd = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  mem_ctrl_csr = _RAND_30[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  mem_ctrl_fence_i = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  wb_ctrl_mem = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  wb_ctrl_wfd = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  wb_ctrl_div = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  wb_ctrl_wxd = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  wb_ctrl_csr = _RAND_36[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  wb_ctrl_fence_i = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  ex_reg_xcpt_interrupt = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  ex_reg_valid = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  ex_reg_rvc = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  ex_reg_btb_resp_entry = _RAND_41[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  ex_reg_btb_resp_bht_history = _RAND_42[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  ex_reg_xcpt = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  ex_reg_flush_pipe = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  ex_reg_load_use = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {2{`RANDOM}};
  ex_reg_cause = _RAND_46[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  ex_reg_replay = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {2{`RANDOM}};
  ex_reg_pc = _RAND_48[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  ex_reg_mem_size = _RAND_49[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  ex_reg_inst = _RAND_50[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  ex_reg_raw_inst = _RAND_51[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  mem_reg_xcpt_interrupt = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  mem_reg_valid = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  mem_reg_rvc = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  mem_reg_btb_resp_entry = _RAND_55[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  mem_reg_btb_resp_bht_history = _RAND_56[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  mem_reg_xcpt = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  mem_reg_replay = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  mem_reg_flush_pipe = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {2{`RANDOM}};
  mem_reg_cause = _RAND_60[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  mem_reg_slow_bypass = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  mem_reg_load = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  mem_reg_store = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  mem_reg_sfence = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {2{`RANDOM}};
  mem_reg_pc = _RAND_65[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  mem_reg_inst = _RAND_66[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  mem_reg_mem_size = _RAND_67[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  mem_reg_raw_inst = _RAND_68[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {2{`RANDOM}};
  mem_reg_wdata = _RAND_69[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {2{`RANDOM}};
  mem_reg_rs2 = _RAND_70[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  mem_br_taken = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  wb_reg_valid = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  wb_reg_xcpt = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  wb_reg_replay = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  wb_reg_flush_pipe = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {2{`RANDOM}};
  wb_reg_cause = _RAND_76[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  wb_reg_sfence = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {2{`RANDOM}};
  wb_reg_pc = _RAND_78[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  wb_reg_mem_size = _RAND_79[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  wb_reg_inst = _RAND_80[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  wb_reg_raw_inst = _RAND_81[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {2{`RANDOM}};
  wb_reg_wdata = _RAND_82[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  id_reg_fence = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  ex_reg_rs_bypass_0 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  ex_reg_rs_bypass_1 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  ex_reg_rs_lsb_0 = _RAND_86[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  ex_reg_rs_lsb_1 = _RAND_87[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {2{`RANDOM}};
  ex_reg_rs_msb_0 = _RAND_88[61:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {2{`RANDOM}};
  ex_reg_rs_msb_1 = _RAND_89[61:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _r = _RAND_90[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  id_stall_fpu__r = _RAND_91[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  blocked = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  div_io_kill_REG = _RAND_93[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  Rocket_state = _RAND_94[19:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1048576; initvar = initvar+1)
    Rocket_cov[initvar] = _RAND_95[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  Rocket_covSum = _RAND_96[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  Rocket_metaAssert = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(rf_MPORT_en & rf_MPORT_mask) begin
      rf[rf_MPORT_addr] <= rf_MPORT_data; // @[RocketCore.scala 1015:15]
    end
    if (metaReset) begin
      id_reg_pause <= 1'h0;
    end else if (unpause) begin
      id_reg_pause <= 1'h0;
    end else if (~ctrl_killd) begin
      id_reg_pause <= _GEN_1;
    end
    if (metaReset) begin
      imem_might_request_reg <= 1'h0;
    end else begin
      imem_might_request_reg <= _io_imem_might_request_imem_might_request_reg_T | io_ptw_customCSRs_csrs_0_value[1];
    end
    if (metaReset) begin
      ex_ctrl_fp <= 1'h0;
    end else if (~ctrl_killd) begin
      ex_ctrl_fp <= id_ctrl_decoder_1;
    end
    if (metaReset) begin
      ex_ctrl_branch <= 1'h0;
    end else if (~ctrl_killd) begin
      ex_ctrl_branch <= id_ctrl_decoder_3;
    end
    if (metaReset) begin
      ex_ctrl_jal <= 1'h0;
    end else if (~ctrl_killd) begin
      ex_ctrl_jal <= id_ctrl_decoder_4;
    end
    if (metaReset) begin
      ex_ctrl_jalr <= 1'h0;
    end else if (~ctrl_killd) begin
      ex_ctrl_jalr <= id_ctrl_decoder_5;
    end
    if (metaReset) begin
      ex_ctrl_rxs2 <= 1'h0;
    end else if (~ctrl_killd) begin
      ex_ctrl_rxs2 <= id_ctrl_decoder_6;
    end
    if (metaReset) begin
      ex_ctrl_sel_alu2 <= 2'h0;
    end else if (~ctrl_killd) begin
      if (id_xcpt) begin
        if (_T_35) begin
          ex_ctrl_sel_alu2 <= 2'h0;
        end else if (_T_32) begin
          ex_ctrl_sel_alu2 <= 2'h1;
        end else begin
          ex_ctrl_sel_alu2 <= 2'h0;
        end
      end else begin
        ex_ctrl_sel_alu2 <= id_ctrl_decoder_9;
      end
    end
    if (metaReset) begin
      ex_ctrl_sel_alu1 <= 2'h0;
    end else if (~ctrl_killd) begin
      if (id_xcpt) begin
        if (_T_35) begin
          ex_ctrl_sel_alu1 <= 2'h2;
        end else if (_T_32) begin
          ex_ctrl_sel_alu1 <= 2'h2;
        end else begin
          ex_ctrl_sel_alu1 <= 2'h1;
        end
      end else begin
        ex_ctrl_sel_alu1 <= id_ctrl_decoder_10;
      end
    end
    if (metaReset) begin
      ex_ctrl_sel_imm <= 3'h0;
    end else if (~ctrl_killd) begin
      ex_ctrl_sel_imm <= id_ctrl_decoder_11;
    end
    if (metaReset) begin
      ex_ctrl_alu_dw <= 1'h0;
    end else if (~ctrl_killd) begin
      ex_ctrl_alu_dw <= _GEN_9;
    end
    if (metaReset) begin
      ex_ctrl_alu_fn <= 4'h0;
    end else if (~ctrl_killd) begin
      if (id_xcpt) begin
        ex_ctrl_alu_fn <= 4'h0;
      end else begin
        ex_ctrl_alu_fn <= id_ctrl_decoder_13;
      end
    end
    if (metaReset) begin
      ex_ctrl_mem <= 1'h0;
    end else if (~ctrl_killd) begin
      ex_ctrl_mem <= id_ctrl_decoder_14;
    end
    if (metaReset) begin
      ex_ctrl_mem_cmd <= 5'h0;
    end else if (~ctrl_killd) begin
      ex_ctrl_mem_cmd <= id_ctrl_decoder_15;
    end
    if (metaReset) begin
      ex_ctrl_wfd <= 1'h0;
    end else if (~ctrl_killd) begin
      ex_ctrl_wfd <= id_ctrl_decoder_19;
    end
    if (metaReset) begin
      ex_ctrl_div <= 1'h0;
    end else if (~ctrl_killd) begin
      ex_ctrl_div <= id_ctrl_decoder_21;
    end
    if (metaReset) begin
      ex_ctrl_wxd <= 1'h0;
    end else if (~ctrl_killd) begin
      ex_ctrl_wxd <= id_ctrl_decoder_22;
    end
    if (metaReset) begin
      ex_ctrl_csr <= 3'h0;
    end else if (~ctrl_killd) begin
      if (id_csr_ren) begin
        ex_ctrl_csr <= 3'h2;
      end else begin
        ex_ctrl_csr <= id_ctrl_decoder_23;
      end
    end
    if (metaReset) begin
      ex_ctrl_fence_i <= 1'h0;
    end else if (~ctrl_killd) begin
      ex_ctrl_fence_i <= id_ctrl_decoder_24;
    end
    if (metaReset) begin
      mem_ctrl_fp <= 1'h0;
    end else if (!(_T_56)) begin
      if (ex_pc_valid) begin
        mem_ctrl_fp <= ex_ctrl_fp;
      end
    end
    if (metaReset) begin
      mem_ctrl_branch <= 1'h0;
    end else if (!(_T_56)) begin
      if (ex_pc_valid) begin
        mem_ctrl_branch <= ex_ctrl_branch;
      end
    end
    if (metaReset) begin
      mem_ctrl_jal <= 1'h0;
    end else if (!(_T_56)) begin
      if (ex_pc_valid) begin
        mem_ctrl_jal <= ex_ctrl_jal;
      end
    end
    if (metaReset) begin
      mem_ctrl_jalr <= 1'h0;
    end else if (!(_T_56)) begin
      if (ex_pc_valid) begin
        mem_ctrl_jalr <= ex_ctrl_jalr;
      end
    end
    if (metaReset) begin
      mem_ctrl_mem <= 1'h0;
    end else if (!(_T_56)) begin
      if (ex_pc_valid) begin
        mem_ctrl_mem <= ex_ctrl_mem;
      end
    end
    if (metaReset) begin
      mem_ctrl_wfd <= 1'h0;
    end else if (!(_T_56)) begin
      if (ex_pc_valid) begin
        mem_ctrl_wfd <= ex_ctrl_wfd;
      end
    end
    if (metaReset) begin
      mem_ctrl_div <= 1'h0;
    end else if (!(_T_56)) begin
      if (ex_pc_valid) begin
        mem_ctrl_div <= ex_ctrl_div;
      end
    end
    if (metaReset) begin
      mem_ctrl_wxd <= 1'h0;
    end else if (!(_T_56)) begin
      if (ex_pc_valid) begin
        mem_ctrl_wxd <= ex_ctrl_wxd;
      end
    end
    if (metaReset) begin
      mem_ctrl_csr <= 3'h0;
    end else if (!(_T_56)) begin
      if (ex_pc_valid) begin
        mem_ctrl_csr <= ex_ctrl_csr;
      end
    end
    if (metaReset) begin
      mem_ctrl_fence_i <= 1'h0;
    end else if (!(_T_56)) begin
      if (ex_pc_valid) begin
        mem_ctrl_fence_i <= _GEN_77;
      end
    end
    if (metaReset) begin
      wb_ctrl_mem <= 1'h0;
    end else if (mem_pc_valid) begin
      wb_ctrl_mem <= mem_ctrl_mem;
    end
    if (metaReset) begin
      wb_ctrl_wfd <= 1'h0;
    end else if (mem_pc_valid) begin
      wb_ctrl_wfd <= mem_ctrl_wfd;
    end
    if (metaReset) begin
      wb_ctrl_div <= 1'h0;
    end else if (mem_pc_valid) begin
      wb_ctrl_div <= mem_ctrl_div;
    end
    if (metaReset) begin
      wb_ctrl_wxd <= 1'h0;
    end else if (mem_pc_valid) begin
      wb_ctrl_wxd <= mem_ctrl_wxd;
    end
    if (metaReset) begin
      wb_ctrl_csr <= 3'h0;
    end else if (mem_pc_valid) begin
      wb_ctrl_csr <= mem_ctrl_csr;
    end
    if (metaReset) begin
      wb_ctrl_fence_i <= 1'h0;
    end else if (mem_pc_valid) begin
      wb_ctrl_fence_i <= mem_ctrl_fence_i;
    end
    if (metaReset) begin
      ex_reg_xcpt_interrupt <= 1'h0;
    end else begin
      ex_reg_xcpt_interrupt <= _ex_reg_replay_T_1 & csr_io_interrupt;
    end
    if (metaReset) begin
      ex_reg_valid <= 1'h0;
    end else begin
      ex_reg_valid <= ~ctrl_killd;
    end
    if (metaReset) begin
      ex_reg_rvc <= 1'h0;
    end else if (~ctrl_killd) begin
      if (id_xcpt) begin
        ex_reg_rvc <= _GEN_5;
      end else begin
        ex_reg_rvc <= ibuf_io_inst_0_bits_rvc;
      end
    end
    if (metaReset) begin
      ex_reg_btb_resp_entry <= 5'h0;
    end else if (_T_45) begin
      ex_reg_btb_resp_entry <= ibuf_io_btb_resp_entry;
    end
    if (metaReset) begin
      ex_reg_btb_resp_bht_history <= 8'h0;
    end else if (_T_45) begin
      ex_reg_btb_resp_bht_history <= ibuf_io_btb_resp_bht_history;
    end
    if (metaReset) begin
      ex_reg_xcpt <= 1'h0;
    end else begin
      ex_reg_xcpt <= ~ctrl_killd & id_xcpt;
    end
    if (metaReset) begin
      ex_reg_flush_pipe <= 1'h0;
    end else if (~ctrl_killd) begin
      ex_reg_flush_pipe <= _ex_reg_flush_pipe_T;
    end
    if (metaReset) begin
      ex_reg_load_use <= 1'h0;
    end else if (~ctrl_killd) begin
      ex_reg_load_use <= id_load_use;
    end
    if (metaReset) begin
      ex_reg_cause <= 64'h0;
    end else if (_T_45) begin
      if (csr_io_interrupt) begin
        ex_reg_cause <= csr_io_interrupt_cause;
      end else begin
        ex_reg_cause <= {{60'd0}, _T_12};
      end
    end
    if (metaReset) begin
      ex_reg_replay <= 1'h0;
    end else begin
      ex_reg_replay <= _ex_reg_replay_T_1 & ibuf_io_inst_0_bits_replay;
    end
    if (metaReset) begin
      ex_reg_pc <= 40'h0;
    end else if (_T_45) begin
      ex_reg_pc <= ibuf_io_pc;
    end
    if (metaReset) begin
      ex_reg_mem_size <= 2'h0;
    end else if (~ctrl_killd) begin
      if (_T_38) begin
        ex_reg_mem_size <= _ex_reg_mem_size_T_1;
      end else begin
        ex_reg_mem_size <= ibuf_io_inst_0_bits_inst_bits[13:12];
      end
    end
    if (metaReset) begin
      ex_reg_inst <= 32'h0;
    end else if (_T_45) begin
      ex_reg_inst <= ibuf_io_inst_0_bits_inst_bits;
    end
    if (metaReset) begin
      ex_reg_raw_inst <= 32'h0;
    end else if (_T_45) begin
      ex_reg_raw_inst <= ibuf_io_inst_0_bits_raw;
    end
    if (metaReset) begin
      mem_reg_xcpt_interrupt <= 1'h0;
    end else begin
      mem_reg_xcpt_interrupt <= ~take_pc_mem_wb & ex_reg_xcpt_interrupt;
    end
    if (metaReset) begin
      mem_reg_valid <= 1'h0;
    end else begin
      mem_reg_valid <= ~ctrl_killx;
    end
    if (metaReset) begin
      mem_reg_rvc <= 1'h0;
    end else if (!(_T_56)) begin
      if (ex_pc_valid) begin
        mem_reg_rvc <= ex_reg_rvc;
      end
    end
    if (metaReset) begin
      mem_reg_btb_resp_entry <= 5'h0;
    end else if (!(_T_56)) begin
      if (ex_pc_valid) begin
        mem_reg_btb_resp_entry <= ex_reg_btb_resp_entry;
      end
    end
    if (metaReset) begin
      mem_reg_btb_resp_bht_history <= 8'h0;
    end else if (!(_T_56)) begin
      if (ex_pc_valid) begin
        mem_reg_btb_resp_bht_history <= ex_reg_btb_resp_bht_history;
      end
    end
    if (metaReset) begin
      mem_reg_xcpt <= 1'h0;
    end else begin
      mem_reg_xcpt <= ~ctrl_killx & ex_xcpt;
    end
    if (metaReset) begin
      mem_reg_replay <= 1'h0;
    end else begin
      mem_reg_replay <= ~take_pc_mem_wb & replay_ex;
    end
    if (metaReset) begin
      mem_reg_flush_pipe <= 1'h0;
    end else if (!(_T_56)) begin
      if (ex_pc_valid) begin
        mem_reg_flush_pipe <= _GEN_78;
      end
    end
    if (metaReset) begin
      mem_reg_cause <= 64'h0;
    end else if (!(_T_56)) begin
      if (ex_pc_valid) begin
        mem_reg_cause <= ex_reg_cause;
      end
    end
    if (metaReset) begin
      mem_reg_slow_bypass <= 1'h0;
    end else if (!(_T_56)) begin
      if (ex_pc_valid) begin
        mem_reg_slow_bypass <= ex_slow_bypass;
      end
    end
    if (metaReset) begin
      mem_reg_load <= 1'h0;
    end else if (!(_T_56)) begin
      if (ex_pc_valid) begin
        mem_reg_load <= _mem_reg_load_T_23;
      end
    end
    if (metaReset) begin
      mem_reg_store <= 1'h0;
    end else if (!(_T_56)) begin
      if (ex_pc_valid) begin
        mem_reg_store <= _mem_reg_store_T_23;
      end
    end
    if (metaReset) begin
      mem_reg_sfence <= 1'h0;
    end else if (_T_56) begin
      mem_reg_sfence <= 1'h0;
    end else if (ex_pc_valid) begin
      mem_reg_sfence <= ex_sfence;
    end
    if (metaReset) begin
      mem_reg_pc <= 40'h0;
    end else if (!(_T_56)) begin
      if (ex_pc_valid) begin
        mem_reg_pc <= ex_reg_pc;
      end
    end
    if (metaReset) begin
      mem_reg_inst <= 32'h0;
    end else if (!(_T_56)) begin
      if (ex_pc_valid) begin
        mem_reg_inst <= ex_reg_inst;
      end
    end
    if (metaReset) begin
      mem_reg_mem_size <= 2'h0;
    end else if (!(_T_56)) begin
      if (ex_pc_valid) begin
        mem_reg_mem_size <= ex_reg_mem_size;
      end
    end
    if (metaReset) begin
      mem_reg_raw_inst <= 32'h0;
    end else if (!(_T_56)) begin
      if (ex_pc_valid) begin
        mem_reg_raw_inst <= ex_reg_raw_inst;
      end
    end
    if (metaReset) begin
      mem_reg_wdata <= 64'h0;
    end else if (!(_T_56)) begin
      if (ex_pc_valid) begin
        mem_reg_wdata <= _mem_reg_wdata_T;
      end
    end
    if (metaReset) begin
      mem_reg_rs2 <= 64'h0;
    end else if (!(_T_56)) begin
      if (ex_pc_valid) begin
        if (_T_59) begin
          if (_mem_reg_rs2_T) begin
            mem_reg_rs2 <= _mem_reg_rs2_T_1;
          end else if (_mem_reg_rs2_T_2) begin
            mem_reg_rs2 <= _mem_reg_rs2_T_3;
          end else if (_mem_reg_rs2_T_4) begin
            mem_reg_rs2 <= _mem_reg_rs2_T_5;
          end else if (ex_reg_rs_bypass_1) begin
            if (_ex_rs_T_11) begin
              mem_reg_rs2 <= io_dmem_resp_bits_data_word_bypass;
            end else if (_ex_rs_T_9) begin
              mem_reg_rs2 <= wb_reg_wdata;
            end else if (_ex_rs_T_7) begin
              mem_reg_rs2 <= mem_reg_wdata;
            end else begin
              mem_reg_rs2 <= 64'h0;
            end
          end else begin
            mem_reg_rs2 <= _ex_rs_T_13;
          end
        end
      end
    end
    if (metaReset) begin
      mem_br_taken <= 1'h0;
    end else if (!(_T_56)) begin
      if (ex_pc_valid) begin
        mem_br_taken <= alu_io_cmp_out;
      end
    end
    if (metaReset) begin
      wb_reg_valid <= 1'h0;
    end else begin
      wb_reg_valid <= ~ctrl_killm;
    end
    if (metaReset) begin
      wb_reg_xcpt <= 1'h0;
    end else begin
      wb_reg_xcpt <= mem_xcpt & ~take_pc_wb;
    end
    if (metaReset) begin
      wb_reg_replay <= 1'h0;
    end else begin
      wb_reg_replay <= replay_mem & ~take_pc_wb;
    end
    if (metaReset) begin
      wb_reg_flush_pipe <= 1'h0;
    end else begin
      wb_reg_flush_pipe <= ~ctrl_killm & mem_reg_flush_pipe;
    end
    if (metaReset) begin
      wb_reg_cause <= 64'h0;
    end else if (mem_pc_valid) begin
      if (_T_61) begin
        wb_reg_cause <= mem_reg_cause;
      end else begin
        wb_reg_cause <= {{60'd0}, _T_65};
      end
    end
    if (metaReset) begin
      wb_reg_sfence <= 1'h0;
    end else if (mem_pc_valid) begin
      wb_reg_sfence <= mem_reg_sfence;
    end
    if (metaReset) begin
      wb_reg_pc <= 40'h0;
    end else if (mem_pc_valid) begin
      wb_reg_pc <= mem_reg_pc;
    end
    if (metaReset) begin
      wb_reg_mem_size <= 2'h0;
    end else if (mem_pc_valid) begin
      wb_reg_mem_size <= mem_reg_mem_size;
    end
    if (metaReset) begin
      wb_reg_inst <= 32'h0;
    end else if (mem_pc_valid) begin
      wb_reg_inst <= mem_reg_inst;
    end
    if (metaReset) begin
      wb_reg_raw_inst <= 32'h0;
    end else if (mem_pc_valid) begin
      wb_reg_raw_inst <= mem_reg_raw_inst;
    end
    if (metaReset) begin
      wb_reg_wdata <= 64'h0;
    end else if (mem_pc_valid) begin
      if (_wb_reg_wdata_T_2) begin
        wb_reg_wdata <= io_fpu_toint_data;
      end else begin
        wb_reg_wdata <= mem_int_wdata;
      end
    end
    if (metaReset) begin
      id_reg_fence <= 1'h0;
    end else if (reset) begin
      id_reg_fence <= 1'h0;
    end else if (~ctrl_killd) begin
      id_reg_fence <= _GEN_2;
    end else if (~id_mem_busy) begin
      id_reg_fence <= 1'h0;
    end
    if (metaReset) begin
      ex_reg_rs_bypass_0 <= 1'h0;
    end else if (~ctrl_killd) begin
      if (id_illegal_insn) begin
        ex_reg_rs_bypass_0 <= 1'h0;
      end else begin
        ex_reg_rs_bypass_0 <= do_bypass;
      end
    end
    if (metaReset) begin
      ex_reg_rs_bypass_1 <= 1'h0;
    end else if (~ctrl_killd) begin
      ex_reg_rs_bypass_1 <= do_bypass_1;
    end
    if (metaReset) begin
      ex_reg_rs_lsb_0 <= 2'h0;
    end else if (~ctrl_killd) begin
      if (id_illegal_insn) begin
        ex_reg_rs_lsb_0 <= inst[1:0];
      end else if (_T_40) begin
        ex_reg_rs_lsb_0 <= id_rs_0[1:0];
      end else if (id_bypass_src_0_0) begin
        ex_reg_rs_lsb_0 <= 2'h0;
      end else if (id_bypass_src_0_1) begin
        ex_reg_rs_lsb_0 <= 2'h1;
      end else if (id_bypass_src_0_2) begin
        ex_reg_rs_lsb_0 <= 2'h2;
      end else begin
        ex_reg_rs_lsb_0 <= 2'h3;
      end
    end
    if (metaReset) begin
      ex_reg_rs_lsb_1 <= 2'h0;
    end else if (~ctrl_killd) begin
      if (_T_42) begin
        ex_reg_rs_lsb_1 <= id_rs_1[1:0];
      end else if (id_bypass_src_1_0) begin
        ex_reg_rs_lsb_1 <= 2'h0;
      end else if (id_bypass_src_1_1) begin
        ex_reg_rs_lsb_1 <= 2'h1;
      end else if (id_bypass_src_1_2) begin
        ex_reg_rs_lsb_1 <= 2'h2;
      end else begin
        ex_reg_rs_lsb_1 <= 2'h3;
      end
    end
    if (metaReset) begin
      ex_reg_rs_msb_0 <= 62'h0;
    end else if (~ctrl_killd) begin
      if (id_illegal_insn) begin
        ex_reg_rs_msb_0 <= {{32'd0}, inst[31:2]};
      end else if (_T_40) begin
        ex_reg_rs_msb_0 <= id_rs_0[63:2];
      end
    end
    if (metaReset) begin
      ex_reg_rs_msb_1 <= 62'h0;
    end else if (~ctrl_killd) begin
      if (_T_42) begin
        ex_reg_rs_msb_1 <= id_rs_1[63:2];
      end
    end
    if (metaReset) begin
      _r <= 32'h0;
    end else if (reset) begin
      _r <= 32'h0;
    end else if (_T_138) begin
      _r <= _T_137;
    end else if (ll_wen) begin
      _r <= _T_132;
    end
    if (metaReset) begin
      id_stall_fpu__r <= 32'h0;
    end else if (reset) begin
      id_stall_fpu__r <= 32'h0;
    end else if (_id_stall_fpu_T_17) begin
      id_stall_fpu__r <= _id_stall_fpu_T_16;
    end else if (_id_stall_fpu_T_12) begin
      id_stall_fpu__r <= _id_stall_fpu_T_11;
    end else if (_id_stall_fpu_T_2) begin
      id_stall_fpu__r <= _id_stall_fpu_T_5;
    end
    if (metaReset) begin
      blocked <= 1'h0;
    end else begin
      blocked <= _dcache_blocked_blocked_T_3 & _dcache_blocked_blocked_T_5;
    end
    if (metaReset) begin
      div_io_kill_REG <= 1'h0;
    end else begin
      div_io_kill_REG <= div_io_req_ready & div_io_req_valid;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_254 & ~reset) begin
          $fwrite(32'h80000002,"%d 0x%x (0x%x) f%d p%d 0xXXXXXXXXXXXXXXXX\n",csr_io_trace_0_priv,csr_io_trace_0_iaddr,csr_io_trace_0_insn,wb_waddr,_T_142); // @[RocketCore.scala 912:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_257 & ~reset) begin
          $fwrite(32'h80000002,"%d 0x%x (0x%x) x%d 0x%x\n",csr_io_trace_0_priv,csr_io_trace_0_iaddr,csr_io_trace_0_insn,wb_waddr,rf_wdata); // @[RocketCore.scala 915:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_262 & ~reset) begin
          $fwrite(32'h80000002,"%d 0x%x (0x%x) x%d p%d 0xXXXXXXXXXXXXXXXX\n",csr_io_trace_0_priv,csr_io_trace_0_iaddr,csr_io_trace_0_insn,wb_waddr,wb_waddr); // @[RocketCore.scala 918:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_268 & ~reset) begin
          $fwrite(32'h80000002,"%d 0x%x (0x%x)\n",csr_io_trace_0_priv,csr_io_trace_0_iaddr,csr_io_trace_0_insn); // @[RocketCore.scala 921:16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_159 & ~reset) begin
          $fwrite(32'h80000002,"x%d p%d 0x%x\n",rf_waddr,rf_waddr,rf_wdata); // @[RocketCore.scala 926:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    Rocket_state <= Rocket_xor0;
    if (!(Rocket_cov_read_data)) begin
      Rocket_covSum <= Rocket_covSum + 1'h1;
    end
    if (metaReset) begin
      Rocket_metaAssert <= 1'h0;
    end else begin
      Rocket_metaAssert <= Rocket_metaAssert | Rocket_or0;
    end
  end
  always @(posedge clock) begin
    if(Rocket_cov_write_en & Rocket_cov_write_mask) begin
      Rocket_cov[Rocket_cov_write_addr] <= Rocket_cov_write_data; // @[Coverage map for Rocket]
    end
  end
endmodule
module TLMonitor_23(
  input         clock,
  input         reset,
  input         io_in_a_ready,
  input         io_in_a_valid,
  input  [2:0]  io_in_a_bits_opcode,
  input  [2:0]  io_in_a_bits_param,
  input  [3:0]  io_in_a_bits_size,
  input         io_in_a_bits_source,
  input  [31:0] io_in_a_bits_address,
  input  [7:0]  io_in_a_bits_mask,
  input         io_in_b_ready,
  input         io_in_b_valid,
  input  [2:0]  io_in_b_bits_opcode,
  input  [1:0]  io_in_b_bits_param,
  input  [3:0]  io_in_b_bits_size,
  input         io_in_b_bits_source,
  input  [31:0] io_in_b_bits_address,
  input  [7:0]  io_in_b_bits_mask,
  input         io_in_b_bits_corrupt,
  input         io_in_c_ready,
  input         io_in_c_valid,
  input  [2:0]  io_in_c_bits_opcode,
  input  [2:0]  io_in_c_bits_param,
  input  [3:0]  io_in_c_bits_size,
  input         io_in_c_bits_source,
  input  [31:0] io_in_c_bits_address,
  input         io_in_d_ready,
  input         io_in_d_valid,
  input  [2:0]  io_in_d_bits_opcode,
  input  [1:0]  io_in_d_bits_param,
  input  [3:0]  io_in_d_bits_size,
  input         io_in_d_bits_source,
  input  [1:0]  io_in_d_bits_sink,
  input         io_in_d_bits_denied,
  input         io_in_d_bits_corrupt,
  input         io_in_e_ready,
  input         io_in_e_valid,
  input  [1:0]  io_in_e_bits_sink,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11]
  wire [31:0] plusarg_reader_1_out; // @[PlusArg.scala 80:11]
  wire  source_ok; // @[Parameters.scala 1125:46]
  wire [26:0] _is_aligned_mask_T_1; // @[package.scala 234:77]
  wire [11:0] is_aligned_mask; // @[package.scala 234:46]
  wire [31:0] _GEN_86; // @[Edges.scala 20:16]
  wire [31:0] _is_aligned_T; // @[Edges.scala 20:16]
  wire  is_aligned; // @[Edges.scala 20:24]
  wire [1:0] mask_sizeOH_shiftAmount; // @[OneHot.scala 64:49]
  wire [3:0] _mask_sizeOH_T_1; // @[OneHot.scala 65:12]
  wire [2:0] mask_sizeOH; // @[Misc.scala 201:81]
  wire  _mask_T; // @[Misc.scala 205:21]
  wire  mask_size; // @[Misc.scala 208:26]
  wire  mask_bit; // @[Misc.scala 209:26]
  wire  mask_nbit; // @[Misc.scala 210:20]
  wire  _mask_acc_T; // @[Misc.scala 214:38]
  wire  mask_acc; // @[Misc.scala 214:29]
  wire  _mask_acc_T_1; // @[Misc.scala 214:38]
  wire  mask_acc_1; // @[Misc.scala 214:29]
  wire  mask_size_1; // @[Misc.scala 208:26]
  wire  mask_bit_1; // @[Misc.scala 209:26]
  wire  mask_nbit_1; // @[Misc.scala 210:20]
  wire  mask_eq_2; // @[Misc.scala 213:27]
  wire  _mask_acc_T_2; // @[Misc.scala 214:38]
  wire  mask_acc_2; // @[Misc.scala 214:29]
  wire  mask_eq_3; // @[Misc.scala 213:27]
  wire  _mask_acc_T_3; // @[Misc.scala 214:38]
  wire  mask_acc_3; // @[Misc.scala 214:29]
  wire  mask_eq_4; // @[Misc.scala 213:27]
  wire  _mask_acc_T_4; // @[Misc.scala 214:38]
  wire  mask_acc_4; // @[Misc.scala 214:29]
  wire  mask_eq_5; // @[Misc.scala 213:27]
  wire  _mask_acc_T_5; // @[Misc.scala 214:38]
  wire  mask_acc_5; // @[Misc.scala 214:29]
  wire  mask_size_2; // @[Misc.scala 208:26]
  wire  mask_bit_2; // @[Misc.scala 209:26]
  wire  mask_nbit_2; // @[Misc.scala 210:20]
  wire  mask_eq_6; // @[Misc.scala 213:27]
  wire  _mask_acc_T_6; // @[Misc.scala 214:38]
  wire  mask_lo_lo_lo; // @[Misc.scala 214:29]
  wire  mask_eq_7; // @[Misc.scala 213:27]
  wire  _mask_acc_T_7; // @[Misc.scala 214:38]
  wire  mask_lo_lo_hi; // @[Misc.scala 214:29]
  wire  mask_eq_8; // @[Misc.scala 213:27]
  wire  _mask_acc_T_8; // @[Misc.scala 214:38]
  wire  mask_lo_hi_lo; // @[Misc.scala 214:29]
  wire  mask_eq_9; // @[Misc.scala 213:27]
  wire  _mask_acc_T_9; // @[Misc.scala 214:38]
  wire  mask_lo_hi_hi; // @[Misc.scala 214:29]
  wire  mask_eq_10; // @[Misc.scala 213:27]
  wire  _mask_acc_T_10; // @[Misc.scala 214:38]
  wire  mask_hi_lo_lo; // @[Misc.scala 214:29]
  wire  mask_eq_11; // @[Misc.scala 213:27]
  wire  _mask_acc_T_11; // @[Misc.scala 214:38]
  wire  mask_hi_lo_hi; // @[Misc.scala 214:29]
  wire  mask_eq_12; // @[Misc.scala 213:27]
  wire  _mask_acc_T_12; // @[Misc.scala 214:38]
  wire  mask_hi_hi_lo; // @[Misc.scala 214:29]
  wire  mask_eq_13; // @[Misc.scala 213:27]
  wire  _mask_acc_T_13; // @[Misc.scala 214:38]
  wire  mask_hi_hi_hi; // @[Misc.scala 214:29]
  wire [7:0] mask; // @[Cat.scala 30:58]
  wire [32:0] _T_7; // @[Parameters.scala 137:49]
  wire  _T_24; // @[Monitor.scala 81:25]
  wire  _T_26; // @[Parameters.scala 92:42]
  wire  _T_31; // @[Parameters.scala 1160:30]
  wire [32:0] _T_37; // @[Parameters.scala 137:52]
  wire  _T_38; // @[Parameters.scala 137:67]
  wire [31:0] _T_39; // @[Parameters.scala 137:31]
  wire [32:0] _T_40; // @[Parameters.scala 137:49]
  wire [32:0] _T_42; // @[Parameters.scala 137:52]
  wire  _T_43; // @[Parameters.scala 137:67]
  wire [31:0] _T_44; // @[Parameters.scala 137:31]
  wire [32:0] _T_45; // @[Parameters.scala 137:49]
  wire [32:0] _T_47; // @[Parameters.scala 137:52]
  wire  _T_48; // @[Parameters.scala 137:67]
  wire [31:0] _T_49; // @[Parameters.scala 137:31]
  wire [32:0] _T_50; // @[Parameters.scala 137:49]
  wire [32:0] _T_52; // @[Parameters.scala 137:52]
  wire  _T_53; // @[Parameters.scala 137:67]
  wire [31:0] _T_54; // @[Parameters.scala 137:31]
  wire [32:0] _T_55; // @[Parameters.scala 137:49]
  wire [32:0] _T_57; // @[Parameters.scala 137:52]
  wire  _T_58; // @[Parameters.scala 137:67]
  wire [31:0] _T_59; // @[Parameters.scala 137:31]
  wire [32:0] _T_60; // @[Parameters.scala 137:49]
  wire [32:0] _T_62; // @[Parameters.scala 137:52]
  wire  _T_63; // @[Parameters.scala 137:67]
  wire  _T_64; // @[Parameters.scala 671:42]
  wire  _T_65; // @[Parameters.scala 671:42]
  wire  _T_66; // @[Parameters.scala 671:42]
  wire  _T_67; // @[Parameters.scala 671:42]
  wire  _T_68; // @[Parameters.scala 671:42]
  wire  _T_71; // @[Parameters.scala 92:42]
  wire [31:0] _T_74; // @[Parameters.scala 137:31]
  wire [32:0] _T_75; // @[Parameters.scala 137:49]
  wire [32:0] _T_77; // @[Parameters.scala 137:52]
  wire  _T_78; // @[Parameters.scala 137:67]
  wire  _T_79; // @[Parameters.scala 670:56]
  wire  _T_82; // @[Monitor.scala 82:72]
  wire  _T_84; // @[Monitor.scala 42:11]
  wire  _T_88; // @[Parameters.scala 91:48]
  wire  _T_89; // @[Mux.scala 27:72]
  wire  _T_136; // @[Parameters.scala 671:42]
  wire  _T_137; // @[Parameters.scala 670:56]
  wire  _T_139; // @[Monitor.scala 83:78]
  wire  _T_141; // @[Monitor.scala 42:11]
  wire  _T_144; // @[Monitor.scala 42:11]
  wire  _T_148; // @[Monitor.scala 42:11]
  wire  _T_151; // @[Monitor.scala 42:11]
  wire  _T_153; // @[Bundles.scala 108:27]
  wire  _T_155; // @[Monitor.scala 42:11]
  wire  _T_158; // @[Monitor.scala 88:31]
  wire  _T_160; // @[Monitor.scala 42:11]
  wire  _T_166; // @[Monitor.scala 92:25]
  wire  _T_299; // @[Monitor.scala 99:31]
  wire  _T_301; // @[Monitor.scala 42:11]
  wire  _T_312; // @[Monitor.scala 104:25]
  wire  _T_322; // @[Monitor.scala 42:11]
  wire  _T_333; // @[Parameters.scala 670:56]
  wire  _T_368; // @[Parameters.scala 671:42]
  wire  _T_369; // @[Parameters.scala 671:42]
  wire  _T_370; // @[Parameters.scala 671:42]
  wire  _T_371; // @[Parameters.scala 671:42]
  wire  _T_372; // @[Parameters.scala 671:42]
  wire  _T_373; // @[Parameters.scala 670:56]
  wire  _T_375; // @[Parameters.scala 672:30]
  wire  _T_377; // @[Monitor.scala 42:11]
  wire  _T_385; // @[Monitor.scala 109:31]
  wire  _T_387; // @[Monitor.scala 42:11]
  wire  _T_389; // @[Monitor.scala 110:30]
  wire  _T_391; // @[Monitor.scala 42:11]
  wire  _T_397; // @[Monitor.scala 114:25]
  wire  _T_440; // @[Parameters.scala 671:42]
  wire  _T_441; // @[Parameters.scala 671:42]
  wire  _T_442; // @[Parameters.scala 671:42]
  wire  _T_443; // @[Parameters.scala 670:56]
  wire  _T_452; // @[Parameters.scala 92:42]
  wire  _T_460; // @[Parameters.scala 670:56]
  wire  _T_462; // @[Parameters.scala 672:30]
  wire  _T_464; // @[Parameters.scala 672:30]
  wire  _T_465; // @[Monitor.scala 115:71]
  wire  _T_467; // @[Monitor.scala 42:11]
  wire  _T_483; // @[Monitor.scala 122:25]
  wire [7:0] _T_566; // @[Monitor.scala 127:31]
  wire  _T_567; // @[Monitor.scala 127:40]
  wire  _T_569; // @[Monitor.scala 42:11]
  wire  _T_571; // @[Monitor.scala 130:25]
  wire  _T_581; // @[Parameters.scala 92:42]
  wire  _T_605; // @[Parameters.scala 671:42]
  wire  _T_606; // @[Parameters.scala 671:42]
  wire  _T_607; // @[Parameters.scala 670:56]
  wire  _T_629; // @[Monitor.scala 131:74]
  wire  _T_631; // @[Monitor.scala 42:11]
  wire  _T_639; // @[Bundles.scala 138:33]
  wire  _T_641; // @[Monitor.scala 42:11]
  wire  _T_647; // @[Monitor.scala 138:25]
  wire  _T_715; // @[Bundles.scala 145:30]
  wire  _T_717; // @[Monitor.scala 42:11]
  wire  _T_723; // @[Monitor.scala 146:25]
  wire  _T_781; // @[Monitor.scala 147:68]
  wire  _T_783; // @[Monitor.scala 42:11]
  wire  _T_791; // @[Bundles.scala 158:28]
  wire  _T_793; // @[Monitor.scala 42:11]
  wire  _T_803; // @[Bundles.scala 42:24]
  wire  _T_805; // @[Monitor.scala 49:11]
  wire  source_ok_1; // @[Parameters.scala 1125:46]
  wire  _T_807; // @[Monitor.scala 310:25]
  wire  _T_809; // @[Monitor.scala 49:11]
  wire  _T_811; // @[Monitor.scala 312:27]
  wire  _T_813; // @[Monitor.scala 49:11]
  wire  _T_815; // @[Monitor.scala 313:28]
  wire  _T_817; // @[Monitor.scala 49:11]
  wire  _T_821; // @[Monitor.scala 49:11]
  wire  _T_825; // @[Monitor.scala 49:11]
  wire  _T_827; // @[Monitor.scala 318:25]
  wire  _T_838; // @[Bundles.scala 102:26]
  wire  _T_840; // @[Monitor.scala 49:11]
  wire  _T_842; // @[Monitor.scala 323:28]
  wire  _T_844; // @[Monitor.scala 49:11]
  wire  _T_855; // @[Monitor.scala 328:25]
  wire  _T_875; // @[Monitor.scala 334:30]
  wire  _T_877; // @[Monitor.scala 49:11]
  wire  _T_884; // @[Monitor.scala 338:25]
  wire  _T_901; // @[Monitor.scala 346:25]
  wire  _T_919; // @[Monitor.scala 354:25]
  wire  _T_936; // @[Bundles.scala 40:24]
  wire  _T_938; // @[Monitor.scala 42:11]
  wire [32:0] _T_943; // @[Parameters.scala 137:49]
  wire [31:0] _address_ok_T; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_1; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_3; // @[Parameters.scala 137:52]
  wire  _address_ok_T_4; // @[Parameters.scala 137:67]
  wire [31:0] _address_ok_T_5; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_6; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_8; // @[Parameters.scala 137:52]
  wire  _address_ok_T_9; // @[Parameters.scala 137:67]
  wire [31:0] _address_ok_T_10; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_11; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_13; // @[Parameters.scala 137:52]
  wire  _address_ok_T_14; // @[Parameters.scala 137:67]
  wire [32:0] _address_ok_T_18; // @[Parameters.scala 137:52]
  wire  _address_ok_T_19; // @[Parameters.scala 137:67]
  wire [31:0] _address_ok_T_20; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_21; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_23; // @[Parameters.scala 137:52]
  wire  _address_ok_T_24; // @[Parameters.scala 137:67]
  wire [31:0] _address_ok_T_25; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_26; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_28; // @[Parameters.scala 137:52]
  wire  _address_ok_T_29; // @[Parameters.scala 137:67]
  wire [31:0] _address_ok_T_30; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_31; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_33; // @[Parameters.scala 137:52]
  wire  _address_ok_T_34; // @[Parameters.scala 137:67]
  wire  _address_ok_T_35; // @[Parameters.scala 622:64]
  wire  _address_ok_T_36; // @[Parameters.scala 622:64]
  wire  _address_ok_T_37; // @[Parameters.scala 622:64]
  wire  _address_ok_T_38; // @[Parameters.scala 622:64]
  wire  _address_ok_T_39; // @[Parameters.scala 622:64]
  wire  address_ok; // @[Parameters.scala 622:64]
  wire [26:0] _is_aligned_mask_T_4; // @[package.scala 234:77]
  wire [11:0] is_aligned_mask_1; // @[package.scala 234:46]
  wire [31:0] _GEN_87; // @[Edges.scala 20:16]
  wire [31:0] _is_aligned_T_1; // @[Edges.scala 20:16]
  wire  is_aligned_1; // @[Edges.scala 20:24]
  wire [1:0] mask_sizeOH_shiftAmount_1; // @[OneHot.scala 64:49]
  wire [3:0] _mask_sizeOH_T_4; // @[OneHot.scala 65:12]
  wire [2:0] mask_sizeOH_1; // @[Misc.scala 201:81]
  wire  _mask_T_1; // @[Misc.scala 205:21]
  wire  mask_size_3; // @[Misc.scala 208:26]
  wire  mask_bit_3; // @[Misc.scala 209:26]
  wire  mask_nbit_3; // @[Misc.scala 210:20]
  wire  _mask_acc_T_14; // @[Misc.scala 214:38]
  wire  mask_acc_6; // @[Misc.scala 214:29]
  wire  _mask_acc_T_15; // @[Misc.scala 214:38]
  wire  mask_acc_7; // @[Misc.scala 214:29]
  wire  mask_size_4; // @[Misc.scala 208:26]
  wire  mask_bit_4; // @[Misc.scala 209:26]
  wire  mask_nbit_4; // @[Misc.scala 210:20]
  wire  mask_eq_16; // @[Misc.scala 213:27]
  wire  _mask_acc_T_16; // @[Misc.scala 214:38]
  wire  mask_acc_8; // @[Misc.scala 214:29]
  wire  mask_eq_17; // @[Misc.scala 213:27]
  wire  _mask_acc_T_17; // @[Misc.scala 214:38]
  wire  mask_acc_9; // @[Misc.scala 214:29]
  wire  mask_eq_18; // @[Misc.scala 213:27]
  wire  _mask_acc_T_18; // @[Misc.scala 214:38]
  wire  mask_acc_10; // @[Misc.scala 214:29]
  wire  mask_eq_19; // @[Misc.scala 213:27]
  wire  _mask_acc_T_19; // @[Misc.scala 214:38]
  wire  mask_acc_11; // @[Misc.scala 214:29]
  wire  mask_size_5; // @[Misc.scala 208:26]
  wire  mask_bit_5; // @[Misc.scala 209:26]
  wire  mask_nbit_5; // @[Misc.scala 210:20]
  wire  mask_eq_20; // @[Misc.scala 213:27]
  wire  _mask_acc_T_20; // @[Misc.scala 214:38]
  wire  mask_lo_lo_lo_1; // @[Misc.scala 214:29]
  wire  mask_eq_21; // @[Misc.scala 213:27]
  wire  _mask_acc_T_21; // @[Misc.scala 214:38]
  wire  mask_lo_lo_hi_1; // @[Misc.scala 214:29]
  wire  mask_eq_22; // @[Misc.scala 213:27]
  wire  _mask_acc_T_22; // @[Misc.scala 214:38]
  wire  mask_lo_hi_lo_1; // @[Misc.scala 214:29]
  wire  mask_eq_23; // @[Misc.scala 213:27]
  wire  _mask_acc_T_23; // @[Misc.scala 214:38]
  wire  mask_lo_hi_hi_1; // @[Misc.scala 214:29]
  wire  mask_eq_24; // @[Misc.scala 213:27]
  wire  _mask_acc_T_24; // @[Misc.scala 214:38]
  wire  mask_hi_lo_lo_1; // @[Misc.scala 214:29]
  wire  mask_eq_25; // @[Misc.scala 213:27]
  wire  _mask_acc_T_25; // @[Misc.scala 214:38]
  wire  mask_hi_lo_hi_1; // @[Misc.scala 214:29]
  wire  mask_eq_26; // @[Misc.scala 213:27]
  wire  _mask_acc_T_26; // @[Misc.scala 214:38]
  wire  mask_hi_hi_lo_1; // @[Misc.scala 214:29]
  wire  mask_eq_27; // @[Misc.scala 213:27]
  wire  _mask_acc_T_27; // @[Misc.scala 214:38]
  wire  mask_hi_hi_hi_1; // @[Misc.scala 214:29]
  wire [7:0] mask_1; // @[Cat.scala 30:58]
  wire  legal_source; // @[Monitor.scala 165:113]
  wire  _T_960; // @[Monitor.scala 167:25]
  wire  _T_963; // @[Parameters.scala 91:48]
  wire  _T_964; // @[Mux.scala 27:72]
  wire  _T_968; // @[Parameters.scala 92:42]
  wire  _T_1006; // @[Parameters.scala 671:42]
  wire  _T_1007; // @[Parameters.scala 671:42]
  wire  _T_1008; // @[Parameters.scala 671:42]
  wire  _T_1009; // @[Parameters.scala 671:42]
  wire  _T_1010; // @[Parameters.scala 671:42]
  wire  _T_1011; // @[Parameters.scala 671:42]
  wire  _T_1012; // @[Parameters.scala 670:56]
  wire  _T_1014; // @[Monitor.scala 168:75]
  wire  _T_1016; // @[Monitor.scala 49:11]
  wire  _T_1019; // @[Monitor.scala 49:11]
  wire  _T_1022; // @[Monitor.scala 49:11]
  wire  _T_1025; // @[Monitor.scala 49:11]
  wire  _T_1027; // @[Bundles.scala 102:26]
  wire  _T_1029; // @[Monitor.scala 49:11]
  wire  _T_1031; // @[Monitor.scala 173:27]
  wire  _T_1033; // @[Monitor.scala 49:11]
  wire  _T_1037; // @[Monitor.scala 49:11]
  wire  _T_1039; // @[Monitor.scala 177:25]
  wire  _T_1100; // @[Monitor.scala 182:31]
  wire  _T_1102; // @[Monitor.scala 42:11]
  wire  _T_1112; // @[Monitor.scala 187:25]
  wire  _T_1181; // @[Monitor.scala 196:25]
  wire [7:0] _T_1247; // @[Monitor.scala 202:31]
  wire  _T_1248; // @[Monitor.scala 202:40]
  wire  _T_1250; // @[Monitor.scala 42:11]
  wire  _T_1252; // @[Monitor.scala 205:25]
  wire  _T_1321; // @[Monitor.scala 214:25]
  wire  _T_1390; // @[Monitor.scala 223:25]
  wire  source_ok_2; // @[Parameters.scala 1125:46]
  wire [26:0] _is_aligned_mask_T_7; // @[package.scala 234:77]
  wire [11:0] is_aligned_mask_2; // @[package.scala 234:46]
  wire [31:0] _GEN_88; // @[Edges.scala 20:16]
  wire [31:0] _is_aligned_T_2; // @[Edges.scala 20:16]
  wire  is_aligned_2; // @[Edges.scala 20:24]
  wire [31:0] _address_ok_T_40; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_41; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_43; // @[Parameters.scala 137:52]
  wire  _address_ok_T_44; // @[Parameters.scala 137:67]
  wire [31:0] _address_ok_T_45; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_46; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_48; // @[Parameters.scala 137:52]
  wire  _address_ok_T_49; // @[Parameters.scala 137:67]
  wire [31:0] _address_ok_T_50; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_51; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_53; // @[Parameters.scala 137:52]
  wire  _address_ok_T_54; // @[Parameters.scala 137:67]
  wire [32:0] _address_ok_T_56; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_58; // @[Parameters.scala 137:52]
  wire  _address_ok_T_59; // @[Parameters.scala 137:67]
  wire [31:0] _address_ok_T_60; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_61; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_63; // @[Parameters.scala 137:52]
  wire  _address_ok_T_64; // @[Parameters.scala 137:67]
  wire [31:0] _address_ok_T_65; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_66; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_68; // @[Parameters.scala 137:52]
  wire  _address_ok_T_69; // @[Parameters.scala 137:67]
  wire [31:0] _address_ok_T_70; // @[Parameters.scala 137:31]
  wire [32:0] _address_ok_T_71; // @[Parameters.scala 137:49]
  wire [32:0] _address_ok_T_73; // @[Parameters.scala 137:52]
  wire  _address_ok_T_74; // @[Parameters.scala 137:67]
  wire  _address_ok_T_75; // @[Parameters.scala 622:64]
  wire  _address_ok_T_76; // @[Parameters.scala 622:64]
  wire  _address_ok_T_77; // @[Parameters.scala 622:64]
  wire  _address_ok_T_78; // @[Parameters.scala 622:64]
  wire  _address_ok_T_79; // @[Parameters.scala 622:64]
  wire  address_ok_1; // @[Parameters.scala 622:64]
  wire  _T_1483; // @[Monitor.scala 242:25]
  wire  _T_1485; // @[Monitor.scala 42:11]
  wire  _T_1488; // @[Monitor.scala 42:11]
  wire  _T_1490; // @[Monitor.scala 245:30]
  wire  _T_1492; // @[Monitor.scala 42:11]
  wire  _T_1495; // @[Monitor.scala 42:11]
  wire  _T_1497; // @[Bundles.scala 120:29]
  wire  _T_1499; // @[Monitor.scala 42:11]
  wire  _T_1505; // @[Monitor.scala 251:25]
  wire  _T_1523; // @[Monitor.scala 259:25]
  wire  _T_1525; // @[Parameters.scala 92:42]
  wire  _T_1530; // @[Parameters.scala 1160:30]
  wire  _T_1563; // @[Parameters.scala 671:42]
  wire  _T_1564; // @[Parameters.scala 671:42]
  wire  _T_1565; // @[Parameters.scala 671:42]
  wire  _T_1566; // @[Parameters.scala 671:42]
  wire  _T_1567; // @[Parameters.scala 671:42]
  wire  _T_1570; // @[Parameters.scala 92:42]
  wire  _T_1578; // @[Parameters.scala 670:56]
  wire  _T_1581; // @[Monitor.scala 260:78]
  wire  _T_1583; // @[Monitor.scala 42:11]
  wire  _T_1587; // @[Parameters.scala 91:48]
  wire  _T_1588; // @[Mux.scala 27:72]
  wire  _T_1635; // @[Parameters.scala 671:42]
  wire  _T_1636; // @[Parameters.scala 670:56]
  wire  _T_1638; // @[Monitor.scala 261:78]
  wire  _T_1640; // @[Monitor.scala 42:11]
  wire  _T_1660; // @[Monitor.scala 269:25]
  wire  _T_1793; // @[Monitor.scala 278:25]
  wire  _T_1803; // @[Monitor.scala 282:31]
  wire  _T_1805; // @[Monitor.scala 42:11]
  wire  _T_1811; // @[Monitor.scala 286:25]
  wire  _T_1825; // @[Monitor.scala 293:25]
  wire  _a_first_T; // @[Decoupled.scala 40:37]
  wire [8:0] a_first_beats1_decode; // @[Edges.scala 219:59]
  wire  a_first_beats1_opdata; // @[Edges.scala 91:28]
  reg [8:0] a_first_counter; // @[Edges.scala 228:27]
  reg [31:0] _RAND_0;
  wire [8:0] a_first_counter1; // @[Edges.scala 229:28]
  wire  a_first; // @[Edges.scala 230:25]
  reg [2:0] opcode; // @[Monitor.scala 384:22]
  reg [31:0] _RAND_1;
  reg [2:0] param; // @[Monitor.scala 385:22]
  reg [31:0] _RAND_2;
  reg [3:0] size; // @[Monitor.scala 386:22]
  reg [31:0] _RAND_3;
  reg  source; // @[Monitor.scala 387:22]
  reg [31:0] _RAND_4;
  reg [31:0] address; // @[Monitor.scala 388:22]
  reg [31:0] _RAND_5;
  wire  _T_1847; // @[Monitor.scala 389:19]
  wire  _T_1848; // @[Monitor.scala 390:32]
  wire  _T_1850; // @[Monitor.scala 42:11]
  wire  _T_1852; // @[Monitor.scala 391:32]
  wire  _T_1854; // @[Monitor.scala 42:11]
  wire  _T_1856; // @[Monitor.scala 392:32]
  wire  _T_1858; // @[Monitor.scala 42:11]
  wire  _T_1860; // @[Monitor.scala 393:32]
  wire  _T_1862; // @[Monitor.scala 42:11]
  wire  _T_1864; // @[Monitor.scala 394:32]
  wire  _T_1866; // @[Monitor.scala 42:11]
  wire  _T_1869; // @[Monitor.scala 396:20]
  wire  _d_first_T; // @[Decoupled.scala 40:37]
  wire [26:0] _d_first_beats1_decode_T_1; // @[package.scala 234:77]
  wire [8:0] d_first_beats1_decode; // @[Edges.scala 219:59]
  wire  d_first_beats1_opdata; // @[Edges.scala 105:36]
  reg [8:0] d_first_counter; // @[Edges.scala 228:27]
  reg [31:0] _RAND_6;
  wire [8:0] d_first_counter1; // @[Edges.scala 229:28]
  wire  d_first; // @[Edges.scala 230:25]
  reg [2:0] opcode_1; // @[Monitor.scala 535:22]
  reg [31:0] _RAND_7;
  reg [1:0] param_1; // @[Monitor.scala 536:22]
  reg [31:0] _RAND_8;
  reg [3:0] size_1; // @[Monitor.scala 537:22]
  reg [31:0] _RAND_9;
  reg  source_1; // @[Monitor.scala 538:22]
  reg [31:0] _RAND_10;
  reg [1:0] sink; // @[Monitor.scala 539:22]
  reg [31:0] _RAND_11;
  reg  denied; // @[Monitor.scala 540:22]
  reg [31:0] _RAND_12;
  wire  _T_1871; // @[Monitor.scala 541:19]
  wire  _T_1872; // @[Monitor.scala 542:29]
  wire  _T_1874; // @[Monitor.scala 49:11]
  wire  _T_1876; // @[Monitor.scala 543:29]
  wire  _T_1878; // @[Monitor.scala 49:11]
  wire  _T_1880; // @[Monitor.scala 544:29]
  wire  _T_1882; // @[Monitor.scala 49:11]
  wire  _T_1884; // @[Monitor.scala 545:29]
  wire  _T_1886; // @[Monitor.scala 49:11]
  wire  _T_1888; // @[Monitor.scala 546:29]
  wire  _T_1890; // @[Monitor.scala 49:11]
  wire  _T_1892; // @[Monitor.scala 547:29]
  wire  _T_1894; // @[Monitor.scala 49:11]
  wire  _T_1897; // @[Monitor.scala 549:20]
  wire  b_first_done; // @[Decoupled.scala 40:37]
  reg [8:0] b_first_counter; // @[Edges.scala 228:27]
  reg [31:0] _RAND_13;
  wire [8:0] b_first_counter1; // @[Edges.scala 229:28]
  wire  b_first; // @[Edges.scala 230:25]
  reg [2:0] opcode_2; // @[Monitor.scala 407:22]
  reg [31:0] _RAND_14;
  reg [1:0] param_2; // @[Monitor.scala 408:22]
  reg [31:0] _RAND_15;
  reg [3:0] size_2; // @[Monitor.scala 409:22]
  reg [31:0] _RAND_16;
  reg  source_2; // @[Monitor.scala 410:22]
  reg [31:0] _RAND_17;
  reg [31:0] address_1; // @[Monitor.scala 411:22]
  reg [31:0] _RAND_18;
  wire  _T_1899; // @[Monitor.scala 412:19]
  wire  _T_1900; // @[Monitor.scala 413:32]
  wire  _T_1902; // @[Monitor.scala 42:11]
  wire  _T_1904; // @[Monitor.scala 414:32]
  wire  _T_1906; // @[Monitor.scala 42:11]
  wire  _T_1908; // @[Monitor.scala 415:32]
  wire  _T_1910; // @[Monitor.scala 42:11]
  wire  _T_1912; // @[Monitor.scala 416:32]
  wire  _T_1914; // @[Monitor.scala 42:11]
  wire  _T_1916; // @[Monitor.scala 417:32]
  wire  _T_1918; // @[Monitor.scala 42:11]
  wire  _T_1921; // @[Monitor.scala 419:20]
  wire  _c_first_T; // @[Decoupled.scala 40:37]
  wire [8:0] c_first_beats1_decode; // @[Edges.scala 219:59]
  wire  c_first_beats1_opdata; // @[Edges.scala 101:36]
  reg [8:0] c_first_counter; // @[Edges.scala 228:27]
  reg [31:0] _RAND_19;
  wire [8:0] c_first_counter1; // @[Edges.scala 229:28]
  wire  c_first; // @[Edges.scala 230:25]
  reg [2:0] opcode_3; // @[Monitor.scala 512:22]
  reg [31:0] _RAND_20;
  reg [2:0] param_3; // @[Monitor.scala 513:22]
  reg [31:0] _RAND_21;
  reg [3:0] size_3; // @[Monitor.scala 514:22]
  reg [31:0] _RAND_22;
  reg  source_3; // @[Monitor.scala 515:22]
  reg [31:0] _RAND_23;
  reg [31:0] address_2; // @[Monitor.scala 516:22]
  reg [31:0] _RAND_24;
  wire  _T_1923; // @[Monitor.scala 517:19]
  wire  _T_1924; // @[Monitor.scala 518:32]
  wire  _T_1926; // @[Monitor.scala 42:11]
  wire  _T_1928; // @[Monitor.scala 519:32]
  wire  _T_1930; // @[Monitor.scala 42:11]
  wire  _T_1932; // @[Monitor.scala 520:32]
  wire  _T_1934; // @[Monitor.scala 42:11]
  wire  _T_1936; // @[Monitor.scala 521:32]
  wire  _T_1938; // @[Monitor.scala 42:11]
  wire  _T_1940; // @[Monitor.scala 522:32]
  wire  _T_1942; // @[Monitor.scala 42:11]
  wire  _T_1945; // @[Monitor.scala 524:20]
  reg [1:0] inflight; // @[Monitor.scala 611:27]
  reg [31:0] _RAND_25;
  reg [7:0] inflight_opcodes; // @[Monitor.scala 613:35]
  reg [31:0] _RAND_26;
  reg [15:0] inflight_sizes; // @[Monitor.scala 615:33]
  reg [31:0] _RAND_27;
  reg [8:0] a_first_counter_1; // @[Edges.scala 228:27]
  reg [31:0] _RAND_28;
  wire [8:0] a_first_counter1_1; // @[Edges.scala 229:28]
  wire  a_first_1; // @[Edges.scala 230:25]
  reg [8:0] d_first_counter_1; // @[Edges.scala 228:27]
  reg [31:0] _RAND_29;
  wire [8:0] d_first_counter1_1; // @[Edges.scala 229:28]
  wire  d_first_1; // @[Edges.scala 230:25]
  wire [2:0] _GEN_89; // @[Monitor.scala 634:69]
  wire [3:0] _a_opcode_lookup_T; // @[Monitor.scala 634:69]
  wire [7:0] _a_opcode_lookup_T_1; // @[Monitor.scala 634:44]
  wire [15:0] _a_opcode_lookup_T_5; // @[Monitor.scala 609:57]
  wire [15:0] _GEN_90; // @[Monitor.scala 634:97]
  wire [15:0] _a_opcode_lookup_T_6; // @[Monitor.scala 634:97]
  wire [15:0] _a_opcode_lookup_T_7; // @[Monitor.scala 634:152]
  wire [3:0] _a_size_lookup_T; // @[Monitor.scala 638:65]
  wire [15:0] _a_size_lookup_T_1; // @[Monitor.scala 638:40]
  wire [15:0] _a_size_lookup_T_5; // @[Monitor.scala 609:57]
  wire [15:0] _a_size_lookup_T_6; // @[Monitor.scala 638:91]
  wire [15:0] _a_size_lookup_T_7; // @[Monitor.scala 638:144]
  wire  _T_1946; // @[Monitor.scala 648:26]
  wire [1:0] _a_set_wo_ready_T; // @[OneHot.scala 58:35]
  wire [1:0] a_set_wo_ready; // @[Monitor.scala 648:71]
  wire  _T_1949; // @[Monitor.scala 652:27]
  wire [3:0] _a_opcodes_set_interm_T; // @[Monitor.scala 654:53]
  wire [3:0] _a_opcodes_set_interm_T_1; // @[Monitor.scala 654:61]
  wire [4:0] _a_sizes_set_interm_T; // @[Monitor.scala 655:51]
  wire [4:0] _a_sizes_set_interm_T_1; // @[Monitor.scala 655:59]
  wire [2:0] _GEN_93; // @[Monitor.scala 656:79]
  wire [3:0] _a_opcodes_set_T; // @[Monitor.scala 656:79]
  wire [3:0] a_opcodes_set_interm; // @[Monitor.scala 652:72]
  wire [18:0] _GEN_94; // @[Monitor.scala 656:54]
  wire [18:0] _a_opcodes_set_T_1; // @[Monitor.scala 656:54]
  wire [3:0] _a_sizes_set_T; // @[Monitor.scala 657:77]
  wire [4:0] a_sizes_set_interm; // @[Monitor.scala 652:72]
  wire [19:0] _GEN_95; // @[Monitor.scala 657:52]
  wire [19:0] _a_sizes_set_T_1; // @[Monitor.scala 657:52]
  wire [1:0] _T_1951; // @[Monitor.scala 658:26]
  wire  _T_1955; // @[Monitor.scala 42:11]
  wire [1:0] a_set; // @[Monitor.scala 652:72]
  wire [18:0] _GEN_31; // @[Monitor.scala 652:72]
  wire [19:0] _GEN_32; // @[Monitor.scala 652:72]
  wire  _T_1957; // @[Monitor.scala 671:26]
  wire  _T_1960; // @[Monitor.scala 671:71]
  wire [1:0] _d_clr_wo_ready_T; // @[OneHot.scala 58:35]
  wire [1:0] d_clr_wo_ready; // @[Monitor.scala 671:90]
  wire  _T_1962; // @[Monitor.scala 675:27]
  wire  _T_1965; // @[Monitor.scala 675:72]
  wire [30:0] _GEN_97; // @[Monitor.scala 677:76]
  wire [30:0] _d_opcodes_clr_T_5; // @[Monitor.scala 677:76]
  wire [30:0] _GEN_98; // @[Monitor.scala 678:74]
  wire [30:0] _d_sizes_clr_T_5; // @[Monitor.scala 678:74]
  wire [1:0] d_clr; // @[Monitor.scala 675:91]
  wire [30:0] _GEN_35; // @[Monitor.scala 675:91]
  wire [30:0] _GEN_36; // @[Monitor.scala 675:91]
  wire  _same_cycle_resp_T_2; // @[Monitor.scala 681:113]
  wire  same_cycle_resp; // @[Monitor.scala 681:88]
  wire [1:0] _T_1970; // @[Monitor.scala 682:25]
  wire  _T_1972; // @[Monitor.scala 682:49]
  wire  _T_1974; // @[Monitor.scala 49:11]
  wire [2:0] _GEN_39; // @[Monitor.scala 685:38]
  wire [2:0] _GEN_40; // @[Monitor.scala 685:38]
  wire [2:0] _GEN_41; // @[Monitor.scala 685:38]
  wire [2:0] _GEN_42; // @[Monitor.scala 685:38]
  wire [2:0] _GEN_43; // @[Monitor.scala 685:38]
  wire [2:0] _GEN_44; // @[Monitor.scala 685:38]
  wire  _T_1976; // @[Monitor.scala 685:38]
  wire [2:0] _GEN_51; // @[Monitor.scala 686:39]
  wire [2:0] _GEN_52; // @[Monitor.scala 686:39]
  wire  _T_1977; // @[Monitor.scala 686:39]
  wire  _T_1978; // @[Monitor.scala 685:77]
  wire  _T_1980; // @[Monitor.scala 49:11]
  wire  _T_1982; // @[Monitor.scala 687:36]
  wire  _T_1984; // @[Monitor.scala 49:11]
  wire [3:0] a_opcode_lookup; // @[Monitor.scala 634:21]
  wire [2:0] _GEN_55; // @[Monitor.scala 689:38]
  wire [2:0] _GEN_56; // @[Monitor.scala 689:38]
  wire [2:0] _GEN_57; // @[Monitor.scala 689:38]
  wire [2:0] _GEN_58; // @[Monitor.scala 689:38]
  wire [2:0] _GEN_59; // @[Monitor.scala 689:38]
  wire [2:0] _GEN_60; // @[Monitor.scala 689:38]
  wire  _T_1987; // @[Monitor.scala 689:38]
  wire [2:0] _GEN_67; // @[Monitor.scala 690:38]
  wire [2:0] _GEN_68; // @[Monitor.scala 690:38]
  wire  _T_1989; // @[Monitor.scala 690:38]
  wire  _T_1990; // @[Monitor.scala 689:72]
  wire  _T_1992; // @[Monitor.scala 49:11]
  wire [7:0] a_size_lookup; // @[Monitor.scala 638:19]
  wire [7:0] _GEN_99; // @[Monitor.scala 691:36]
  wire  _T_1994; // @[Monitor.scala 691:36]
  wire  _T_1996; // @[Monitor.scala 49:11]
  wire  _T_1999; // @[Monitor.scala 694:36]
  wire  _T_2000; // @[Monitor.scala 694:47]
  wire  _T_2002; // @[Monitor.scala 694:65]
  wire  _T_2004; // @[Monitor.scala 694:116]
  wire  _T_2006; // @[Monitor.scala 695:32]
  wire  _T_2008; // @[Monitor.scala 49:11]
  wire  _T_2010; // @[Monitor.scala 699:29]
  wire  _T_2011; // @[Monitor.scala 699:67]
  wire  _T_2013; // @[Monitor.scala 699:48]
  wire  _T_2015; // @[Monitor.scala 49:11]
  wire [1:0] _inflight_T; // @[Monitor.scala 702:27]
  wire [1:0] _inflight_T_2; // @[Monitor.scala 702:36]
  wire [7:0] a_opcodes_set; // @[Monitor.scala 656:28]
  wire [7:0] _inflight_opcodes_T; // @[Monitor.scala 703:43]
  wire [7:0] d_opcodes_clr; // @[Monitor.scala 677:21]
  wire [7:0] _inflight_opcodes_T_2; // @[Monitor.scala 703:60]
  wire [15:0] a_sizes_set; // @[Monitor.scala 657:28]
  wire [15:0] _inflight_sizes_T; // @[Monitor.scala 704:39]
  wire [15:0] d_sizes_clr; // @[Monitor.scala 678:21]
  wire [15:0] _inflight_sizes_T_2; // @[Monitor.scala 704:54]
  reg [31:0] watchdog; // @[Monitor.scala 706:27]
  reg [31:0] _RAND_30;
  wire  _T_2017; // @[Monitor.scala 709:26]
  wire  _T_2019; // @[Monitor.scala 709:39]
  wire  _T_2020; // @[Monitor.scala 709:30]
  wire  _T_2021; // @[Monitor.scala 709:59]
  wire  _T_2022; // @[Monitor.scala 709:47]
  wire  _T_2024; // @[Monitor.scala 42:11]
  wire [31:0] _watchdog_T_1; // @[Monitor.scala 711:26]
  wire  _T_2028; // @[Monitor.scala 712:27]
  reg [1:0] inflight_1; // @[Monitor.scala 723:35]
  reg [31:0] _RAND_31;
  reg [15:0] inflight_sizes_1; // @[Monitor.scala 725:35]
  reg [31:0] _RAND_32;
  reg [8:0] c_first_counter_1; // @[Edges.scala 228:27]
  reg [31:0] _RAND_33;
  wire [8:0] c_first_counter1_1; // @[Edges.scala 229:28]
  wire  c_first_1; // @[Edges.scala 230:25]
  reg [8:0] d_first_counter_2; // @[Edges.scala 228:27]
  reg [31:0] _RAND_34;
  wire [8:0] d_first_counter1_2; // @[Edges.scala 229:28]
  wire  d_first_2; // @[Edges.scala 230:25]
  wire [15:0] _c_size_lookup_T_1; // @[Monitor.scala 747:42]
  wire [15:0] _c_size_lookup_T_6; // @[Monitor.scala 747:93]
  wire [15:0] _c_size_lookup_T_7; // @[Monitor.scala 747:146]
  wire  _T_2029; // @[Monitor.scala 756:26]
  wire  _T_2032; // @[Edges.scala 67:40]
  wire  _T_2033; // @[Monitor.scala 756:37]
  wire [1:0] _c_set_wo_ready_T; // @[OneHot.scala 58:35]
  wire [1:0] c_set_wo_ready; // @[Monitor.scala 756:71]
  wire  _T_2035; // @[Monitor.scala 760:27]
  wire  _T_2039; // @[Monitor.scala 760:38]
  wire [4:0] _c_sizes_set_interm_T; // @[Monitor.scala 763:51]
  wire [4:0] _c_sizes_set_interm_T_1; // @[Monitor.scala 763:59]
  wire [3:0] _c_sizes_set_T; // @[Monitor.scala 765:77]
  wire [4:0] c_sizes_set_interm; // @[Monitor.scala 760:72]
  wire [19:0] _GEN_106; // @[Monitor.scala 765:52]
  wire [19:0] _c_sizes_set_T_1; // @[Monitor.scala 765:52]
  wire [1:0] _T_2040; // @[Monitor.scala 766:26]
  wire  _T_2044; // @[Monitor.scala 42:11]
  wire [1:0] c_set; // @[Monitor.scala 760:72]
  wire [19:0] _GEN_77; // @[Monitor.scala 760:72]
  wire  _T_2046; // @[Monitor.scala 779:26]
  wire  _T_2048; // @[Monitor.scala 779:71]
  wire [1:0] d_clr_wo_ready_1; // @[Monitor.scala 779:89]
  wire  _T_2050; // @[Monitor.scala 783:27]
  wire  _T_2052; // @[Monitor.scala 783:72]
  wire [1:0] d_clr_1; // @[Monitor.scala 783:90]
  wire [30:0] _GEN_81; // @[Monitor.scala 783:90]
  wire  _same_cycle_resp_T_8; // @[Monitor.scala 790:113]
  wire  same_cycle_resp_1; // @[Monitor.scala 790:88]
  wire [1:0] _T_2056; // @[Monitor.scala 791:25]
  wire  _T_2058; // @[Monitor.scala 791:49]
  wire  _T_2060; // @[Monitor.scala 49:11]
  wire  _T_2062; // @[Monitor.scala 793:36]
  wire  _T_2064; // @[Monitor.scala 49:11]
  wire [7:0] c_size_lookup; // @[Monitor.scala 747:21]
  wire  _T_2066; // @[Monitor.scala 795:36]
  wire  _T_2068; // @[Monitor.scala 49:11]
  wire  _T_2071; // @[Monitor.scala 799:36]
  wire  _T_2072; // @[Monitor.scala 799:47]
  wire  _T_2074; // @[Monitor.scala 799:65]
  wire  _T_2075; // @[Monitor.scala 799:116]
  wire  _T_2077; // @[Monitor.scala 800:32]
  wire  _T_2079; // @[Monitor.scala 49:11]
  wire  _T_2081; // @[Monitor.scala 804:28]
  wire  _T_2082; // @[Monitor.scala 805:31]
  wire  _T_2084; // @[Monitor.scala 49:11]
  wire [1:0] _inflight_T_3; // @[Monitor.scala 809:35]
  wire [1:0] _inflight_T_5; // @[Monitor.scala 809:44]
  wire [15:0] c_sizes_set; // @[Monitor.scala 765:28]
  wire [15:0] _inflight_sizes_T_3; // @[Monitor.scala 811:41]
  wire [15:0] d_sizes_clr_1; // @[Monitor.scala 786:21]
  wire [15:0] _inflight_sizes_T_5; // @[Monitor.scala 811:56]
  reg [31:0] watchdog_1; // @[Monitor.scala 813:27]
  reg [31:0] _RAND_35;
  wire  _T_2086; // @[Monitor.scala 816:26]
  wire  _T_2088; // @[Monitor.scala 816:39]
  wire  _T_2089; // @[Monitor.scala 816:30]
  wire  _T_2090; // @[Monitor.scala 816:59]
  wire  _T_2091; // @[Monitor.scala 816:47]
  wire  _T_2093; // @[Monitor.scala 42:11]
  wire [31:0] _watchdog_T_3; // @[Monitor.scala 818:26]
  wire  _T_2097; // @[Monitor.scala 819:27]
  reg [3:0] inflight_2; // @[Monitor.scala 823:27]
  reg [31:0] _RAND_36;
  reg [8:0] d_first_counter_3; // @[Edges.scala 228:27]
  reg [31:0] _RAND_37;
  wire [8:0] d_first_counter1_3; // @[Edges.scala 229:28]
  wire  d_first_3; // @[Edges.scala 230:25]
  wire  _T_2099; // @[Monitor.scala 829:27]
  wire  _T_2103; // @[Edges.scala 70:40]
  wire  _T_2104; // @[Monitor.scala 829:38]
  wire [3:0] _d_set_T; // @[OneHot.scala 58:35]
  wire [3:0] _T_2105; // @[Monitor.scala 831:23]
  wire  _T_2109; // @[Monitor.scala 49:11]
  wire [3:0] d_set; // @[Monitor.scala 829:72]
  wire  _T_2111; // @[Decoupled.scala 40:37]
  wire [3:0] _e_clr_T; // @[OneHot.scala 58:35]
  wire [3:0] _T_2114; // @[Monitor.scala 837:24]
  wire [3:0] _T_2115; // @[Monitor.scala 837:35]
  wire  _T_2118; // @[Monitor.scala 42:11]
  wire [3:0] e_clr; // @[Monitor.scala 835:73]
  wire [3:0] _inflight_T_6; // @[Monitor.scala 842:27]
  wire [3:0] _inflight_T_8; // @[Monitor.scala 842:36]
  wire  _GEN_111; // @[Monitor.scala 42:11]
  wire  _GEN_125; // @[Monitor.scala 42:11]
  wire  _GEN_141; // @[Monitor.scala 42:11]
  wire  _GEN_153; // @[Monitor.scala 42:11]
  wire  _GEN_163; // @[Monitor.scala 42:11]
  wire  _GEN_173; // @[Monitor.scala 42:11]
  wire  _GEN_183; // @[Monitor.scala 42:11]
  wire  _GEN_193; // @[Monitor.scala 42:11]
  wire  _GEN_203; // @[Monitor.scala 49:11]
  wire  _GEN_213; // @[Monitor.scala 49:11]
  wire  _GEN_223; // @[Monitor.scala 49:11]
  wire  _GEN_233; // @[Monitor.scala 49:11]
  wire  _GEN_239; // @[Monitor.scala 49:11]
  wire  _GEN_245; // @[Monitor.scala 49:11]
  wire  _GEN_251; // @[Monitor.scala 49:11]
  wire  _GEN_265; // @[Monitor.scala 42:11]
  wire  _GEN_279; // @[Monitor.scala 42:11]
  wire  _GEN_291; // @[Monitor.scala 42:11]
  wire  _GEN_303; // @[Monitor.scala 42:11]
  wire  _GEN_313; // @[Monitor.scala 42:11]
  wire  _GEN_323; // @[Monitor.scala 42:11]
  wire  _GEN_335; // @[Monitor.scala 42:11]
  wire  _GEN_345; // @[Monitor.scala 42:11]
  wire  _GEN_355; // @[Monitor.scala 42:11]
  wire  _GEN_367; // @[Monitor.scala 42:11]
  wire  _GEN_379; // @[Monitor.scala 42:11]
  wire  _GEN_387; // @[Monitor.scala 42:11]
  wire  _GEN_395; // @[Monitor.scala 42:11]
  wire  _GEN_403; // @[Monitor.scala 49:11]
  wire  _GEN_408; // @[Monitor.scala 49:11]
  wire  _GEN_415; // @[Monitor.scala 49:11]
  wire  _GEN_418; // @[Monitor.scala 49:11]
  wire [29:0] TLMonitor_23_covSum;
  wire  stopEn0;
  wire  stopEn1;
  wire  stopEn2;
  wire  stopEn3;
  wire  stopEn4;
  wire  stopEn5;
  wire  stopEn6;
  wire  stopEn7;
  wire  stopEn8;
  wire  stopEn9;
  wire  stopEn10;
  wire  stopEn11;
  wire  stopEn12;
  wire  stopEn13;
  wire  stopEn14;
  wire  stopEn15;
  wire  stopEn16;
  wire  stopEn17;
  wire  stopEn18;
  wire  stopEn19;
  wire  stopEn20;
  wire  stopEn21;
  wire  stopEn22;
  wire  stopEn23;
  wire  stopEn24;
  wire  stopEn25;
  wire  stopEn26;
  wire  stopEn27;
  wire  stopEn28;
  wire  stopEn29;
  wire  stopEn30;
  wire  stopEn31;
  wire  stopEn32;
  wire  stopEn33;
  wire  stopEn34;
  wire  stopEn35;
  wire  stopEn36;
  wire  stopEn37;
  wire  stopEn38;
  wire  stopEn39;
  wire  stopEn40;
  wire  stopEn41;
  wire  stopEn42;
  wire  stopEn43;
  wire  stopEn44;
  wire  stopEn45;
  wire  stopEn46;
  wire  stopEn47;
  wire  stopEn48;
  wire  stopEn49;
  wire  stopEn50;
  wire  stopEn51;
  wire  stopEn52;
  wire  stopEn53;
  wire  stopEn54;
  wire  stopEn55;
  wire  stopEn56;
  wire  stopEn57;
  wire  stopEn58;
  wire  stopEn59;
  wire  stopEn60;
  wire  stopEn61;
  wire  stopEn62;
  wire  stopEn63;
  wire  stopEn64;
  wire  stopEn65;
  wire  stopEn66;
  wire  stopEn67;
  wire  stopEn68;
  wire  stopEn69;
  wire  stopEn70;
  wire  stopEn71;
  wire  stopEn72;
  wire  stopEn73;
  wire  stopEn74;
  wire  stopEn75;
  wire  stopEn76;
  wire  stopEn77;
  wire  stopEn78;
  wire  stopEn79;
  wire  stopEn80;
  wire  stopEn81;
  wire  stopEn82;
  wire  stopEn83;
  wire  stopEn84;
  wire  stopEn85;
  wire  stopEn86;
  wire  stopEn87;
  wire  stopEn88;
  wire  stopEn89;
  wire  stopEn90;
  wire  stopEn91;
  wire  stopEn92;
  wire  stopEn93;
  wire  stopEn94;
  wire  stopEn95;
  wire  stopEn96;
  wire  stopEn97;
  wire  stopEn98;
  wire  stopEn99;
  wire  stopEn100;
  wire  stopEn101;
  wire  stopEn102;
  wire  stopEn103;
  wire  stopEn104;
  wire  stopEn105;
  wire  stopEn106;
  wire  stopEn107;
  wire  stopEn108;
  wire  stopEn109;
  wire  stopEn110;
  wire  stopEn111;
  wire  stopEn112;
  wire  stopEn113;
  wire  stopEn114;
  wire  stopEn115;
  wire  stopEn116;
  wire  stopEn117;
  wire  stopEn118;
  wire  stopEn119;
  wire  stopEn120;
  wire  stopEn121;
  wire  stopEn122;
  wire  stopEn123;
  wire  stopEn124;
  wire  stopEn125;
  wire  stopEn126;
  wire  stopEn127;
  wire  stopEn128;
  wire  stopEn129;
  wire  stopEn130;
  wire  stopEn131;
  wire  stopEn132;
  wire  stopEn133;
  wire  stopEn134;
  wire  stopEn135;
  wire  stopEn136;
  wire  stopEn137;
  wire  stopEn138;
  wire  stopEn139;
  wire  stopEn140;
  wire  stopEn141;
  wire  stopEn142;
  wire  stopEn143;
  wire  stopEn144;
  wire  stopEn145;
  wire  stopEn146;
  wire  stopEn147;
  wire  stopEn148;
  wire  stopEn149;
  wire  stopEn150;
  wire  stopEn151;
  wire  stopEn152;
  wire  stopEn153;
  wire  stopEn154;
  wire  stopEn155;
  wire  stopEn156;
  wire  stopEn157;
  wire  stopEn158;
  wire  stopEn159;
  wire  stopEn160;
  wire  stopEn161;
  wire  stopEn162;
  wire  stopEn163;
  wire  stopEn164;
  wire  stopEn165;
  wire  stopEn166;
  wire  stopEn167;
  wire  stopEn168;
  wire  stopEn169;
  wire  stopEn170;
  wire  stopEn171;
  wire  stopEn172;
  wire  stopEn173;
  wire  stopEn174;
  wire  stopEn175;
  wire  stopEn176;
  wire  stopEn177;
  wire  stopEn178;
  wire  stopEn179;
  wire  stopEn180;
  wire  stopEn181;
  wire  stopEn182;
  wire  stopEn183;
  wire  stopEn184;
  wire  stopEn185;
  wire  stopEn186;
  wire  plusarg_reader_metaAssert_wire;
  wire  plusarg_reader_1_metaAssert_wire;
  wire  TLMonitor_23_or63;
  wire  TLMonitor_23_or130;
  wire  TLMonitor_23_or64;
  wire  TLMonitor_23_or31;
  wire  TLMonitor_23_or132;
  wire  TLMonitor_23_or65;
  wire  TLMonitor_23_or134;
  wire  TLMonitor_23_or66;
  wire  TLMonitor_23_or32;
  wire  TLMonitor_23_or15;
  wire  TLMonitor_23_or136;
  wire  TLMonitor_23_or67;
  wire  TLMonitor_23_or138;
  wire  TLMonitor_23_or68;
  wire  TLMonitor_23_or33;
  wire  TLMonitor_23_or140;
  wire  TLMonitor_23_or69;
  wire  TLMonitor_23_or142;
  wire  TLMonitor_23_or70;
  wire  TLMonitor_23_or34;
  wire  TLMonitor_23_or16;
  wire  TLMonitor_23_or7;
  wire  TLMonitor_23_or144;
  wire  TLMonitor_23_or71;
  wire  TLMonitor_23_or146;
  wire  TLMonitor_23_or72;
  wire  TLMonitor_23_or35;
  wire  TLMonitor_23_or148;
  wire  TLMonitor_23_or73;
  wire  TLMonitor_23_or150;
  wire  TLMonitor_23_or74;
  wire  TLMonitor_23_or36;
  wire  TLMonitor_23_or17;
  wire  TLMonitor_23_or152;
  wire  TLMonitor_23_or75;
  wire  TLMonitor_23_or154;
  wire  TLMonitor_23_or76;
  wire  TLMonitor_23_or37;
  wire  TLMonitor_23_or156;
  wire  TLMonitor_23_or77;
  wire  TLMonitor_23_or158;
  wire  TLMonitor_23_or78;
  wire  TLMonitor_23_or38;
  wire  TLMonitor_23_or18;
  wire  TLMonitor_23_or8;
  wire  TLMonitor_23_or3;
  wire  TLMonitor_23_or79;
  wire  TLMonitor_23_or162;
  wire  TLMonitor_23_or80;
  wire  TLMonitor_23_or39;
  wire  TLMonitor_23_or164;
  wire  TLMonitor_23_or81;
  wire  TLMonitor_23_or166;
  wire  TLMonitor_23_or82;
  wire  TLMonitor_23_or40;
  wire  TLMonitor_23_or19;
  wire  TLMonitor_23_or168;
  wire  TLMonitor_23_or83;
  wire  TLMonitor_23_or170;
  wire  TLMonitor_23_or84;
  wire  TLMonitor_23_or41;
  wire  TLMonitor_23_or172;
  wire  TLMonitor_23_or85;
  wire  TLMonitor_23_or174;
  wire  TLMonitor_23_or86;
  wire  TLMonitor_23_or42;
  wire  TLMonitor_23_or20;
  wire  TLMonitor_23_or9;
  wire  TLMonitor_23_or176;
  wire  TLMonitor_23_or87;
  wire  TLMonitor_23_or178;
  wire  TLMonitor_23_or88;
  wire  TLMonitor_23_or43;
  wire  TLMonitor_23_or180;
  wire  TLMonitor_23_or89;
  wire  TLMonitor_23_or182;
  wire  TLMonitor_23_or90;
  wire  TLMonitor_23_or44;
  wire  TLMonitor_23_or21;
  wire  TLMonitor_23_or184;
  wire  TLMonitor_23_or91;
  wire  TLMonitor_23_or186;
  wire  TLMonitor_23_or92;
  wire  TLMonitor_23_or45;
  wire  TLMonitor_23_or188;
  wire  TLMonitor_23_or93;
  wire  TLMonitor_23_or190;
  wire  TLMonitor_23_or94;
  wire  TLMonitor_23_or46;
  wire  TLMonitor_23_or22;
  wire  TLMonitor_23_or10;
  wire  TLMonitor_23_or4;
  wire  TLMonitor_23_or1;
  wire  TLMonitor_23_or95;
  wire  TLMonitor_23_or194;
  wire  TLMonitor_23_or96;
  wire  TLMonitor_23_or47;
  wire  TLMonitor_23_or196;
  wire  TLMonitor_23_or97;
  wire  TLMonitor_23_or198;
  wire  TLMonitor_23_or98;
  wire  TLMonitor_23_or48;
  wire  TLMonitor_23_or23;
  wire  TLMonitor_23_or200;
  wire  TLMonitor_23_or99;
  wire  TLMonitor_23_or202;
  wire  TLMonitor_23_or100;
  wire  TLMonitor_23_or49;
  wire  TLMonitor_23_or204;
  wire  TLMonitor_23_or101;
  wire  TLMonitor_23_or206;
  wire  TLMonitor_23_or102;
  wire  TLMonitor_23_or50;
  wire  TLMonitor_23_or24;
  wire  TLMonitor_23_or11;
  wire  TLMonitor_23_or208;
  wire  TLMonitor_23_or103;
  wire  TLMonitor_23_or210;
  wire  TLMonitor_23_or104;
  wire  TLMonitor_23_or51;
  wire  TLMonitor_23_or212;
  wire  TLMonitor_23_or105;
  wire  TLMonitor_23_or214;
  wire  TLMonitor_23_or106;
  wire  TLMonitor_23_or52;
  wire  TLMonitor_23_or25;
  wire  TLMonitor_23_or216;
  wire  TLMonitor_23_or107;
  wire  TLMonitor_23_or218;
  wire  TLMonitor_23_or108;
  wire  TLMonitor_23_or53;
  wire  TLMonitor_23_or220;
  wire  TLMonitor_23_or109;
  wire  TLMonitor_23_or222;
  wire  TLMonitor_23_or110;
  wire  TLMonitor_23_or54;
  wire  TLMonitor_23_or26;
  wire  TLMonitor_23_or12;
  wire  TLMonitor_23_or5;
  wire  TLMonitor_23_or224;
  wire  TLMonitor_23_or111;
  wire  TLMonitor_23_or226;
  wire  TLMonitor_23_or112;
  wire  TLMonitor_23_or55;
  wire  TLMonitor_23_or228;
  wire  TLMonitor_23_or113;
  wire  TLMonitor_23_or230;
  wire  TLMonitor_23_or114;
  wire  TLMonitor_23_or56;
  wire  TLMonitor_23_or27;
  wire  TLMonitor_23_or232;
  wire  TLMonitor_23_or115;
  wire  TLMonitor_23_or234;
  wire  TLMonitor_23_or116;
  wire  TLMonitor_23_or57;
  wire  TLMonitor_23_or236;
  wire  TLMonitor_23_or117;
  wire  TLMonitor_23_or238;
  wire  TLMonitor_23_or118;
  wire  TLMonitor_23_or58;
  wire  TLMonitor_23_or28;
  wire  TLMonitor_23_or13;
  wire  TLMonitor_23_or240;
  wire  TLMonitor_23_or119;
  wire  TLMonitor_23_or242;
  wire  TLMonitor_23_or120;
  wire  TLMonitor_23_or59;
  wire  TLMonitor_23_or244;
  wire  TLMonitor_23_or121;
  wire  TLMonitor_23_or246;
  wire  TLMonitor_23_or122;
  wire  TLMonitor_23_or60;
  wire  TLMonitor_23_or29;
  wire  TLMonitor_23_or248;
  wire  TLMonitor_23_or123;
  wire  TLMonitor_23_or250;
  wire  TLMonitor_23_or124;
  wire  TLMonitor_23_or61;
  wire  TLMonitor_23_or252;
  wire  TLMonitor_23_or125;
  wire  TLMonitor_23_or254;
  wire  TLMonitor_23_or126;
  wire  TLMonitor_23_or62;
  wire  TLMonitor_23_or30;
  wire  TLMonitor_23_or14;
  wire  TLMonitor_23_or6;
  wire  TLMonitor_23_or2;
  wire  TLMonitor_23_or0;
  reg  TLMonitor_23_metaAssert;
  reg [31:0] _RAND_38;
//  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11]
//    .out(plusarg_reader_out)
//  );
//  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 ( // @[PlusArg.scala 80:11]
//    .out(plusarg_reader_1_out)
//  );
  assign source_ok = ~io_in_a_bits_source | io_in_a_bits_source; // @[Parameters.scala 1125:46]
  assign _is_aligned_mask_T_1 = 27'hfff << io_in_a_bits_size; // @[package.scala 234:77]
  assign is_aligned_mask = ~_is_aligned_mask_T_1[11:0]; // @[package.scala 234:46]
  assign _GEN_86 = {{20'd0}, is_aligned_mask}; // @[Edges.scala 20:16]
  assign _is_aligned_T = io_in_a_bits_address & _GEN_86; // @[Edges.scala 20:16]
  assign is_aligned = _is_aligned_T == 32'h0; // @[Edges.scala 20:24]
  assign mask_sizeOH_shiftAmount = io_in_a_bits_size[1:0]; // @[OneHot.scala 64:49]
  assign _mask_sizeOH_T_1 = 4'h1 << mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12]
  assign mask_sizeOH = _mask_sizeOH_T_1[2:0] | 3'h1; // @[Misc.scala 201:81]
  assign _mask_T = io_in_a_bits_size >= 4'h3; // @[Misc.scala 205:21]
  assign mask_size = mask_sizeOH[2]; // @[Misc.scala 208:26]
  assign mask_bit = io_in_a_bits_address[2]; // @[Misc.scala 209:26]
  assign mask_nbit = ~mask_bit; // @[Misc.scala 210:20]
  assign _mask_acc_T = mask_size & mask_nbit; // @[Misc.scala 214:38]
  assign mask_acc = _mask_T | _mask_acc_T; // @[Misc.scala 214:29]
  assign _mask_acc_T_1 = mask_size & mask_bit; // @[Misc.scala 214:38]
  assign mask_acc_1 = _mask_T | _mask_acc_T_1; // @[Misc.scala 214:29]
  assign mask_size_1 = mask_sizeOH[1]; // @[Misc.scala 208:26]
  assign mask_bit_1 = io_in_a_bits_address[1]; // @[Misc.scala 209:26]
  assign mask_nbit_1 = ~mask_bit_1; // @[Misc.scala 210:20]
  assign mask_eq_2 = mask_nbit & mask_nbit_1; // @[Misc.scala 213:27]
  assign _mask_acc_T_2 = mask_size_1 & mask_eq_2; // @[Misc.scala 214:38]
  assign mask_acc_2 = mask_acc | _mask_acc_T_2; // @[Misc.scala 214:29]
  assign mask_eq_3 = mask_nbit & mask_bit_1; // @[Misc.scala 213:27]
  assign _mask_acc_T_3 = mask_size_1 & mask_eq_3; // @[Misc.scala 214:38]
  assign mask_acc_3 = mask_acc | _mask_acc_T_3; // @[Misc.scala 214:29]
  assign mask_eq_4 = mask_bit & mask_nbit_1; // @[Misc.scala 213:27]
  assign _mask_acc_T_4 = mask_size_1 & mask_eq_4; // @[Misc.scala 214:38]
  assign mask_acc_4 = mask_acc_1 | _mask_acc_T_4; // @[Misc.scala 214:29]
  assign mask_eq_5 = mask_bit & mask_bit_1; // @[Misc.scala 213:27]
  assign _mask_acc_T_5 = mask_size_1 & mask_eq_5; // @[Misc.scala 214:38]
  assign mask_acc_5 = mask_acc_1 | _mask_acc_T_5; // @[Misc.scala 214:29]
  assign mask_size_2 = mask_sizeOH[0]; // @[Misc.scala 208:26]
  assign mask_bit_2 = io_in_a_bits_address[0]; // @[Misc.scala 209:26]
  assign mask_nbit_2 = ~mask_bit_2; // @[Misc.scala 210:20]
  assign mask_eq_6 = mask_eq_2 & mask_nbit_2; // @[Misc.scala 213:27]
  assign _mask_acc_T_6 = mask_size_2 & mask_eq_6; // @[Misc.scala 214:38]
  assign mask_lo_lo_lo = mask_acc_2 | _mask_acc_T_6; // @[Misc.scala 214:29]
  assign mask_eq_7 = mask_eq_2 & mask_bit_2; // @[Misc.scala 213:27]
  assign _mask_acc_T_7 = mask_size_2 & mask_eq_7; // @[Misc.scala 214:38]
  assign mask_lo_lo_hi = mask_acc_2 | _mask_acc_T_7; // @[Misc.scala 214:29]
  assign mask_eq_8 = mask_eq_3 & mask_nbit_2; // @[Misc.scala 213:27]
  assign _mask_acc_T_8 = mask_size_2 & mask_eq_8; // @[Misc.scala 214:38]
  assign mask_lo_hi_lo = mask_acc_3 | _mask_acc_T_8; // @[Misc.scala 214:29]
  assign mask_eq_9 = mask_eq_3 & mask_bit_2; // @[Misc.scala 213:27]
  assign _mask_acc_T_9 = mask_size_2 & mask_eq_9; // @[Misc.scala 214:38]
  assign mask_lo_hi_hi = mask_acc_3 | _mask_acc_T_9; // @[Misc.scala 214:29]
  assign mask_eq_10 = mask_eq_4 & mask_nbit_2; // @[Misc.scala 213:27]
  assign _mask_acc_T_10 = mask_size_2 & mask_eq_10; // @[Misc.scala 214:38]
  assign mask_hi_lo_lo = mask_acc_4 | _mask_acc_T_10; // @[Misc.scala 214:29]
  assign mask_eq_11 = mask_eq_4 & mask_bit_2; // @[Misc.scala 213:27]
  assign _mask_acc_T_11 = mask_size_2 & mask_eq_11; // @[Misc.scala 214:38]
  assign mask_hi_lo_hi = mask_acc_4 | _mask_acc_T_11; // @[Misc.scala 214:29]
  assign mask_eq_12 = mask_eq_5 & mask_nbit_2; // @[Misc.scala 213:27]
  assign _mask_acc_T_12 = mask_size_2 & mask_eq_12; // @[Misc.scala 214:38]
  assign mask_hi_hi_lo = mask_acc_5 | _mask_acc_T_12; // @[Misc.scala 214:29]
  assign mask_eq_13 = mask_eq_5 & mask_bit_2; // @[Misc.scala 213:27]
  assign _mask_acc_T_13 = mask_size_2 & mask_eq_13; // @[Misc.scala 214:38]
  assign mask_hi_hi_hi = mask_acc_5 | _mask_acc_T_13; // @[Misc.scala 214:29]
  assign mask = {mask_hi_hi_hi,mask_hi_hi_lo,mask_hi_lo_hi,mask_hi_lo_lo,mask_lo_hi_hi,mask_lo_hi_lo,mask_lo_lo_hi,mask_lo_lo_lo}; // @[Cat.scala 30:58]
  assign _T_7 = {1'b0,$signed(io_in_a_bits_address)}; // @[Parameters.scala 137:49]
  assign _T_24 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 81:25]
  assign _T_26 = io_in_a_bits_size <= 4'hc; // @[Parameters.scala 92:42]
  assign _T_31 = _T_26 & source_ok; // @[Parameters.scala 1160:30]
  assign _T_37 = $signed(_T_7) & -33'sh1000; // @[Parameters.scala 137:52]
  assign _T_38 = $signed(_T_37) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_39 = io_in_a_bits_address ^ 32'h3000; // @[Parameters.scala 137:31]
  assign _T_40 = {1'b0,$signed(_T_39)}; // @[Parameters.scala 137:49]
  assign _T_42 = $signed(_T_40) & -33'sh1000; // @[Parameters.scala 137:52]
  assign _T_43 = $signed(_T_42) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_44 = io_in_a_bits_address ^ 32'h10000; // @[Parameters.scala 137:31]
  assign _T_45 = {1'b0,$signed(_T_44)}; // @[Parameters.scala 137:49]
  assign _T_47 = $signed(_T_45) & -33'sh10000; // @[Parameters.scala 137:52]
  assign _T_48 = $signed(_T_47) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_49 = io_in_a_bits_address ^ 32'h2000000; // @[Parameters.scala 137:31]
  assign _T_50 = {1'b0,$signed(_T_49)}; // @[Parameters.scala 137:49]
  assign _T_52 = $signed(_T_50) & -33'sh10000; // @[Parameters.scala 137:52]
  assign _T_53 = $signed(_T_52) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_54 = io_in_a_bits_address ^ 32'hc000000; // @[Parameters.scala 137:31]
  assign _T_55 = {1'b0,$signed(_T_54)}; // @[Parameters.scala 137:49]
  assign _T_57 = $signed(_T_55) & -33'sh4000000; // @[Parameters.scala 137:52]
  assign _T_58 = $signed(_T_57) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_59 = io_in_a_bits_address ^ 32'h60000000; // @[Parameters.scala 137:31]
  assign _T_60 = {1'b0,$signed(_T_59)}; // @[Parameters.scala 137:49]
  assign _T_62 = $signed(_T_60) & -33'sh20000000; // @[Parameters.scala 137:52]
  assign _T_63 = $signed(_T_62) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_64 = _T_38 | _T_43; // @[Parameters.scala 671:42]
  assign _T_65 = _T_64 | _T_48; // @[Parameters.scala 671:42]
  assign _T_66 = _T_65 | _T_53; // @[Parameters.scala 671:42]
  assign _T_67 = _T_66 | _T_58; // @[Parameters.scala 671:42]
  assign _T_68 = _T_67 | _T_63; // @[Parameters.scala 671:42]
  assign _T_71 = io_in_a_bits_size <= 4'h6; // @[Parameters.scala 92:42]
  assign _T_74 = io_in_a_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31]
  assign _T_75 = {1'b0,$signed(_T_74)}; // @[Parameters.scala 137:49]
  assign _T_77 = $signed(_T_75) & -33'sh10000000; // @[Parameters.scala 137:52]
  assign _T_78 = $signed(_T_77) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_79 = _T_71 & _T_78; // @[Parameters.scala 670:56]
  assign _T_82 = _T_31 & _T_79; // @[Monitor.scala 82:72]
  assign _T_84 = _T_82 | reset; // @[Monitor.scala 42:11]
  assign _T_88 = 4'h6 == io_in_a_bits_size; // @[Parameters.scala 91:48]
  assign _T_89 = ~io_in_a_bits_source & _T_88; // @[Mux.scala 27:72]
  assign _T_136 = _T_68 | _T_78; // @[Parameters.scala 671:42]
  assign _T_137 = _T_26 & _T_136; // @[Parameters.scala 670:56]
  assign _T_139 = _T_89 & _T_137; // @[Monitor.scala 83:78]
  assign _T_141 = _T_139 | reset; // @[Monitor.scala 42:11]
  assign _T_144 = source_ok | reset; // @[Monitor.scala 42:11]
  assign _T_148 = _mask_T | reset; // @[Monitor.scala 42:11]
  assign _T_151 = is_aligned | reset; // @[Monitor.scala 42:11]
  assign _T_153 = io_in_a_bits_param <= 3'h2; // @[Bundles.scala 108:27]
  assign _T_155 = _T_153 | reset; // @[Monitor.scala 42:11]
  assign _T_158 = ~io_in_a_bits_mask == 8'h0; // @[Monitor.scala 88:31]
  assign _T_160 = _T_158 | reset; // @[Monitor.scala 42:11]
  assign _T_166 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 92:25]
  assign _T_299 = io_in_a_bits_param != 3'h0; // @[Monitor.scala 99:31]
  assign _T_301 = _T_299 | reset; // @[Monitor.scala 42:11]
  assign _T_312 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 104:25]
  assign _T_322 = _T_31 | reset; // @[Monitor.scala 42:11]
  assign _T_333 = _T_26 & _T_43; // @[Parameters.scala 670:56]
  assign _T_368 = _T_38 | _T_48; // @[Parameters.scala 671:42]
  assign _T_369 = _T_368 | _T_53; // @[Parameters.scala 671:42]
  assign _T_370 = _T_369 | _T_58; // @[Parameters.scala 671:42]
  assign _T_371 = _T_370 | _T_63; // @[Parameters.scala 671:42]
  assign _T_372 = _T_371 | _T_78; // @[Parameters.scala 671:42]
  assign _T_373 = _T_71 & _T_372; // @[Parameters.scala 670:56]
  assign _T_375 = _T_333 | _T_373; // @[Parameters.scala 672:30]
  assign _T_377 = _T_375 | reset; // @[Monitor.scala 42:11]
  assign _T_385 = io_in_a_bits_param == 3'h0; // @[Monitor.scala 109:31]
  assign _T_387 = _T_385 | reset; // @[Monitor.scala 42:11]
  assign _T_389 = io_in_a_bits_mask == mask; // @[Monitor.scala 110:30]
  assign _T_391 = _T_389 | reset; // @[Monitor.scala 42:11]
  assign _T_397 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 114:25]
  assign _T_440 = _T_38 | _T_53; // @[Parameters.scala 671:42]
  assign _T_441 = _T_440 | _T_58; // @[Parameters.scala 671:42]
  assign _T_442 = _T_441 | _T_78; // @[Parameters.scala 671:42]
  assign _T_443 = _T_71 & _T_442; // @[Parameters.scala 670:56]
  assign _T_452 = io_in_a_bits_size <= 4'h8; // @[Parameters.scala 92:42]
  assign _T_460 = _T_452 & _T_63; // @[Parameters.scala 670:56]
  assign _T_462 = _T_333 | _T_443; // @[Parameters.scala 672:30]
  assign _T_464 = _T_462 | _T_460; // @[Parameters.scala 672:30]
  assign _T_465 = _T_31 & _T_464; // @[Monitor.scala 115:71]
  assign _T_467 = _T_465 | reset; // @[Monitor.scala 42:11]
  assign _T_483 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 122:25]
  assign _T_566 = io_in_a_bits_mask & ~mask; // @[Monitor.scala 127:31]
  assign _T_567 = _T_566 == 8'h0; // @[Monitor.scala 127:40]
  assign _T_569 = _T_567 | reset; // @[Monitor.scala 42:11]
  assign _T_571 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 130:25]
  assign _T_581 = io_in_a_bits_size <= 4'h3; // @[Parameters.scala 92:42]
  assign _T_605 = _T_64 | _T_53; // @[Parameters.scala 671:42]
  assign _T_606 = _T_605 | _T_58; // @[Parameters.scala 671:42]
  assign _T_607 = _T_581 & _T_606; // @[Parameters.scala 670:56]
  assign _T_629 = _T_31 & _T_607; // @[Monitor.scala 131:74]
  assign _T_631 = _T_629 | reset; // @[Monitor.scala 42:11]
  assign _T_639 = io_in_a_bits_param <= 3'h4; // @[Bundles.scala 138:33]
  assign _T_641 = _T_639 | reset; // @[Monitor.scala 42:11]
  assign _T_647 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 138:25]
  assign _T_715 = io_in_a_bits_param <= 3'h3; // @[Bundles.scala 145:30]
  assign _T_717 = _T_715 | reset; // @[Monitor.scala 42:11]
  assign _T_723 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 146:25]
  assign _T_781 = _T_31 & _T_333; // @[Monitor.scala 147:68]
  assign _T_783 = _T_781 | reset; // @[Monitor.scala 42:11]
  assign _T_791 = io_in_a_bits_param <= 3'h1; // @[Bundles.scala 158:28]
  assign _T_793 = _T_791 | reset; // @[Monitor.scala 42:11]
  assign _T_803 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 42:24]
  assign _T_805 = _T_803 | reset; // @[Monitor.scala 49:11]
  assign source_ok_1 = ~io_in_d_bits_source | io_in_d_bits_source; // @[Parameters.scala 1125:46]
  assign _T_807 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25]
  assign _T_809 = source_ok_1 | reset; // @[Monitor.scala 49:11]
  assign _T_811 = io_in_d_bits_size >= 4'h3; // @[Monitor.scala 312:27]
  assign _T_813 = _T_811 | reset; // @[Monitor.scala 49:11]
  assign _T_815 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 313:28]
  assign _T_817 = _T_815 | reset; // @[Monitor.scala 49:11]
  assign _T_821 = ~io_in_d_bits_corrupt | reset; // @[Monitor.scala 49:11]
  assign _T_825 = ~io_in_d_bits_denied | reset; // @[Monitor.scala 49:11]
  assign _T_827 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25]
  assign _T_838 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 102:26]
  assign _T_840 = _T_838 | reset; // @[Monitor.scala 49:11]
  assign _T_842 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 323:28]
  assign _T_844 = _T_842 | reset; // @[Monitor.scala 49:11]
  assign _T_855 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25]
  assign _T_875 = ~io_in_d_bits_denied | io_in_d_bits_corrupt; // @[Monitor.scala 334:30]
  assign _T_877 = _T_875 | reset; // @[Monitor.scala 49:11]
  assign _T_884 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25]
  assign _T_901 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25]
  assign _T_919 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25]
  assign _T_936 = io_in_b_bits_opcode <= 3'h6; // @[Bundles.scala 40:24]
  assign _T_938 = _T_936 | reset; // @[Monitor.scala 42:11]
  assign _T_943 = {1'b0,$signed(io_in_b_bits_address)}; // @[Parameters.scala 137:49]
  assign _address_ok_T = io_in_b_bits_address ^ 32'h3000; // @[Parameters.scala 137:31]
  assign _address_ok_T_1 = {1'b0,$signed(_address_ok_T)}; // @[Parameters.scala 137:49]
  assign _address_ok_T_3 = $signed(_address_ok_T_1) & -33'sh1000; // @[Parameters.scala 137:52]
  assign _address_ok_T_4 = $signed(_address_ok_T_3) == 33'sh0; // @[Parameters.scala 137:67]
  assign _address_ok_T_5 = io_in_b_bits_address ^ 32'hc000000; // @[Parameters.scala 137:31]
  assign _address_ok_T_6 = {1'b0,$signed(_address_ok_T_5)}; // @[Parameters.scala 137:49]
  assign _address_ok_T_8 = $signed(_address_ok_T_6) & -33'sh4000000; // @[Parameters.scala 137:52]
  assign _address_ok_T_9 = $signed(_address_ok_T_8) == 33'sh0; // @[Parameters.scala 137:67]
  assign _address_ok_T_10 = io_in_b_bits_address ^ 32'h2000000; // @[Parameters.scala 137:31]
  assign _address_ok_T_11 = {1'b0,$signed(_address_ok_T_10)}; // @[Parameters.scala 137:49]
  assign _address_ok_T_13 = $signed(_address_ok_T_11) & -33'sh10000; // @[Parameters.scala 137:52]
  assign _address_ok_T_14 = $signed(_address_ok_T_13) == 33'sh0; // @[Parameters.scala 137:67]
  assign _address_ok_T_18 = $signed(_T_943) & -33'sh1000; // @[Parameters.scala 137:52]
  assign _address_ok_T_19 = $signed(_address_ok_T_18) == 33'sh0; // @[Parameters.scala 137:67]
  assign _address_ok_T_20 = io_in_b_bits_address ^ 32'h10000; // @[Parameters.scala 137:31]
  assign _address_ok_T_21 = {1'b0,$signed(_address_ok_T_20)}; // @[Parameters.scala 137:49]
  assign _address_ok_T_23 = $signed(_address_ok_T_21) & -33'sh10000; // @[Parameters.scala 137:52]
  assign _address_ok_T_24 = $signed(_address_ok_T_23) == 33'sh0; // @[Parameters.scala 137:67]
  assign _address_ok_T_25 = io_in_b_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31]
  assign _address_ok_T_26 = {1'b0,$signed(_address_ok_T_25)}; // @[Parameters.scala 137:49]
  assign _address_ok_T_28 = $signed(_address_ok_T_26) & -33'sh10000000; // @[Parameters.scala 137:52]
  assign _address_ok_T_29 = $signed(_address_ok_T_28) == 33'sh0; // @[Parameters.scala 137:67]
  assign _address_ok_T_30 = io_in_b_bits_address ^ 32'h60000000; // @[Parameters.scala 137:31]
  assign _address_ok_T_31 = {1'b0,$signed(_address_ok_T_30)}; // @[Parameters.scala 137:49]
  assign _address_ok_T_33 = $signed(_address_ok_T_31) & -33'sh20000000; // @[Parameters.scala 137:52]
  assign _address_ok_T_34 = $signed(_address_ok_T_33) == 33'sh0; // @[Parameters.scala 137:67]
  assign _address_ok_T_35 = _address_ok_T_4 | _address_ok_T_9; // @[Parameters.scala 622:64]
  assign _address_ok_T_36 = _address_ok_T_35 | _address_ok_T_14; // @[Parameters.scala 622:64]
  assign _address_ok_T_37 = _address_ok_T_36 | _address_ok_T_19; // @[Parameters.scala 622:64]
  assign _address_ok_T_38 = _address_ok_T_37 | _address_ok_T_24; // @[Parameters.scala 622:64]
  assign _address_ok_T_39 = _address_ok_T_38 | _address_ok_T_29; // @[Parameters.scala 622:64]
  assign address_ok = _address_ok_T_39 | _address_ok_T_34; // @[Parameters.scala 622:64]
  assign _is_aligned_mask_T_4 = 27'hfff << io_in_b_bits_size; // @[package.scala 234:77]
  assign is_aligned_mask_1 = ~_is_aligned_mask_T_4[11:0]; // @[package.scala 234:46]
  assign _GEN_87 = {{20'd0}, is_aligned_mask_1}; // @[Edges.scala 20:16]
  assign _is_aligned_T_1 = io_in_b_bits_address & _GEN_87; // @[Edges.scala 20:16]
  assign is_aligned_1 = _is_aligned_T_1 == 32'h0; // @[Edges.scala 20:24]
  assign mask_sizeOH_shiftAmount_1 = io_in_b_bits_size[1:0]; // @[OneHot.scala 64:49]
  assign _mask_sizeOH_T_4 = 4'h1 << mask_sizeOH_shiftAmount_1; // @[OneHot.scala 65:12]
  assign mask_sizeOH_1 = _mask_sizeOH_T_4[2:0] | 3'h1; // @[Misc.scala 201:81]
  assign _mask_T_1 = io_in_b_bits_size >= 4'h3; // @[Misc.scala 205:21]
  assign mask_size_3 = mask_sizeOH_1[2]; // @[Misc.scala 208:26]
  assign mask_bit_3 = io_in_b_bits_address[2]; // @[Misc.scala 209:26]
  assign mask_nbit_3 = ~mask_bit_3; // @[Misc.scala 210:20]
  assign _mask_acc_T_14 = mask_size_3 & mask_nbit_3; // @[Misc.scala 214:38]
  assign mask_acc_6 = _mask_T_1 | _mask_acc_T_14; // @[Misc.scala 214:29]
  assign _mask_acc_T_15 = mask_size_3 & mask_bit_3; // @[Misc.scala 214:38]
  assign mask_acc_7 = _mask_T_1 | _mask_acc_T_15; // @[Misc.scala 214:29]
  assign mask_size_4 = mask_sizeOH_1[1]; // @[Misc.scala 208:26]
  assign mask_bit_4 = io_in_b_bits_address[1]; // @[Misc.scala 209:26]
  assign mask_nbit_4 = ~mask_bit_4; // @[Misc.scala 210:20]
  assign mask_eq_16 = mask_nbit_3 & mask_nbit_4; // @[Misc.scala 213:27]
  assign _mask_acc_T_16 = mask_size_4 & mask_eq_16; // @[Misc.scala 214:38]
  assign mask_acc_8 = mask_acc_6 | _mask_acc_T_16; // @[Misc.scala 214:29]
  assign mask_eq_17 = mask_nbit_3 & mask_bit_4; // @[Misc.scala 213:27]
  assign _mask_acc_T_17 = mask_size_4 & mask_eq_17; // @[Misc.scala 214:38]
  assign mask_acc_9 = mask_acc_6 | _mask_acc_T_17; // @[Misc.scala 214:29]
  assign mask_eq_18 = mask_bit_3 & mask_nbit_4; // @[Misc.scala 213:27]
  assign _mask_acc_T_18 = mask_size_4 & mask_eq_18; // @[Misc.scala 214:38]
  assign mask_acc_10 = mask_acc_7 | _mask_acc_T_18; // @[Misc.scala 214:29]
  assign mask_eq_19 = mask_bit_3 & mask_bit_4; // @[Misc.scala 213:27]
  assign _mask_acc_T_19 = mask_size_4 & mask_eq_19; // @[Misc.scala 214:38]
  assign mask_acc_11 = mask_acc_7 | _mask_acc_T_19; // @[Misc.scala 214:29]
  assign mask_size_5 = mask_sizeOH_1[0]; // @[Misc.scala 208:26]
  assign mask_bit_5 = io_in_b_bits_address[0]; // @[Misc.scala 209:26]
  assign mask_nbit_5 = ~mask_bit_5; // @[Misc.scala 210:20]
  assign mask_eq_20 = mask_eq_16 & mask_nbit_5; // @[Misc.scala 213:27]
  assign _mask_acc_T_20 = mask_size_5 & mask_eq_20; // @[Misc.scala 214:38]
  assign mask_lo_lo_lo_1 = mask_acc_8 | _mask_acc_T_20; // @[Misc.scala 214:29]
  assign mask_eq_21 = mask_eq_16 & mask_bit_5; // @[Misc.scala 213:27]
  assign _mask_acc_T_21 = mask_size_5 & mask_eq_21; // @[Misc.scala 214:38]
  assign mask_lo_lo_hi_1 = mask_acc_8 | _mask_acc_T_21; // @[Misc.scala 214:29]
  assign mask_eq_22 = mask_eq_17 & mask_nbit_5; // @[Misc.scala 213:27]
  assign _mask_acc_T_22 = mask_size_5 & mask_eq_22; // @[Misc.scala 214:38]
  assign mask_lo_hi_lo_1 = mask_acc_9 | _mask_acc_T_22; // @[Misc.scala 214:29]
  assign mask_eq_23 = mask_eq_17 & mask_bit_5; // @[Misc.scala 213:27]
  assign _mask_acc_T_23 = mask_size_5 & mask_eq_23; // @[Misc.scala 214:38]
  assign mask_lo_hi_hi_1 = mask_acc_9 | _mask_acc_T_23; // @[Misc.scala 214:29]
  assign mask_eq_24 = mask_eq_18 & mask_nbit_5; // @[Misc.scala 213:27]
  assign _mask_acc_T_24 = mask_size_5 & mask_eq_24; // @[Misc.scala 214:38]
  assign mask_hi_lo_lo_1 = mask_acc_10 | _mask_acc_T_24; // @[Misc.scala 214:29]
  assign mask_eq_25 = mask_eq_18 & mask_bit_5; // @[Misc.scala 213:27]
  assign _mask_acc_T_25 = mask_size_5 & mask_eq_25; // @[Misc.scala 214:38]
  assign mask_hi_lo_hi_1 = mask_acc_10 | _mask_acc_T_25; // @[Misc.scala 214:29]
  assign mask_eq_26 = mask_eq_19 & mask_nbit_5; // @[Misc.scala 213:27]
  assign _mask_acc_T_26 = mask_size_5 & mask_eq_26; // @[Misc.scala 214:38]
  assign mask_hi_hi_lo_1 = mask_acc_11 | _mask_acc_T_26; // @[Misc.scala 214:29]
  assign mask_eq_27 = mask_eq_19 & mask_bit_5; // @[Misc.scala 213:27]
  assign _mask_acc_T_27 = mask_size_5 & mask_eq_27; // @[Misc.scala 214:38]
  assign mask_hi_hi_hi_1 = mask_acc_11 | _mask_acc_T_27; // @[Misc.scala 214:29]
  assign mask_1 = {mask_hi_hi_hi_1,mask_hi_hi_lo_1,mask_hi_lo_hi_1,mask_hi_lo_lo_1,mask_lo_hi_hi_1,mask_lo_hi_lo_1,mask_lo_lo_hi_1,mask_lo_lo_lo_1}; // @[Cat.scala 30:58]
  assign legal_source = io_in_b_bits_source == io_in_b_bits_source; // @[Monitor.scala 165:113]
  assign _T_960 = io_in_b_bits_opcode == 3'h6; // @[Monitor.scala 167:25]
  assign _T_963 = 4'h6 == io_in_b_bits_size; // @[Parameters.scala 91:48]
  assign _T_964 = ~io_in_b_bits_source & _T_963; // @[Mux.scala 27:72]
  assign _T_968 = io_in_b_bits_size <= 4'hc; // @[Parameters.scala 92:42]
  assign _T_1006 = _address_ok_T_19 | _address_ok_T_4; // @[Parameters.scala 671:42]
  assign _T_1007 = _T_1006 | _address_ok_T_24; // @[Parameters.scala 671:42]
  assign _T_1008 = _T_1007 | _address_ok_T_14; // @[Parameters.scala 671:42]
  assign _T_1009 = _T_1008 | _address_ok_T_9; // @[Parameters.scala 671:42]
  assign _T_1010 = _T_1009 | _address_ok_T_34; // @[Parameters.scala 671:42]
  assign _T_1011 = _T_1010 | _address_ok_T_29; // @[Parameters.scala 671:42]
  assign _T_1012 = _T_968 & _T_1011; // @[Parameters.scala 670:56]
  assign _T_1014 = _T_964 & _T_1012; // @[Monitor.scala 168:75]
  assign _T_1016 = _T_1014 | reset; // @[Monitor.scala 49:11]
  assign _T_1019 = address_ok | reset; // @[Monitor.scala 49:11]
  assign _T_1022 = legal_source | reset; // @[Monitor.scala 49:11]
  assign _T_1025 = is_aligned_1 | reset; // @[Monitor.scala 49:11]
  assign _T_1027 = io_in_b_bits_param <= 2'h2; // @[Bundles.scala 102:26]
  assign _T_1029 = _T_1027 | reset; // @[Monitor.scala 49:11]
  assign _T_1031 = io_in_b_bits_mask == mask_1; // @[Monitor.scala 173:27]
  assign _T_1033 = _T_1031 | reset; // @[Monitor.scala 49:11]
  assign _T_1037 = ~io_in_b_bits_corrupt | reset; // @[Monitor.scala 49:11]
  assign _T_1039 = io_in_b_bits_opcode == 3'h4; // @[Monitor.scala 177:25]
  assign _T_1100 = io_in_b_bits_param == 2'h0; // @[Monitor.scala 182:31]
  assign _T_1102 = _T_1100 | reset; // @[Monitor.scala 42:11]
  assign _T_1112 = io_in_b_bits_opcode == 3'h0; // @[Monitor.scala 187:25]
  assign _T_1181 = io_in_b_bits_opcode == 3'h1; // @[Monitor.scala 196:25]
  assign _T_1247 = io_in_b_bits_mask & ~mask_1; // @[Monitor.scala 202:31]
  assign _T_1248 = _T_1247 == 8'h0; // @[Monitor.scala 202:40]
  assign _T_1250 = _T_1248 | reset; // @[Monitor.scala 42:11]
  assign _T_1252 = io_in_b_bits_opcode == 3'h2; // @[Monitor.scala 205:25]
  assign _T_1321 = io_in_b_bits_opcode == 3'h3; // @[Monitor.scala 214:25]
  assign _T_1390 = io_in_b_bits_opcode == 3'h5; // @[Monitor.scala 223:25]
  assign source_ok_2 = ~io_in_c_bits_source | io_in_c_bits_source; // @[Parameters.scala 1125:46]
  assign _is_aligned_mask_T_7 = 27'hfff << io_in_c_bits_size; // @[package.scala 234:77]
  assign is_aligned_mask_2 = ~_is_aligned_mask_T_7[11:0]; // @[package.scala 234:46]
  assign _GEN_88 = {{20'd0}, is_aligned_mask_2}; // @[Edges.scala 20:16]
  assign _is_aligned_T_2 = io_in_c_bits_address & _GEN_88; // @[Edges.scala 20:16]
  assign is_aligned_2 = _is_aligned_T_2 == 32'h0; // @[Edges.scala 20:24]
  assign _address_ok_T_40 = io_in_c_bits_address ^ 32'h3000; // @[Parameters.scala 137:31]
  assign _address_ok_T_41 = {1'b0,$signed(_address_ok_T_40)}; // @[Parameters.scala 137:49]
  assign _address_ok_T_43 = $signed(_address_ok_T_41) & -33'sh1000; // @[Parameters.scala 137:52]
  assign _address_ok_T_44 = $signed(_address_ok_T_43) == 33'sh0; // @[Parameters.scala 137:67]
  assign _address_ok_T_45 = io_in_c_bits_address ^ 32'hc000000; // @[Parameters.scala 137:31]
  assign _address_ok_T_46 = {1'b0,$signed(_address_ok_T_45)}; // @[Parameters.scala 137:49]
  assign _address_ok_T_48 = $signed(_address_ok_T_46) & -33'sh4000000; // @[Parameters.scala 137:52]
  assign _address_ok_T_49 = $signed(_address_ok_T_48) == 33'sh0; // @[Parameters.scala 137:67]
  assign _address_ok_T_50 = io_in_c_bits_address ^ 32'h2000000; // @[Parameters.scala 137:31]
  assign _address_ok_T_51 = {1'b0,$signed(_address_ok_T_50)}; // @[Parameters.scala 137:49]
  assign _address_ok_T_53 = $signed(_address_ok_T_51) & -33'sh10000; // @[Parameters.scala 137:52]
  assign _address_ok_T_54 = $signed(_address_ok_T_53) == 33'sh0; // @[Parameters.scala 137:67]
  assign _address_ok_T_56 = {1'b0,$signed(io_in_c_bits_address)}; // @[Parameters.scala 137:49]
  assign _address_ok_T_58 = $signed(_address_ok_T_56) & -33'sh1000; // @[Parameters.scala 137:52]
  assign _address_ok_T_59 = $signed(_address_ok_T_58) == 33'sh0; // @[Parameters.scala 137:67]
  assign _address_ok_T_60 = io_in_c_bits_address ^ 32'h10000; // @[Parameters.scala 137:31]
  assign _address_ok_T_61 = {1'b0,$signed(_address_ok_T_60)}; // @[Parameters.scala 137:49]
  assign _address_ok_T_63 = $signed(_address_ok_T_61) & -33'sh10000; // @[Parameters.scala 137:52]
  assign _address_ok_T_64 = $signed(_address_ok_T_63) == 33'sh0; // @[Parameters.scala 137:67]
  assign _address_ok_T_65 = io_in_c_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31]
  assign _address_ok_T_66 = {1'b0,$signed(_address_ok_T_65)}; // @[Parameters.scala 137:49]
  assign _address_ok_T_68 = $signed(_address_ok_T_66) & -33'sh10000000; // @[Parameters.scala 137:52]
  assign _address_ok_T_69 = $signed(_address_ok_T_68) == 33'sh0; // @[Parameters.scala 137:67]
  assign _address_ok_T_70 = io_in_c_bits_address ^ 32'h60000000; // @[Parameters.scala 137:31]
  assign _address_ok_T_71 = {1'b0,$signed(_address_ok_T_70)}; // @[Parameters.scala 137:49]
  assign _address_ok_T_73 = $signed(_address_ok_T_71) & -33'sh20000000; // @[Parameters.scala 137:52]
  assign _address_ok_T_74 = $signed(_address_ok_T_73) == 33'sh0; // @[Parameters.scala 137:67]
  assign _address_ok_T_75 = _address_ok_T_44 | _address_ok_T_49; // @[Parameters.scala 622:64]
  assign _address_ok_T_76 = _address_ok_T_75 | _address_ok_T_54; // @[Parameters.scala 622:64]
  assign _address_ok_T_77 = _address_ok_T_76 | _address_ok_T_59; // @[Parameters.scala 622:64]
  assign _address_ok_T_78 = _address_ok_T_77 | _address_ok_T_64; // @[Parameters.scala 622:64]
  assign _address_ok_T_79 = _address_ok_T_78 | _address_ok_T_69; // @[Parameters.scala 622:64]
  assign address_ok_1 = _address_ok_T_79 | _address_ok_T_74; // @[Parameters.scala 622:64]
  assign _T_1483 = io_in_c_bits_opcode == 3'h4; // @[Monitor.scala 242:25]
  assign _T_1485 = address_ok_1 | reset; // @[Monitor.scala 42:11]
  assign _T_1488 = source_ok_2 | reset; // @[Monitor.scala 42:11]
  assign _T_1490 = io_in_c_bits_size >= 4'h3; // @[Monitor.scala 245:30]
  assign _T_1492 = _T_1490 | reset; // @[Monitor.scala 42:11]
  assign _T_1495 = is_aligned_2 | reset; // @[Monitor.scala 42:11]
  assign _T_1497 = io_in_c_bits_param <= 3'h5; // @[Bundles.scala 120:29]
  assign _T_1499 = _T_1497 | reset; // @[Monitor.scala 42:11]
  assign _T_1505 = io_in_c_bits_opcode == 3'h5; // @[Monitor.scala 251:25]
  assign _T_1523 = io_in_c_bits_opcode == 3'h6; // @[Monitor.scala 259:25]
  assign _T_1525 = io_in_c_bits_size <= 4'hc; // @[Parameters.scala 92:42]
  assign _T_1530 = _T_1525 & source_ok_2; // @[Parameters.scala 1160:30]
  assign _T_1563 = _address_ok_T_59 | _address_ok_T_44; // @[Parameters.scala 671:42]
  assign _T_1564 = _T_1563 | _address_ok_T_64; // @[Parameters.scala 671:42]
  assign _T_1565 = _T_1564 | _address_ok_T_54; // @[Parameters.scala 671:42]
  assign _T_1566 = _T_1565 | _address_ok_T_49; // @[Parameters.scala 671:42]
  assign _T_1567 = _T_1566 | _address_ok_T_74; // @[Parameters.scala 671:42]
  assign _T_1570 = io_in_c_bits_size <= 4'h6; // @[Parameters.scala 92:42]
  assign _T_1578 = _T_1570 & _address_ok_T_69; // @[Parameters.scala 670:56]
  assign _T_1581 = _T_1530 & _T_1578; // @[Monitor.scala 260:78]
  assign _T_1583 = _T_1581 | reset; // @[Monitor.scala 42:11]
  assign _T_1587 = 4'h6 == io_in_c_bits_size; // @[Parameters.scala 91:48]
  assign _T_1588 = ~io_in_c_bits_source & _T_1587; // @[Mux.scala 27:72]
  assign _T_1635 = _T_1567 | _address_ok_T_69; // @[Parameters.scala 671:42]
  assign _T_1636 = _T_1525 & _T_1635; // @[Parameters.scala 670:56]
  assign _T_1638 = _T_1588 & _T_1636; // @[Monitor.scala 261:78]
  assign _T_1640 = _T_1638 | reset; // @[Monitor.scala 42:11]
  assign _T_1660 = io_in_c_bits_opcode == 3'h7; // @[Monitor.scala 269:25]
  assign _T_1793 = io_in_c_bits_opcode == 3'h0; // @[Monitor.scala 278:25]
  assign _T_1803 = io_in_c_bits_param == 3'h0; // @[Monitor.scala 282:31]
  assign _T_1805 = _T_1803 | reset; // @[Monitor.scala 42:11]
  assign _T_1811 = io_in_c_bits_opcode == 3'h1; // @[Monitor.scala 286:25]
  assign _T_1825 = io_in_c_bits_opcode == 3'h2; // @[Monitor.scala 293:25]
  assign _a_first_T = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37]
  assign a_first_beats1_decode = is_aligned_mask[11:3]; // @[Edges.scala 219:59]
  assign a_first_beats1_opdata = ~io_in_a_bits_opcode[2]; // @[Edges.scala 91:28]
  assign a_first_counter1 = a_first_counter - 9'h1; // @[Edges.scala 229:28]
  assign a_first = a_first_counter == 9'h0; // @[Edges.scala 230:25]
  assign _T_1847 = io_in_a_valid & ~a_first; // @[Monitor.scala 389:19]
  assign _T_1848 = io_in_a_bits_opcode == opcode; // @[Monitor.scala 390:32]
  assign _T_1850 = _T_1848 | reset; // @[Monitor.scala 42:11]
  assign _T_1852 = io_in_a_bits_param == param; // @[Monitor.scala 391:32]
  assign _T_1854 = _T_1852 | reset; // @[Monitor.scala 42:11]
  assign _T_1856 = io_in_a_bits_size == size; // @[Monitor.scala 392:32]
  assign _T_1858 = _T_1856 | reset; // @[Monitor.scala 42:11]
  assign _T_1860 = io_in_a_bits_source == source; // @[Monitor.scala 393:32]
  assign _T_1862 = _T_1860 | reset; // @[Monitor.scala 42:11]
  assign _T_1864 = io_in_a_bits_address == address; // @[Monitor.scala 394:32]
  assign _T_1866 = _T_1864 | reset; // @[Monitor.scala 42:11]
  assign _T_1869 = _a_first_T & a_first; // @[Monitor.scala 396:20]
  assign _d_first_T = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37]
  assign _d_first_beats1_decode_T_1 = 27'hfff << io_in_d_bits_size; // @[package.scala 234:77]
  assign d_first_beats1_decode = ~_d_first_beats1_decode_T_1[11:3]; // @[Edges.scala 219:59]
  assign d_first_beats1_opdata = io_in_d_bits_opcode[0]; // @[Edges.scala 105:36]
  assign d_first_counter1 = d_first_counter - 9'h1; // @[Edges.scala 229:28]
  assign d_first = d_first_counter == 9'h0; // @[Edges.scala 230:25]
  assign _T_1871 = io_in_d_valid & ~d_first; // @[Monitor.scala 541:19]
  assign _T_1872 = io_in_d_bits_opcode == opcode_1; // @[Monitor.scala 542:29]
  assign _T_1874 = _T_1872 | reset; // @[Monitor.scala 49:11]
  assign _T_1876 = io_in_d_bits_param == param_1; // @[Monitor.scala 543:29]
  assign _T_1878 = _T_1876 | reset; // @[Monitor.scala 49:11]
  assign _T_1880 = io_in_d_bits_size == size_1; // @[Monitor.scala 544:29]
  assign _T_1882 = _T_1880 | reset; // @[Monitor.scala 49:11]
  assign _T_1884 = io_in_d_bits_source == source_1; // @[Monitor.scala 545:29]
  assign _T_1886 = _T_1884 | reset; // @[Monitor.scala 49:11]
  assign _T_1888 = io_in_d_bits_sink == sink; // @[Monitor.scala 546:29]
  assign _T_1890 = _T_1888 | reset; // @[Monitor.scala 49:11]
  assign _T_1892 = io_in_d_bits_denied == denied; // @[Monitor.scala 547:29]
  assign _T_1894 = _T_1892 | reset; // @[Monitor.scala 49:11]
  assign _T_1897 = _d_first_T & d_first; // @[Monitor.scala 549:20]
  assign b_first_done = io_in_b_ready & io_in_b_valid; // @[Decoupled.scala 40:37]
  assign b_first_counter1 = b_first_counter - 9'h1; // @[Edges.scala 229:28]
  assign b_first = b_first_counter == 9'h0; // @[Edges.scala 230:25]
  assign _T_1899 = io_in_b_valid & ~b_first; // @[Monitor.scala 412:19]
  assign _T_1900 = io_in_b_bits_opcode == opcode_2; // @[Monitor.scala 413:32]
  assign _T_1902 = _T_1900 | reset; // @[Monitor.scala 42:11]
  assign _T_1904 = io_in_b_bits_param == param_2; // @[Monitor.scala 414:32]
  assign _T_1906 = _T_1904 | reset; // @[Monitor.scala 42:11]
  assign _T_1908 = io_in_b_bits_size == size_2; // @[Monitor.scala 415:32]
  assign _T_1910 = _T_1908 | reset; // @[Monitor.scala 42:11]
  assign _T_1912 = io_in_b_bits_source == source_2; // @[Monitor.scala 416:32]
  assign _T_1914 = _T_1912 | reset; // @[Monitor.scala 42:11]
  assign _T_1916 = io_in_b_bits_address == address_1; // @[Monitor.scala 417:32]
  assign _T_1918 = _T_1916 | reset; // @[Monitor.scala 42:11]
  assign _T_1921 = b_first_done & b_first; // @[Monitor.scala 419:20]
  assign _c_first_T = io_in_c_ready & io_in_c_valid; // @[Decoupled.scala 40:37]
  assign c_first_beats1_decode = is_aligned_mask_2[11:3]; // @[Edges.scala 219:59]
  assign c_first_beats1_opdata = io_in_c_bits_opcode[0]; // @[Edges.scala 101:36]
  assign c_first_counter1 = c_first_counter - 9'h1; // @[Edges.scala 229:28]
  assign c_first = c_first_counter == 9'h0; // @[Edges.scala 230:25]
  assign _T_1923 = io_in_c_valid & ~c_first; // @[Monitor.scala 517:19]
  assign _T_1924 = io_in_c_bits_opcode == opcode_3; // @[Monitor.scala 518:32]
  assign _T_1926 = _T_1924 | reset; // @[Monitor.scala 42:11]
  assign _T_1928 = io_in_c_bits_param == param_3; // @[Monitor.scala 519:32]
  assign _T_1930 = _T_1928 | reset; // @[Monitor.scala 42:11]
  assign _T_1932 = io_in_c_bits_size == size_3; // @[Monitor.scala 520:32]
  assign _T_1934 = _T_1932 | reset; // @[Monitor.scala 42:11]
  assign _T_1936 = io_in_c_bits_source == source_3; // @[Monitor.scala 521:32]
  assign _T_1938 = _T_1936 | reset; // @[Monitor.scala 42:11]
  assign _T_1940 = io_in_c_bits_address == address_2; // @[Monitor.scala 522:32]
  assign _T_1942 = _T_1940 | reset; // @[Monitor.scala 42:11]
  assign _T_1945 = _c_first_T & c_first; // @[Monitor.scala 524:20]
  assign a_first_counter1_1 = a_first_counter_1 - 9'h1; // @[Edges.scala 229:28]
  assign a_first_1 = a_first_counter_1 == 9'h0; // @[Edges.scala 230:25]
  assign d_first_counter1_1 = d_first_counter_1 - 9'h1; // @[Edges.scala 229:28]
  assign d_first_1 = d_first_counter_1 == 9'h0; // @[Edges.scala 230:25]
  assign _GEN_89 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 634:69]
  assign _a_opcode_lookup_T = {{1'd0}, _GEN_89}; // @[Monitor.scala 634:69]
  assign _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T; // @[Monitor.scala 634:44]
  assign _a_opcode_lookup_T_5 = 16'h10 - 16'h1; // @[Monitor.scala 609:57]
  assign _GEN_90 = {{8'd0}, _a_opcode_lookup_T_1}; // @[Monitor.scala 634:97]
  assign _a_opcode_lookup_T_6 = _GEN_90 & _a_opcode_lookup_T_5; // @[Monitor.scala 634:97]
  assign _a_opcode_lookup_T_7 = {{1'd0}, _a_opcode_lookup_T_6[15:1]}; // @[Monitor.scala 634:152]
  assign _a_size_lookup_T = {io_in_d_bits_source, 3'h0}; // @[Monitor.scala 638:65]
  assign _a_size_lookup_T_1 = inflight_sizes >> _a_size_lookup_T; // @[Monitor.scala 638:40]
  assign _a_size_lookup_T_5 = 16'h100 - 16'h1; // @[Monitor.scala 609:57]
  assign _a_size_lookup_T_6 = _a_size_lookup_T_1 & _a_size_lookup_T_5; // @[Monitor.scala 638:91]
  assign _a_size_lookup_T_7 = {{1'd0}, _a_size_lookup_T_6[15:1]}; // @[Monitor.scala 638:144]
  assign _T_1946 = io_in_a_valid & a_first_1; // @[Monitor.scala 648:26]
  assign _a_set_wo_ready_T = 2'h1 << io_in_a_bits_source; // @[OneHot.scala 58:35]
  assign a_set_wo_ready = _T_1946 ? _a_set_wo_ready_T : 2'h0; // @[Monitor.scala 648:71]
  assign _T_1949 = _a_first_T & a_first_1; // @[Monitor.scala 652:27]
  assign _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 654:53]
  assign _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1; // @[Monitor.scala 654:61]
  assign _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 655:51]
  assign _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 5'h1; // @[Monitor.scala 655:59]
  assign _GEN_93 = {io_in_a_bits_source, 2'h0}; // @[Monitor.scala 656:79]
  assign _a_opcodes_set_T = {{1'd0}, _GEN_93}; // @[Monitor.scala 656:79]
  assign a_opcodes_set_interm = _T_1949 ? _a_opcodes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72]
  assign _GEN_94 = {{15'd0}, a_opcodes_set_interm}; // @[Monitor.scala 656:54]
  assign _a_opcodes_set_T_1 = _GEN_94 << _a_opcodes_set_T; // @[Monitor.scala 656:54]
  assign _a_sizes_set_T = {io_in_a_bits_source, 3'h0}; // @[Monitor.scala 657:77]
  assign a_sizes_set_interm = _T_1949 ? _a_sizes_set_interm_T_1 : 5'h0; // @[Monitor.scala 652:72]
  assign _GEN_95 = {{15'd0}, a_sizes_set_interm}; // @[Monitor.scala 657:52]
  assign _a_sizes_set_T_1 = _GEN_95 << _a_sizes_set_T; // @[Monitor.scala 657:52]
  assign _T_1951 = inflight >> io_in_a_bits_source; // @[Monitor.scala 658:26]
  assign _T_1955 = ~_T_1951[0] | reset; // @[Monitor.scala 42:11]
  assign a_set = _T_1949 ? _a_set_wo_ready_T : 2'h0; // @[Monitor.scala 652:72]
  assign _GEN_31 = _T_1949 ? _a_opcodes_set_T_1 : 19'h0; // @[Monitor.scala 652:72]
  assign _GEN_32 = _T_1949 ? _a_sizes_set_T_1 : 20'h0; // @[Monitor.scala 652:72]
  assign _T_1957 = io_in_d_valid & d_first_1; // @[Monitor.scala 671:26]
  assign _T_1960 = _T_1957 & ~_T_807; // @[Monitor.scala 671:71]
  assign _d_clr_wo_ready_T = 2'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35]
  assign d_clr_wo_ready = _T_1960 ? _d_clr_wo_ready_T : 2'h0; // @[Monitor.scala 671:90]
  assign _T_1962 = _d_first_T & d_first_1; // @[Monitor.scala 675:27]
  assign _T_1965 = _T_1962 & ~_T_807; // @[Monitor.scala 675:72]
  assign _GEN_97 = {{15'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 677:76]
  assign _d_opcodes_clr_T_5 = _GEN_97 << _a_opcode_lookup_T; // @[Monitor.scala 677:76]
  assign _GEN_98 = {{15'd0}, _a_size_lookup_T_5}; // @[Monitor.scala 678:74]
  assign _d_sizes_clr_T_5 = _GEN_98 << _a_size_lookup_T; // @[Monitor.scala 678:74]
  assign d_clr = _T_1965 ? _d_clr_wo_ready_T : 2'h0; // @[Monitor.scala 675:91]
  assign _GEN_35 = _T_1965 ? _d_opcodes_clr_T_5 : 31'h0; // @[Monitor.scala 675:91]
  assign _GEN_36 = _T_1965 ? _d_sizes_clr_T_5 : 31'h0; // @[Monitor.scala 675:91]
  assign _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:113]
  assign same_cycle_resp = _T_1946 & _same_cycle_resp_T_2; // @[Monitor.scala 681:88]
  assign _T_1970 = inflight >> io_in_d_bits_source; // @[Monitor.scala 682:25]
  assign _T_1972 = _T_1970[0] | same_cycle_resp; // @[Monitor.scala 682:49]
  assign _T_1974 = _T_1972 | reset; // @[Monitor.scala 49:11]
  assign _GEN_39 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 685:38]
  assign _GEN_40 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_39; // @[Monitor.scala 685:38]
  assign _GEN_41 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_40; // @[Monitor.scala 685:38]
  assign _GEN_42 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_41; // @[Monitor.scala 685:38]
  assign _GEN_43 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_42; // @[Monitor.scala 685:38]
  assign _GEN_44 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_43; // @[Monitor.scala 685:38]
  assign _T_1976 = io_in_d_bits_opcode == _GEN_44; // @[Monitor.scala 685:38]
  assign _GEN_51 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_42; // @[Monitor.scala 686:39]
  assign _GEN_52 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_51; // @[Monitor.scala 686:39]
  assign _T_1977 = io_in_d_bits_opcode == _GEN_52; // @[Monitor.scala 686:39]
  assign _T_1978 = _T_1976 | _T_1977; // @[Monitor.scala 685:77]
  assign _T_1980 = _T_1978 | reset; // @[Monitor.scala 49:11]
  assign _T_1982 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 687:36]
  assign _T_1984 = _T_1982 | reset; // @[Monitor.scala 49:11]
  assign a_opcode_lookup = _a_opcode_lookup_T_7[3:0]; // @[Monitor.scala 634:21]
  assign _GEN_55 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 689:38]
  assign _GEN_56 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_55; // @[Monitor.scala 689:38]
  assign _GEN_57 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_56; // @[Monitor.scala 689:38]
  assign _GEN_58 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_57; // @[Monitor.scala 689:38]
  assign _GEN_59 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_58; // @[Monitor.scala 689:38]
  assign _GEN_60 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_59; // @[Monitor.scala 689:38]
  assign _T_1987 = io_in_d_bits_opcode == _GEN_60; // @[Monitor.scala 689:38]
  assign _GEN_67 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_58; // @[Monitor.scala 690:38]
  assign _GEN_68 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_67; // @[Monitor.scala 690:38]
  assign _T_1989 = io_in_d_bits_opcode == _GEN_68; // @[Monitor.scala 690:38]
  assign _T_1990 = _T_1987 | _T_1989; // @[Monitor.scala 689:72]
  assign _T_1992 = _T_1990 | reset; // @[Monitor.scala 49:11]
  assign a_size_lookup = _a_size_lookup_T_7[7:0]; // @[Monitor.scala 638:19]
  assign _GEN_99 = {{4'd0}, io_in_d_bits_size}; // @[Monitor.scala 691:36]
  assign _T_1994 = _GEN_99 == a_size_lookup; // @[Monitor.scala 691:36]
  assign _T_1996 = _T_1994 | reset; // @[Monitor.scala 49:11]
  assign _T_1999 = _T_1957 & a_first_1; // @[Monitor.scala 694:36]
  assign _T_2000 = _T_1999 & io_in_a_valid; // @[Monitor.scala 694:47]
  assign _T_2002 = _T_2000 & _same_cycle_resp_T_2; // @[Monitor.scala 694:65]
  assign _T_2004 = _T_2002 & ~_T_807; // @[Monitor.scala 694:116]
  assign _T_2006 = ~io_in_d_ready | io_in_a_ready; // @[Monitor.scala 695:32]
  assign _T_2008 = _T_2006 | reset; // @[Monitor.scala 49:11]
  assign _T_2010 = a_set_wo_ready != d_clr_wo_ready; // @[Monitor.scala 699:29]
  assign _T_2011 = |a_set_wo_ready; // @[Monitor.scala 699:67]
  assign _T_2013 = _T_2010 | ~_T_2011; // @[Monitor.scala 699:48]
  assign _T_2015 = _T_2013 | reset; // @[Monitor.scala 49:11]
  assign _inflight_T = inflight | a_set; // @[Monitor.scala 702:27]
  assign _inflight_T_2 = _inflight_T & ~d_clr; // @[Monitor.scala 702:36]
  assign a_opcodes_set = _GEN_31[7:0]; // @[Monitor.scala 656:28]
  assign _inflight_opcodes_T = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 703:43]
  assign d_opcodes_clr = _GEN_35[7:0]; // @[Monitor.scala 677:21]
  assign _inflight_opcodes_T_2 = _inflight_opcodes_T & ~d_opcodes_clr; // @[Monitor.scala 703:60]
  assign a_sizes_set = _GEN_32[15:0]; // @[Monitor.scala 657:28]
  assign _inflight_sizes_T = inflight_sizes | a_sizes_set; // @[Monitor.scala 704:39]
  assign d_sizes_clr = _GEN_36[15:0]; // @[Monitor.scala 678:21]
  assign _inflight_sizes_T_2 = _inflight_sizes_T & ~d_sizes_clr; // @[Monitor.scala 704:54]
  assign _T_2017 = |inflight; // @[Monitor.scala 709:26]
  assign _T_2019 = plusarg_reader_out == 32'h0; // @[Monitor.scala 709:39]
  assign _T_2020 = ~_T_2017 | _T_2019; // @[Monitor.scala 709:30]
  assign _T_2021 = watchdog < plusarg_reader_out; // @[Monitor.scala 709:59]
  assign _T_2022 = _T_2020 | _T_2021; // @[Monitor.scala 709:47]
  assign _T_2024 = _T_2022 | reset; // @[Monitor.scala 42:11]
  assign _watchdog_T_1 = watchdog + 32'h1; // @[Monitor.scala 711:26]
  assign _T_2028 = _a_first_T | _d_first_T; // @[Monitor.scala 712:27]
  assign c_first_counter1_1 = c_first_counter_1 - 9'h1; // @[Edges.scala 229:28]
  assign c_first_1 = c_first_counter_1 == 9'h0; // @[Edges.scala 230:25]
  assign d_first_counter1_2 = d_first_counter_2 - 9'h1; // @[Edges.scala 229:28]
  assign d_first_2 = d_first_counter_2 == 9'h0; // @[Edges.scala 230:25]
  assign _c_size_lookup_T_1 = inflight_sizes_1 >> _a_size_lookup_T; // @[Monitor.scala 747:42]
  assign _c_size_lookup_T_6 = _c_size_lookup_T_1 & _a_size_lookup_T_5; // @[Monitor.scala 747:93]
  assign _c_size_lookup_T_7 = {{1'd0}, _c_size_lookup_T_6[15:1]}; // @[Monitor.scala 747:146]
  assign _T_2029 = io_in_c_valid & c_first_1; // @[Monitor.scala 756:26]
  assign _T_2032 = io_in_c_bits_opcode[2] & io_in_c_bits_opcode[1]; // @[Edges.scala 67:40]
  assign _T_2033 = _T_2029 & _T_2032; // @[Monitor.scala 756:37]
  assign _c_set_wo_ready_T = 2'h1 << io_in_c_bits_source; // @[OneHot.scala 58:35]
  assign c_set_wo_ready = _T_2033 ? _c_set_wo_ready_T : 2'h0; // @[Monitor.scala 756:71]
  assign _T_2035 = _c_first_T & c_first_1; // @[Monitor.scala 760:27]
  assign _T_2039 = _T_2035 & _T_2032; // @[Monitor.scala 760:38]
  assign _c_sizes_set_interm_T = {io_in_c_bits_size, 1'h0}; // @[Monitor.scala 763:51]
  assign _c_sizes_set_interm_T_1 = _c_sizes_set_interm_T | 5'h1; // @[Monitor.scala 763:59]
  assign _c_sizes_set_T = {io_in_c_bits_source, 3'h0}; // @[Monitor.scala 765:77]
  assign c_sizes_set_interm = _T_2039 ? _c_sizes_set_interm_T_1 : 5'h0; // @[Monitor.scala 760:72]
  assign _GEN_106 = {{15'd0}, c_sizes_set_interm}; // @[Monitor.scala 765:52]
  assign _c_sizes_set_T_1 = _GEN_106 << _c_sizes_set_T; // @[Monitor.scala 765:52]
  assign _T_2040 = inflight_1 >> io_in_c_bits_source; // @[Monitor.scala 766:26]
  assign _T_2044 = ~_T_2040[0] | reset; // @[Monitor.scala 42:11]
  assign c_set = _T_2039 ? _c_set_wo_ready_T : 2'h0; // @[Monitor.scala 760:72]
  assign _GEN_77 = _T_2039 ? _c_sizes_set_T_1 : 20'h0; // @[Monitor.scala 760:72]
  assign _T_2046 = io_in_d_valid & d_first_2; // @[Monitor.scala 779:26]
  assign _T_2048 = _T_2046 & _T_807; // @[Monitor.scala 779:71]
  assign d_clr_wo_ready_1 = _T_2048 ? _d_clr_wo_ready_T : 2'h0; // @[Monitor.scala 779:89]
  assign _T_2050 = _d_first_T & d_first_2; // @[Monitor.scala 783:27]
  assign _T_2052 = _T_2050 & _T_807; // @[Monitor.scala 783:72]
  assign d_clr_1 = _T_2052 ? _d_clr_wo_ready_T : 2'h0; // @[Monitor.scala 783:90]
  assign _GEN_81 = _T_2052 ? _d_sizes_clr_T_5 : 31'h0; // @[Monitor.scala 783:90]
  assign _same_cycle_resp_T_8 = io_in_c_bits_source == io_in_d_bits_source; // @[Monitor.scala 790:113]
  assign same_cycle_resp_1 = _T_2033 & _same_cycle_resp_T_8; // @[Monitor.scala 790:88]
  assign _T_2056 = inflight_1 >> io_in_d_bits_source; // @[Monitor.scala 791:25]
  assign _T_2058 = _T_2056[0] | same_cycle_resp_1; // @[Monitor.scala 791:49]
  assign _T_2060 = _T_2058 | reset; // @[Monitor.scala 49:11]
  assign _T_2062 = io_in_d_bits_size == io_in_c_bits_size; // @[Monitor.scala 793:36]
  assign _T_2064 = _T_2062 | reset; // @[Monitor.scala 49:11]
  assign c_size_lookup = _c_size_lookup_T_7[7:0]; // @[Monitor.scala 747:21]
  assign _T_2066 = _GEN_99 == c_size_lookup; // @[Monitor.scala 795:36]
  assign _T_2068 = _T_2066 | reset; // @[Monitor.scala 49:11]
  assign _T_2071 = _T_2046 & c_first_1; // @[Monitor.scala 799:36]
  assign _T_2072 = _T_2071 & io_in_c_valid; // @[Monitor.scala 799:47]
  assign _T_2074 = _T_2072 & _same_cycle_resp_T_8; // @[Monitor.scala 799:65]
  assign _T_2075 = _T_2074 & _T_807; // @[Monitor.scala 799:116]
  assign _T_2077 = ~io_in_d_ready | io_in_c_ready; // @[Monitor.scala 800:32]
  assign _T_2079 = _T_2077 | reset; // @[Monitor.scala 49:11]
  assign _T_2081 = |c_set_wo_ready; // @[Monitor.scala 804:28]
  assign _T_2082 = c_set_wo_ready != d_clr_wo_ready_1; // @[Monitor.scala 805:31]
  assign _T_2084 = _T_2082 | reset; // @[Monitor.scala 49:11]
  assign _inflight_T_3 = inflight_1 | c_set; // @[Monitor.scala 809:35]
  assign _inflight_T_5 = _inflight_T_3 & ~d_clr_1; // @[Monitor.scala 809:44]
  assign c_sizes_set = _GEN_77[15:0]; // @[Monitor.scala 765:28]
  assign _inflight_sizes_T_3 = inflight_sizes_1 | c_sizes_set; // @[Monitor.scala 811:41]
  assign d_sizes_clr_1 = _GEN_81[15:0]; // @[Monitor.scala 786:21]
  assign _inflight_sizes_T_5 = _inflight_sizes_T_3 & ~d_sizes_clr_1; // @[Monitor.scala 811:56]
  assign _T_2086 = |inflight_1; // @[Monitor.scala 816:26]
  assign _T_2088 = plusarg_reader_1_out == 32'h0; // @[Monitor.scala 816:39]
  assign _T_2089 = ~_T_2086 | _T_2088; // @[Monitor.scala 816:30]
  assign _T_2090 = watchdog_1 < plusarg_reader_1_out; // @[Monitor.scala 816:59]
  assign _T_2091 = _T_2089 | _T_2090; // @[Monitor.scala 816:47]
  assign _T_2093 = _T_2091 | reset; // @[Monitor.scala 42:11]
  assign _watchdog_T_3 = watchdog_1 + 32'h1; // @[Monitor.scala 818:26]
  assign _T_2097 = _c_first_T | _d_first_T; // @[Monitor.scala 819:27]
  assign d_first_counter1_3 = d_first_counter_3 - 9'h1; // @[Edges.scala 229:28]
  assign d_first_3 = d_first_counter_3 == 9'h0; // @[Edges.scala 230:25]
  assign _T_2099 = _d_first_T & d_first_3; // @[Monitor.scala 829:27]
  assign _T_2103 = io_in_d_bits_opcode[2] & ~io_in_d_bits_opcode[1]; // @[Edges.scala 70:40]
  assign _T_2104 = _T_2099 & _T_2103; // @[Monitor.scala 829:38]
  assign _d_set_T = 4'h1 << io_in_d_bits_sink; // @[OneHot.scala 58:35]
  assign _T_2105 = inflight_2 >> io_in_d_bits_sink; // @[Monitor.scala 831:23]
  assign _T_2109 = ~_T_2105[0] | reset; // @[Monitor.scala 49:11]
  assign d_set = _T_2104 ? _d_set_T : 4'h0; // @[Monitor.scala 829:72]
  assign _T_2111 = io_in_e_ready & io_in_e_valid; // @[Decoupled.scala 40:37]
  assign _e_clr_T = 4'h1 << io_in_e_bits_sink; // @[OneHot.scala 58:35]
  assign _T_2114 = d_set | inflight_2; // @[Monitor.scala 837:24]
  assign _T_2115 = _T_2114 >> io_in_e_bits_sink; // @[Monitor.scala 837:35]
  assign _T_2118 = _T_2115[0] | reset; // @[Monitor.scala 42:11]
  assign e_clr = _T_2111 ? _e_clr_T : 4'h0; // @[Monitor.scala 835:73]
  assign _inflight_T_6 = inflight_2 | d_set; // @[Monitor.scala 842:27]
  assign _inflight_T_8 = _inflight_T_6 & ~e_clr; // @[Monitor.scala 842:36]
  assign _GEN_111 = io_in_a_valid & _T_24; // @[Monitor.scala 42:11]
  assign _GEN_125 = io_in_a_valid & _T_166; // @[Monitor.scala 42:11]
  assign _GEN_141 = io_in_a_valid & _T_312; // @[Monitor.scala 42:11]
  assign _GEN_153 = io_in_a_valid & _T_397; // @[Monitor.scala 42:11]
  assign _GEN_163 = io_in_a_valid & _T_483; // @[Monitor.scala 42:11]
  assign _GEN_173 = io_in_a_valid & _T_571; // @[Monitor.scala 42:11]
  assign _GEN_183 = io_in_a_valid & _T_647; // @[Monitor.scala 42:11]
  assign _GEN_193 = io_in_a_valid & _T_723; // @[Monitor.scala 42:11]
  assign _GEN_203 = io_in_d_valid & _T_807; // @[Monitor.scala 49:11]
  assign _GEN_213 = io_in_d_valid & _T_827; // @[Monitor.scala 49:11]
  assign _GEN_223 = io_in_d_valid & _T_855; // @[Monitor.scala 49:11]
  assign _GEN_233 = io_in_d_valid & _T_884; // @[Monitor.scala 49:11]
  assign _GEN_239 = io_in_d_valid & _T_901; // @[Monitor.scala 49:11]
  assign _GEN_245 = io_in_d_valid & _T_919; // @[Monitor.scala 49:11]
  assign _GEN_251 = io_in_b_valid & _T_960; // @[Monitor.scala 49:11]
  assign _GEN_265 = io_in_b_valid & _T_1039; // @[Monitor.scala 42:11]
  assign _GEN_279 = io_in_b_valid & _T_1112; // @[Monitor.scala 42:11]
  assign _GEN_291 = io_in_b_valid & _T_1181; // @[Monitor.scala 42:11]
  assign _GEN_303 = io_in_b_valid & _T_1252; // @[Monitor.scala 42:11]
  assign _GEN_313 = io_in_b_valid & _T_1321; // @[Monitor.scala 42:11]
  assign _GEN_323 = io_in_b_valid & _T_1390; // @[Monitor.scala 42:11]
  assign _GEN_335 = io_in_c_valid & _T_1483; // @[Monitor.scala 42:11]
  assign _GEN_345 = io_in_c_valid & _T_1505; // @[Monitor.scala 42:11]
  assign _GEN_355 = io_in_c_valid & _T_1523; // @[Monitor.scala 42:11]
  assign _GEN_367 = io_in_c_valid & _T_1660; // @[Monitor.scala 42:11]
  assign _GEN_379 = io_in_c_valid & _T_1793; // @[Monitor.scala 42:11]
  assign _GEN_387 = io_in_c_valid & _T_1811; // @[Monitor.scala 42:11]
  assign _GEN_395 = io_in_c_valid & _T_1825; // @[Monitor.scala 42:11]
  assign _GEN_403 = _T_1960 & same_cycle_resp; // @[Monitor.scala 49:11]
  assign _GEN_408 = _T_1960 & ~same_cycle_resp; // @[Monitor.scala 49:11]
  assign _GEN_415 = _T_2048 & same_cycle_resp_1; // @[Monitor.scala 49:11]
  assign _GEN_418 = _T_2048 & ~same_cycle_resp_1; // @[Monitor.scala 49:11]
  assign TLMonitor_23_covSum = 30'h0;
  assign io_covSum = TLMonitor_23_covSum;
  assign stopEn0 = _GEN_111 & ~_T_84;
  assign stopEn1 = _GEN_111 & ~_T_141;
  assign stopEn2 = _GEN_111 & ~_T_144;
  assign stopEn3 = _GEN_111 & ~_T_148;
  assign stopEn4 = _GEN_111 & ~_T_151;
  assign stopEn5 = _GEN_111 & ~_T_155;
  assign stopEn6 = _GEN_111 & ~_T_160;
  assign stopEn7 = _GEN_125 & ~_T_84;
  assign stopEn8 = _GEN_125 & ~_T_141;
  assign stopEn9 = _GEN_125 & ~_T_144;
  assign stopEn10 = _GEN_125 & ~_T_148;
  assign stopEn11 = _GEN_125 & ~_T_151;
  assign stopEn12 = _GEN_125 & ~_T_155;
  assign stopEn13 = _GEN_125 & ~_T_301;
  assign stopEn14 = _GEN_125 & ~_T_160;
  assign stopEn15 = _GEN_141 & ~_T_322;
  assign stopEn16 = _GEN_141 & ~_T_377;
  assign stopEn17 = _GEN_141 & ~_T_144;
  assign stopEn18 = _GEN_141 & ~_T_151;
  assign stopEn19 = _GEN_141 & ~_T_387;
  assign stopEn20 = _GEN_141 & ~_T_391;
  assign stopEn21 = _GEN_153 & ~_T_467;
  assign stopEn22 = _GEN_153 & ~_T_144;
  assign stopEn23 = _GEN_153 & ~_T_151;
  assign stopEn24 = _GEN_153 & ~_T_387;
  assign stopEn25 = _GEN_153 & ~_T_391;
  assign stopEn26 = _GEN_163 & ~_T_467;
  assign stopEn27 = _GEN_163 & ~_T_144;
  assign stopEn28 = _GEN_163 & ~_T_151;
  assign stopEn29 = _GEN_163 & ~_T_387;
  assign stopEn30 = _GEN_163 & ~_T_569;
  assign stopEn31 = _GEN_173 & ~_T_631;
  assign stopEn32 = _GEN_173 & ~_T_144;
  assign stopEn33 = _GEN_173 & ~_T_151;
  assign stopEn34 = _GEN_173 & ~_T_641;
  assign stopEn35 = _GEN_173 & ~_T_391;
  assign stopEn36 = _GEN_183 & ~_T_631;
  assign stopEn37 = _GEN_183 & ~_T_144;
  assign stopEn38 = _GEN_183 & ~_T_151;
  assign stopEn39 = _GEN_183 & ~_T_717;
  assign stopEn40 = _GEN_183 & ~_T_391;
  assign stopEn41 = _GEN_193 & ~_T_783;
  assign stopEn42 = _GEN_193 & ~_T_144;
  assign stopEn43 = _GEN_193 & ~_T_151;
  assign stopEn44 = _GEN_193 & ~_T_793;
  assign stopEn45 = _GEN_193 & ~_T_391;
  assign stopEn46 = io_in_d_valid & ~_T_805;
  assign stopEn47 = _GEN_203 & ~_T_809;
  assign stopEn48 = _GEN_203 & ~_T_813;
  assign stopEn49 = _GEN_203 & ~_T_817;
  assign stopEn50 = _GEN_203 & ~_T_821;
  assign stopEn51 = _GEN_203 & ~_T_825;
  assign stopEn52 = _GEN_213 & ~_T_809;
  assign stopEn53 = _GEN_213 & ~_T_813;
  assign stopEn54 = _GEN_213 & ~_T_840;
  assign stopEn55 = _GEN_213 & ~_T_844;
  assign stopEn56 = _GEN_213 & ~_T_821;
  assign stopEn57 = _GEN_223 & ~_T_809;
  assign stopEn58 = _GEN_223 & ~_T_813;
  assign stopEn59 = _GEN_223 & ~_T_840;
  assign stopEn60 = _GEN_223 & ~_T_844;
  assign stopEn61 = _GEN_223 & ~_T_877;
  assign stopEn62 = _GEN_233 & ~_T_809;
  assign stopEn63 = _GEN_233 & ~_T_817;
  assign stopEn64 = _GEN_233 & ~_T_821;
  assign stopEn65 = _GEN_239 & ~_T_809;
  assign stopEn66 = _GEN_239 & ~_T_817;
  assign stopEn67 = _GEN_239 & ~_T_877;
  assign stopEn68 = _GEN_245 & ~_T_809;
  assign stopEn69 = _GEN_245 & ~_T_817;
  assign stopEn70 = _GEN_245 & ~_T_821;
  assign stopEn71 = io_in_b_valid & ~_T_938;
  assign stopEn72 = _GEN_251 & ~_T_1016;
  assign stopEn73 = _GEN_251 & ~_T_1019;
  assign stopEn74 = _GEN_251 & ~_T_1022;
  assign stopEn75 = _GEN_251 & ~_T_1025;
  assign stopEn76 = _GEN_251 & ~_T_1029;
  assign stopEn77 = _GEN_251 & ~_T_1033;
  assign stopEn78 = _GEN_251 & ~_T_1037;
  assign stopEn79 = _GEN_265 & ~reset;
  assign stopEn80 = _GEN_265 & ~_T_1019;
  assign stopEn81 = _GEN_265 & ~_T_1022;
  assign stopEn82 = _GEN_265 & ~_T_1025;
  assign stopEn83 = _GEN_265 & ~_T_1102;
  assign stopEn84 = _GEN_265 & ~_T_1033;
  assign stopEn85 = _GEN_265 & ~_T_1037;
  assign stopEn86 = _GEN_279 & ~reset;
  assign stopEn87 = _GEN_279 & ~_T_1019;
  assign stopEn88 = _GEN_279 & ~_T_1022;
  assign stopEn89 = _GEN_279 & ~_T_1025;
  assign stopEn90 = _GEN_279 & ~_T_1102;
  assign stopEn91 = _GEN_279 & ~_T_1033;
  assign stopEn92 = _GEN_291 & ~reset;
  assign stopEn93 = _GEN_291 & ~_T_1019;
  assign stopEn94 = _GEN_291 & ~_T_1022;
  assign stopEn95 = _GEN_291 & ~_T_1025;
  assign stopEn96 = _GEN_291 & ~_T_1102;
  assign stopEn97 = _GEN_291 & ~_T_1250;
  assign stopEn98 = _GEN_303 & ~reset;
  assign stopEn99 = _GEN_303 & ~_T_1019;
  assign stopEn100 = _GEN_303 & ~_T_1022;
  assign stopEn101 = _GEN_303 & ~_T_1025;
  assign stopEn102 = _GEN_303 & ~_T_1033;
  assign stopEn103 = _GEN_313 & ~reset;
  assign stopEn104 = _GEN_313 & ~_T_1019;
  assign stopEn105 = _GEN_313 & ~_T_1022;
  assign stopEn106 = _GEN_313 & ~_T_1025;
  assign stopEn107 = _GEN_313 & ~_T_1033;
  assign stopEn108 = _GEN_323 & ~reset;
  assign stopEn109 = _GEN_323 & ~_T_1019;
  assign stopEn110 = _GEN_323 & ~_T_1022;
  assign stopEn111 = _GEN_323 & ~_T_1025;
  assign stopEn112 = _GEN_323 & ~_T_1033;
  assign stopEn113 = _GEN_323 & ~_T_1037;
  assign stopEn114 = _GEN_335 & ~_T_1485;
  assign stopEn115 = _GEN_335 & ~_T_1488;
  assign stopEn116 = _GEN_335 & ~_T_1492;
  assign stopEn117 = _GEN_335 & ~_T_1495;
  assign stopEn118 = _GEN_335 & ~_T_1499;
  assign stopEn119 = _GEN_345 & ~_T_1485;
  assign stopEn120 = _GEN_345 & ~_T_1488;
  assign stopEn121 = _GEN_345 & ~_T_1492;
  assign stopEn122 = _GEN_345 & ~_T_1495;
  assign stopEn123 = _GEN_345 & ~_T_1499;
  assign stopEn124 = _GEN_355 & ~_T_1583;
  assign stopEn125 = _GEN_355 & ~_T_1640;
  assign stopEn126 = _GEN_355 & ~_T_1488;
  assign stopEn127 = _GEN_355 & ~_T_1492;
  assign stopEn128 = _GEN_355 & ~_T_1495;
  assign stopEn129 = _GEN_355 & ~_T_1499;
  assign stopEn130 = _GEN_367 & ~_T_1583;
  assign stopEn131 = _GEN_367 & ~_T_1640;
  assign stopEn132 = _GEN_367 & ~_T_1488;
  assign stopEn133 = _GEN_367 & ~_T_1492;
  assign stopEn134 = _GEN_367 & ~_T_1495;
  assign stopEn135 = _GEN_367 & ~_T_1499;
  assign stopEn136 = _GEN_379 & ~_T_1485;
  assign stopEn137 = _GEN_379 & ~_T_1488;
  assign stopEn138 = _GEN_379 & ~_T_1495;
  assign stopEn139 = _GEN_379 & ~_T_1805;
  assign stopEn140 = _GEN_387 & ~_T_1485;
  assign stopEn141 = _GEN_387 & ~_T_1488;
  assign stopEn142 = _GEN_387 & ~_T_1495;
  assign stopEn143 = _GEN_387 & ~_T_1805;
  assign stopEn144 = _GEN_395 & ~_T_1485;
  assign stopEn145 = _GEN_395 & ~_T_1488;
  assign stopEn146 = _GEN_395 & ~_T_1495;
  assign stopEn147 = _GEN_395 & ~_T_1805;
  assign stopEn148 = _T_1847 & ~_T_1850;
  assign stopEn149 = _T_1847 & ~_T_1854;
  assign stopEn150 = _T_1847 & ~_T_1858;
  assign stopEn151 = _T_1847 & ~_T_1862;
  assign stopEn152 = _T_1847 & ~_T_1866;
  assign stopEn153 = _T_1871 & ~_T_1874;
  assign stopEn154 = _T_1871 & ~_T_1878;
  assign stopEn155 = _T_1871 & ~_T_1882;
  assign stopEn156 = _T_1871 & ~_T_1886;
  assign stopEn157 = _T_1871 & ~_T_1890;
  assign stopEn158 = _T_1871 & ~_T_1894;
  assign stopEn159 = _T_1899 & ~_T_1902;
  assign stopEn160 = _T_1899 & ~_T_1906;
  assign stopEn161 = _T_1899 & ~_T_1910;
  assign stopEn162 = _T_1899 & ~_T_1914;
  assign stopEn163 = _T_1899 & ~_T_1918;
  assign stopEn164 = _T_1923 & ~_T_1926;
  assign stopEn165 = _T_1923 & ~_T_1930;
  assign stopEn166 = _T_1923 & ~_T_1934;
  assign stopEn167 = _T_1923 & ~_T_1938;
  assign stopEn168 = _T_1923 & ~_T_1942;
  assign stopEn169 = _T_1949 & ~_T_1955;
  assign stopEn170 = _T_1960 & ~_T_1974;
  assign stopEn171 = _GEN_403 & ~_T_1980;
  assign stopEn172 = _GEN_403 & ~_T_1984;
  assign stopEn173 = _GEN_408 & ~_T_1992;
  assign stopEn174 = _GEN_408 & ~_T_1996;
  assign stopEn175 = _T_2004 & ~_T_2008;
  assign stopEn176 = ~_T_2015;
  assign stopEn177 = ~_T_2024;
  assign stopEn178 = _T_2039 & ~_T_2044;
  assign stopEn179 = _T_2048 & ~_T_2060;
  assign stopEn180 = _GEN_415 & ~_T_2064;
  assign stopEn181 = _GEN_418 & ~_T_2068;
  assign stopEn182 = _T_2075 & ~_T_2079;
  assign stopEn183 = _T_2081 & ~_T_2084;
  assign stopEn184 = ~_T_2093;
  assign stopEn185 = _T_2104 & ~_T_2109;
  assign stopEn186 = _T_2111 & ~_T_2118;
//  assign plusarg_reader_metaAssert_wire = plusarg_reader_metaAssert;
//  assign plusarg_reader_1_metaAssert_wire = plusarg_reader_1_metaAssert;
  assign TLMonitor_23_or63 = stopEn0 | stopEn1;
  assign TLMonitor_23_or130 = stopEn3 | stopEn4;
  assign TLMonitor_23_or64 = stopEn2 | TLMonitor_23_or130;
  assign TLMonitor_23_or31 = TLMonitor_23_or63 | TLMonitor_23_or64;
  assign TLMonitor_23_or132 = stopEn6 | stopEn7;
  assign TLMonitor_23_or65 = stopEn5 | TLMonitor_23_or132;
  assign TLMonitor_23_or134 = stopEn9 | stopEn10;
  assign TLMonitor_23_or66 = stopEn8 | TLMonitor_23_or134;
  assign TLMonitor_23_or32 = TLMonitor_23_or65 | TLMonitor_23_or66;
  assign TLMonitor_23_or15 = TLMonitor_23_or31 | TLMonitor_23_or32;
  assign TLMonitor_23_or136 = stopEn12 | stopEn13;
  assign TLMonitor_23_or67 = stopEn11 | TLMonitor_23_or136;
  assign TLMonitor_23_or138 = stopEn15 | stopEn16;
  assign TLMonitor_23_or68 = stopEn14 | TLMonitor_23_or138;
  assign TLMonitor_23_or33 = TLMonitor_23_or67 | TLMonitor_23_or68;
  assign TLMonitor_23_or140 = stopEn18 | stopEn19;
  assign TLMonitor_23_or69 = stopEn17 | TLMonitor_23_or140;
  assign TLMonitor_23_or142 = stopEn21 | stopEn22;
  assign TLMonitor_23_or70 = stopEn20 | TLMonitor_23_or142;
  assign TLMonitor_23_or34 = TLMonitor_23_or69 | TLMonitor_23_or70;
  assign TLMonitor_23_or16 = TLMonitor_23_or33 | TLMonitor_23_or34;
  assign TLMonitor_23_or7 = TLMonitor_23_or15 | TLMonitor_23_or16;
  assign TLMonitor_23_or144 = stopEn24 | stopEn25;
  assign TLMonitor_23_or71 = stopEn23 | TLMonitor_23_or144;
  assign TLMonitor_23_or146 = stopEn27 | stopEn28;
  assign TLMonitor_23_or72 = stopEn26 | TLMonitor_23_or146;
  assign TLMonitor_23_or35 = TLMonitor_23_or71 | TLMonitor_23_or72;
  assign TLMonitor_23_or148 = stopEn30 | stopEn31;
  assign TLMonitor_23_or73 = stopEn29 | TLMonitor_23_or148;
  assign TLMonitor_23_or150 = stopEn33 | stopEn34;
  assign TLMonitor_23_or74 = stopEn32 | TLMonitor_23_or150;
  assign TLMonitor_23_or36 = TLMonitor_23_or73 | TLMonitor_23_or74;
  assign TLMonitor_23_or17 = TLMonitor_23_or35 | TLMonitor_23_or36;
  assign TLMonitor_23_or152 = stopEn36 | stopEn37;
  assign TLMonitor_23_or75 = stopEn35 | TLMonitor_23_or152;
  assign TLMonitor_23_or154 = stopEn39 | stopEn40;
  assign TLMonitor_23_or76 = stopEn38 | TLMonitor_23_or154;
  assign TLMonitor_23_or37 = TLMonitor_23_or75 | TLMonitor_23_or76;
  assign TLMonitor_23_or156 = stopEn42 | stopEn43;
  assign TLMonitor_23_or77 = stopEn41 | TLMonitor_23_or156;
  assign TLMonitor_23_or158 = stopEn45 | stopEn46;
  assign TLMonitor_23_or78 = stopEn44 | TLMonitor_23_or158;
  assign TLMonitor_23_or38 = TLMonitor_23_or77 | TLMonitor_23_or78;
  assign TLMonitor_23_or18 = TLMonitor_23_or37 | TLMonitor_23_or38;
  assign TLMonitor_23_or8 = TLMonitor_23_or17 | TLMonitor_23_or18;
  assign TLMonitor_23_or3 = TLMonitor_23_or7 | TLMonitor_23_or8;
  assign TLMonitor_23_or79 = stopEn47 | stopEn48;
  assign TLMonitor_23_or162 = stopEn50 | stopEn51;
  assign TLMonitor_23_or80 = stopEn49 | TLMonitor_23_or162;
  assign TLMonitor_23_or39 = TLMonitor_23_or79 | TLMonitor_23_or80;
  assign TLMonitor_23_or164 = stopEn53 | stopEn54;
  assign TLMonitor_23_or81 = stopEn52 | TLMonitor_23_or164;
  assign TLMonitor_23_or166 = stopEn56 | stopEn57;
  assign TLMonitor_23_or82 = stopEn55 | TLMonitor_23_or166;
  assign TLMonitor_23_or40 = TLMonitor_23_or81 | TLMonitor_23_or82;
  assign TLMonitor_23_or19 = TLMonitor_23_or39 | TLMonitor_23_or40;
  assign TLMonitor_23_or168 = stopEn59 | stopEn60;
  assign TLMonitor_23_or83 = stopEn58 | TLMonitor_23_or168;
  assign TLMonitor_23_or170 = stopEn62 | stopEn63;
  assign TLMonitor_23_or84 = stopEn61 | TLMonitor_23_or170;
  assign TLMonitor_23_or41 = TLMonitor_23_or83 | TLMonitor_23_or84;
  assign TLMonitor_23_or172 = stopEn65 | stopEn66;
  assign TLMonitor_23_or85 = stopEn64 | TLMonitor_23_or172;
  assign TLMonitor_23_or174 = stopEn68 | stopEn69;
  assign TLMonitor_23_or86 = stopEn67 | TLMonitor_23_or174;
  assign TLMonitor_23_or42 = TLMonitor_23_or85 | TLMonitor_23_or86;
  assign TLMonitor_23_or20 = TLMonitor_23_or41 | TLMonitor_23_or42;
  assign TLMonitor_23_or9 = TLMonitor_23_or19 | TLMonitor_23_or20;
  assign TLMonitor_23_or176 = stopEn71 | stopEn72;
  assign TLMonitor_23_or87 = stopEn70 | TLMonitor_23_or176;
  assign TLMonitor_23_or178 = stopEn74 | stopEn75;
  assign TLMonitor_23_or88 = stopEn73 | TLMonitor_23_or178;
  assign TLMonitor_23_or43 = TLMonitor_23_or87 | TLMonitor_23_or88;
  assign TLMonitor_23_or180 = stopEn77 | stopEn78;
  assign TLMonitor_23_or89 = stopEn76 | TLMonitor_23_or180;
  assign TLMonitor_23_or182 = stopEn80 | stopEn81;
  assign TLMonitor_23_or90 = stopEn79 | TLMonitor_23_or182;
  assign TLMonitor_23_or44 = TLMonitor_23_or89 | TLMonitor_23_or90;
  assign TLMonitor_23_or21 = TLMonitor_23_or43 | TLMonitor_23_or44;
  assign TLMonitor_23_or184 = stopEn83 | stopEn84;
  assign TLMonitor_23_or91 = stopEn82 | TLMonitor_23_or184;
  assign TLMonitor_23_or186 = stopEn86 | stopEn87;
  assign TLMonitor_23_or92 = stopEn85 | TLMonitor_23_or186;
  assign TLMonitor_23_or45 = TLMonitor_23_or91 | TLMonitor_23_or92;
  assign TLMonitor_23_or188 = stopEn89 | stopEn90;
  assign TLMonitor_23_or93 = stopEn88 | TLMonitor_23_or188;
  assign TLMonitor_23_or190 = stopEn92 | stopEn93;
  assign TLMonitor_23_or94 = stopEn91 | TLMonitor_23_or190;
  assign TLMonitor_23_or46 = TLMonitor_23_or93 | TLMonitor_23_or94;
  assign TLMonitor_23_or22 = TLMonitor_23_or45 | TLMonitor_23_or46;
  assign TLMonitor_23_or10 = TLMonitor_23_or21 | TLMonitor_23_or22;
  assign TLMonitor_23_or4 = TLMonitor_23_or9 | TLMonitor_23_or10;
  assign TLMonitor_23_or1 = TLMonitor_23_or3 | TLMonitor_23_or4;
  assign TLMonitor_23_or95 = stopEn94 | stopEn95;
  assign TLMonitor_23_or194 = stopEn97 | stopEn98;
  assign TLMonitor_23_or96 = stopEn96 | TLMonitor_23_or194;
  assign TLMonitor_23_or47 = TLMonitor_23_or95 | TLMonitor_23_or96;
  assign TLMonitor_23_or196 = stopEn100 | stopEn101;
  assign TLMonitor_23_or97 = stopEn99 | TLMonitor_23_or196;
  assign TLMonitor_23_or198 = stopEn103 | stopEn104;
  assign TLMonitor_23_or98 = stopEn102 | TLMonitor_23_or198;
  assign TLMonitor_23_or48 = TLMonitor_23_or97 | TLMonitor_23_or98;
  assign TLMonitor_23_or23 = TLMonitor_23_or47 | TLMonitor_23_or48;
  assign TLMonitor_23_or200 = stopEn106 | stopEn107;
  assign TLMonitor_23_or99 = stopEn105 | TLMonitor_23_or200;
  assign TLMonitor_23_or202 = stopEn109 | stopEn110;
  assign TLMonitor_23_or100 = stopEn108 | TLMonitor_23_or202;
  assign TLMonitor_23_or49 = TLMonitor_23_or99 | TLMonitor_23_or100;
  assign TLMonitor_23_or204 = stopEn112 | stopEn113;
  assign TLMonitor_23_or101 = stopEn111 | TLMonitor_23_or204;
  assign TLMonitor_23_or206 = stopEn115 | stopEn116;
  assign TLMonitor_23_or102 = stopEn114 | TLMonitor_23_or206;
  assign TLMonitor_23_or50 = TLMonitor_23_or101 | TLMonitor_23_or102;
  assign TLMonitor_23_or24 = TLMonitor_23_or49 | TLMonitor_23_or50;
  assign TLMonitor_23_or11 = TLMonitor_23_or23 | TLMonitor_23_or24;
  assign TLMonitor_23_or208 = stopEn118 | stopEn119;
  assign TLMonitor_23_or103 = stopEn117 | TLMonitor_23_or208;
  assign TLMonitor_23_or210 = stopEn121 | stopEn122;
  assign TLMonitor_23_or104 = stopEn120 | TLMonitor_23_or210;
  assign TLMonitor_23_or51 = TLMonitor_23_or103 | TLMonitor_23_or104;
  assign TLMonitor_23_or212 = stopEn124 | stopEn125;
  assign TLMonitor_23_or105 = stopEn123 | TLMonitor_23_or212;
  assign TLMonitor_23_or214 = stopEn127 | stopEn128;
  assign TLMonitor_23_or106 = stopEn126 | TLMonitor_23_or214;
  assign TLMonitor_23_or52 = TLMonitor_23_or105 | TLMonitor_23_or106;
  assign TLMonitor_23_or25 = TLMonitor_23_or51 | TLMonitor_23_or52;
  assign TLMonitor_23_or216 = stopEn130 | stopEn131;
  assign TLMonitor_23_or107 = stopEn129 | TLMonitor_23_or216;
  assign TLMonitor_23_or218 = stopEn133 | stopEn134;
  assign TLMonitor_23_or108 = stopEn132 | TLMonitor_23_or218;
  assign TLMonitor_23_or53 = TLMonitor_23_or107 | TLMonitor_23_or108;
  assign TLMonitor_23_or220 = stopEn136 | stopEn137;
  assign TLMonitor_23_or109 = stopEn135 | TLMonitor_23_or220;
  assign TLMonitor_23_or222 = stopEn139 | stopEn140;
  assign TLMonitor_23_or110 = stopEn138 | TLMonitor_23_or222;
  assign TLMonitor_23_or54 = TLMonitor_23_or109 | TLMonitor_23_or110;
  assign TLMonitor_23_or26 = TLMonitor_23_or53 | TLMonitor_23_or54;
  assign TLMonitor_23_or12 = TLMonitor_23_or25 | TLMonitor_23_or26;
  assign TLMonitor_23_or5 = TLMonitor_23_or11 | TLMonitor_23_or12;
  assign TLMonitor_23_or224 = stopEn142 | stopEn143;
  assign TLMonitor_23_or111 = stopEn141 | TLMonitor_23_or224;
  assign TLMonitor_23_or226 = stopEn145 | stopEn146;
  assign TLMonitor_23_or112 = stopEn144 | TLMonitor_23_or226;
  assign TLMonitor_23_or55 = TLMonitor_23_or111 | TLMonitor_23_or112;
  assign TLMonitor_23_or228 = stopEn148 | stopEn149;
  assign TLMonitor_23_or113 = stopEn147 | TLMonitor_23_or228;
  assign TLMonitor_23_or230 = stopEn151 | stopEn152;
  assign TLMonitor_23_or114 = stopEn150 | TLMonitor_23_or230;
  assign TLMonitor_23_or56 = TLMonitor_23_or113 | TLMonitor_23_or114;
  assign TLMonitor_23_or27 = TLMonitor_23_or55 | TLMonitor_23_or56;
  assign TLMonitor_23_or232 = stopEn154 | stopEn155;
  assign TLMonitor_23_or115 = stopEn153 | TLMonitor_23_or232;
  assign TLMonitor_23_or234 = stopEn157 | stopEn158;
  assign TLMonitor_23_or116 = stopEn156 | TLMonitor_23_or234;
  assign TLMonitor_23_or57 = TLMonitor_23_or115 | TLMonitor_23_or116;
  assign TLMonitor_23_or236 = stopEn160 | stopEn161;
  assign TLMonitor_23_or117 = stopEn159 | TLMonitor_23_or236;
  assign TLMonitor_23_or238 = stopEn163 | stopEn164;
  assign TLMonitor_23_or118 = stopEn162 | TLMonitor_23_or238;
  assign TLMonitor_23_or58 = TLMonitor_23_or117 | TLMonitor_23_or118;
  assign TLMonitor_23_or28 = TLMonitor_23_or57 | TLMonitor_23_or58;
  assign TLMonitor_23_or13 = TLMonitor_23_or27 | TLMonitor_23_or28;
  assign TLMonitor_23_or240 = stopEn166 | stopEn167;
  assign TLMonitor_23_or119 = stopEn165 | TLMonitor_23_or240;
  assign TLMonitor_23_or242 = stopEn169 | stopEn170;
  assign TLMonitor_23_or120 = stopEn168 | TLMonitor_23_or242;
  assign TLMonitor_23_or59 = TLMonitor_23_or119 | TLMonitor_23_or120;
  assign TLMonitor_23_or244 = stopEn172 | stopEn173;
  assign TLMonitor_23_or121 = stopEn171 | TLMonitor_23_or244;
  assign TLMonitor_23_or246 = stopEn175 | stopEn176;
  assign TLMonitor_23_or122 = stopEn174 | TLMonitor_23_or246;
  assign TLMonitor_23_or60 = TLMonitor_23_or121 | TLMonitor_23_or122;
  assign TLMonitor_23_or29 = TLMonitor_23_or59 | TLMonitor_23_or60;
  assign TLMonitor_23_or248 = stopEn178 | stopEn179;
  assign TLMonitor_23_or123 = stopEn177 | TLMonitor_23_or248;
  assign TLMonitor_23_or250 = stopEn181 | stopEn182;
  assign TLMonitor_23_or124 = stopEn180 | TLMonitor_23_or250;
  assign TLMonitor_23_or61 = TLMonitor_23_or123 | TLMonitor_23_or124;
  assign TLMonitor_23_or252 = stopEn184 | stopEn185;
  assign TLMonitor_23_or125 = stopEn183 | TLMonitor_23_or252;
  assign TLMonitor_23_or254 = plusarg_reader_metaAssert_wire | plusarg_reader_1_metaAssert_wire;
  assign TLMonitor_23_or126 = stopEn186 | TLMonitor_23_or254;
  assign TLMonitor_23_or62 = TLMonitor_23_or125 | TLMonitor_23_or126;
  assign TLMonitor_23_or30 = TLMonitor_23_or61 | TLMonitor_23_or62;
  assign TLMonitor_23_or14 = TLMonitor_23_or29 | TLMonitor_23_or30;
  assign TLMonitor_23_or6 = TLMonitor_23_or13 | TLMonitor_23_or14;
  assign TLMonitor_23_or2 = TLMonitor_23_or5 | TLMonitor_23_or6;
  assign TLMonitor_23_or0 = TLMonitor_23_or1 | TLMonitor_23_or2;
  assign metaAssert = TLMonitor_23_metaAssert;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  opcode = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  param = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  size = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  source = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  address = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  d_first_counter = _RAND_6[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  opcode_1 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  param_1 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  size_1 = _RAND_9[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  source_1 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  sink = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  denied = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  b_first_counter = _RAND_13[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  opcode_2 = _RAND_14[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  param_2 = _RAND_15[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  size_2 = _RAND_16[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  source_2 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  address_1 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  c_first_counter = _RAND_19[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  opcode_3 = _RAND_20[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  param_3 = _RAND_21[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  size_3 = _RAND_22[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  source_3 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  address_2 = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  inflight = _RAND_25[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  inflight_opcodes = _RAND_26[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  inflight_sizes = _RAND_27[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  a_first_counter_1 = _RAND_28[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  d_first_counter_1 = _RAND_29[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  watchdog = _RAND_30[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  inflight_1 = _RAND_31[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  inflight_sizes_1 = _RAND_32[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  c_first_counter_1 = _RAND_33[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  d_first_counter_2 = _RAND_34[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  watchdog_1 = _RAND_35[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  inflight_2 = _RAND_36[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  d_first_counter_3 = _RAND_37[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  TLMonitor_23_metaAssert = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      a_first_counter <= 9'h0;
    end else if (reset) begin
      a_first_counter <= 9'h0;
    end else if (_a_first_T) begin
      if (a_first) begin
        if (a_first_beats1_opdata) begin
          a_first_counter <= a_first_beats1_decode;
        end else begin
          a_first_counter <= 9'h0;
        end
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (metaReset) begin
      opcode <= 3'h0;
    end else if (_T_1869) begin
      opcode <= io_in_a_bits_opcode;
    end
    if (metaReset) begin
      param <= 3'h0;
    end else if (_T_1869) begin
      param <= io_in_a_bits_param;
    end
    if (metaReset) begin
      size <= 4'h0;
    end else if (_T_1869) begin
      size <= io_in_a_bits_size;
    end
    if (metaReset) begin
      source <= 1'h0;
    end else if (_T_1869) begin
      source <= io_in_a_bits_source;
    end
    if (metaReset) begin
      address <= 32'h0;
    end else if (_T_1869) begin
      address <= io_in_a_bits_address;
    end
    if (metaReset) begin
      d_first_counter <= 9'h0;
    end else if (reset) begin
      d_first_counter <= 9'h0;
    end else if (_d_first_T) begin
      if (d_first) begin
        if (d_first_beats1_opdata) begin
          d_first_counter <= d_first_beats1_decode;
        end else begin
          d_first_counter <= 9'h0;
        end
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    if (metaReset) begin
      opcode_1 <= 3'h0;
    end else if (_T_1897) begin
      opcode_1 <= io_in_d_bits_opcode;
    end
    if (metaReset) begin
      param_1 <= 2'h0;
    end else if (_T_1897) begin
      param_1 <= io_in_d_bits_param;
    end
    if (metaReset) begin
      size_1 <= 4'h0;
    end else if (_T_1897) begin
      size_1 <= io_in_d_bits_size;
    end
    if (metaReset) begin
      source_1 <= 1'h0;
    end else if (_T_1897) begin
      source_1 <= io_in_d_bits_source;
    end
    if (metaReset) begin
      sink <= 2'h0;
    end else if (_T_1897) begin
      sink <= io_in_d_bits_sink;
    end
    if (metaReset) begin
      denied <= 1'h0;
    end else if (_T_1897) begin
      denied <= io_in_d_bits_denied;
    end
    if (metaReset) begin
      b_first_counter <= 9'h0;
    end else if (reset) begin
      b_first_counter <= 9'h0;
    end else if (b_first_done) begin
      if (b_first) begin
        b_first_counter <= 9'h0;
      end else begin
        b_first_counter <= b_first_counter1;
      end
    end
    if (metaReset) begin
      opcode_2 <= 3'h0;
    end else if (_T_1921) begin
      opcode_2 <= io_in_b_bits_opcode;
    end
    if (metaReset) begin
      param_2 <= 2'h0;
    end else if (_T_1921) begin
      param_2 <= io_in_b_bits_param;
    end
    if (metaReset) begin
      size_2 <= 4'h0;
    end else if (_T_1921) begin
      size_2 <= io_in_b_bits_size;
    end
    if (metaReset) begin
      source_2 <= 1'h0;
    end else if (_T_1921) begin
      source_2 <= io_in_b_bits_source;
    end
    if (metaReset) begin
      address_1 <= 32'h0;
    end else if (_T_1921) begin
      address_1 <= io_in_b_bits_address;
    end
    if (metaReset) begin
      c_first_counter <= 9'h0;
    end else if (reset) begin
      c_first_counter <= 9'h0;
    end else if (_c_first_T) begin
      if (c_first) begin
        if (c_first_beats1_opdata) begin
          c_first_counter <= c_first_beats1_decode;
        end else begin
          c_first_counter <= 9'h0;
        end
      end else begin
        c_first_counter <= c_first_counter1;
      end
    end
    if (metaReset) begin
      opcode_3 <= 3'h0;
    end else if (_T_1945) begin
      opcode_3 <= io_in_c_bits_opcode;
    end
    if (metaReset) begin
      param_3 <= 3'h0;
    end else if (_T_1945) begin
      param_3 <= io_in_c_bits_param;
    end
    if (metaReset) begin
      size_3 <= 4'h0;
    end else if (_T_1945) begin
      size_3 <= io_in_c_bits_size;
    end
    if (metaReset) begin
      source_3 <= 1'h0;
    end else if (_T_1945) begin
      source_3 <= io_in_c_bits_source;
    end
    if (metaReset) begin
      address_2 <= 32'h0;
    end else if (_T_1945) begin
      address_2 <= io_in_c_bits_address;
    end
    if (metaReset) begin
      inflight <= 2'h0;
    end else if (reset) begin
      inflight <= 2'h0;
    end else begin
      inflight <= _inflight_T_2;
    end
    if (metaReset) begin
      inflight_opcodes <= 8'h0;
    end else if (reset) begin
      inflight_opcodes <= 8'h0;
    end else begin
      inflight_opcodes <= _inflight_opcodes_T_2;
    end
    if (metaReset) begin
      inflight_sizes <= 16'h0;
    end else if (reset) begin
      inflight_sizes <= 16'h0;
    end else begin
      inflight_sizes <= _inflight_sizes_T_2;
    end
    if (metaReset) begin
      a_first_counter_1 <= 9'h0;
    end else if (reset) begin
      a_first_counter_1 <= 9'h0;
    end else if (_a_first_T) begin
      if (a_first_1) begin
        if (a_first_beats1_opdata) begin
          a_first_counter_1 <= a_first_beats1_decode;
        end else begin
          a_first_counter_1 <= 9'h0;
        end
      end else begin
        a_first_counter_1 <= a_first_counter1_1;
      end
    end
    if (metaReset) begin
      d_first_counter_1 <= 9'h0;
    end else if (reset) begin
      d_first_counter_1 <= 9'h0;
    end else if (_d_first_T) begin
      if (d_first_1) begin
        if (d_first_beats1_opdata) begin
          d_first_counter_1 <= d_first_beats1_decode;
        end else begin
          d_first_counter_1 <= 9'h0;
        end
      end else begin
        d_first_counter_1 <= d_first_counter1_1;
      end
    end
    if (metaReset) begin
      watchdog <= 32'h0;
    end else if (reset) begin
      watchdog <= 32'h0;
    end else if (_T_2028) begin
      watchdog <= 32'h0;
    end else begin
      watchdog <= _watchdog_T_1;
    end
    if (metaReset) begin
      inflight_1 <= 2'h0;
    end else if (reset) begin
      inflight_1 <= 2'h0;
    end else begin
      inflight_1 <= _inflight_T_5;
    end
    if (metaReset) begin
      inflight_sizes_1 <= 16'h0;
    end else if (reset) begin
      inflight_sizes_1 <= 16'h0;
    end else begin
      inflight_sizes_1 <= _inflight_sizes_T_5;
    end
    if (metaReset) begin
      c_first_counter_1 <= 9'h0;
    end else if (reset) begin
      c_first_counter_1 <= 9'h0;
    end else if (_c_first_T) begin
      if (c_first_1) begin
        if (c_first_beats1_opdata) begin
          c_first_counter_1 <= c_first_beats1_decode;
        end else begin
          c_first_counter_1 <= 9'h0;
        end
      end else begin
        c_first_counter_1 <= c_first_counter1_1;
      end
    end
    if (metaReset) begin
      d_first_counter_2 <= 9'h0;
    end else if (reset) begin
      d_first_counter_2 <= 9'h0;
    end else if (_d_first_T) begin
      if (d_first_2) begin
        if (d_first_beats1_opdata) begin
          d_first_counter_2 <= d_first_beats1_decode;
        end else begin
          d_first_counter_2 <= 9'h0;
        end
      end else begin
        d_first_counter_2 <= d_first_counter1_2;
      end
    end
    if (metaReset) begin
      watchdog_1 <= 32'h0;
    end else if (reset) begin
      watchdog_1 <= 32'h0;
    end else if (_T_2097) begin
      watchdog_1 <= 32'h0;
    end else begin
      watchdog_1 <= _watchdog_T_3;
    end
    if (metaReset) begin
      inflight_2 <= 4'h0;
    end else if (reset) begin
      inflight_2 <= 4'h0;
    end else begin
      inflight_2 <= _inflight_T_8;
    end
    if (metaReset) begin
      d_first_counter_3 <= 9'h0;
    end else if (reset) begin
      d_first_counter_3 <= 9'h0;
    end else if (_d_first_T) begin
      if (d_first_3) begin
        if (d_first_beats1_opdata) begin
          d_first_counter_3 <= d_first_beats1_decode;
        end else begin
          d_first_counter_3 <= 9'h0;
        end
      end else begin
        d_first_counter_3 <= d_first_counter1_3;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_111 & ~_T_84) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_111 & ~_T_84) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_111 & ~_T_141) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_111 & ~_T_141) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_111 & ~_T_144) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_111 & ~_T_144) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_111 & ~_T_148) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_111 & ~_T_148) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_111 & ~_T_151) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_111 & ~_T_151) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_111 & ~_T_155) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_111 & ~_T_155) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_111 & ~_T_160) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_111 & ~_T_160) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & ~_T_84) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & ~_T_84) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & ~_T_141) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & ~_T_141) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & ~_T_144) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & ~_T_144) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & ~_T_148) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & ~_T_148) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & ~_T_151) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & ~_T_151) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & ~_T_155) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & ~_T_155) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & ~_T_301) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & ~_T_301) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_125 & ~_T_160) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_125 & ~_T_160) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & ~_T_322) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & ~_T_322) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & ~_T_377) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & ~_T_377) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & ~_T_144) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & ~_T_144) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & ~_T_151) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & ~_T_151) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & ~_T_387) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & ~_T_387) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & ~_T_391) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get contains invalid mask (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & ~_T_391) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_153 & ~_T_467) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_153 & ~_T_467) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_153 & ~_T_144) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_153 & ~_T_144) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_153 & ~_T_151) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_153 & ~_T_151) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_153 & ~_T_387) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_153 & ~_T_387) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_153 & ~_T_391) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull contains invalid mask (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_153 & ~_T_391) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_163 & ~_T_467) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_163 & ~_T_467) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_163 & ~_T_144) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_163 & ~_T_144) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_163 & ~_T_151) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_163 & ~_T_151) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_163 & ~_T_387) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_163 & ~_T_387) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_163 & ~_T_569) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial contains invalid mask (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_163 & ~_T_569) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_173 & ~_T_631) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_173 & ~_T_631) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_173 & ~_T_144) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_173 & ~_T_144) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_173 & ~_T_151) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_173 & ~_T_151) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_173 & ~_T_641) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_173 & ~_T_641) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_173 & ~_T_391) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_173 & ~_T_391) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_183 & ~_T_631) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_183 & ~_T_631) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_183 & ~_T_144) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_183 & ~_T_144) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_183 & ~_T_151) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_183 & ~_T_151) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_183 & ~_T_717) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid opcode param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_183 & ~_T_717) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_183 & ~_T_391) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical contains invalid mask (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_183 & ~_T_391) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_193 & ~_T_783) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_193 & ~_T_783) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_193 & ~_T_144) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_193 & ~_T_144) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_193 & ~_T_151) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_193 & ~_T_151) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_193 & ~_T_793) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint carries invalid opcode param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_193 & ~_T_793) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_193 & ~_T_391) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint contains invalid mask (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_193 & ~_T_391) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & ~_T_805) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel has invalid opcode (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & ~_T_805) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_203 & ~_T_809) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & ~_T_809) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_203 & ~_T_813) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & ~_T_813) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_203 & ~_T_817) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & ~_T_817) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_203 & ~_T_821) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is corrupt (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & ~_T_821) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_203 & ~_T_825) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is denied (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & ~_T_825) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_213 & ~_T_809) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_213 & ~_T_809) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_213 & ~_T_813) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant smaller than a beat (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_213 & ~_T_813) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_213 & ~_T_840) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid cap param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_213 & ~_T_840) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_213 & ~_T_844) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries toN param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_213 & ~_T_844) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_213 & ~_T_821) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is corrupt (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_213 & ~_T_821) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & ~_T_809) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & ~_T_809) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & ~_T_813) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData smaller than a beat (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & ~_T_813) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & ~_T_840) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid cap param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & ~_T_840) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & ~_T_844) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries toN param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & ~_T_844) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & ~_T_877) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & ~_T_877) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & ~_T_809) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & ~_T_809) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & ~_T_817) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & ~_T_817) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & ~_T_821) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is corrupt (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & ~_T_821) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_239 & ~_T_809) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_239 & ~_T_809) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_239 & ~_T_817) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_239 & ~_T_817) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_239 & ~_T_877) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_239 & ~_T_877) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_245 & ~_T_809) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_245 & ~_T_809) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_245 & ~_T_817) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_245 & ~_T_817) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_245 & ~_T_821) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is corrupt (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_245 & ~_T_821) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_b_valid & ~_T_938) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel has invalid opcode (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_b_valid & ~_T_938) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_251 & ~_T_1016) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Probe type which is unexpected using diplomatic parameters (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_251 & ~_T_1016) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_251 & ~_T_1019) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries unmanaged address (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_251 & ~_T_1019) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_251 & ~_T_1022) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries source that is not first source (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_251 & ~_T_1022) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_251 & ~_T_1025) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_251 & ~_T_1025) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_251 & ~_T_1029) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries invalid cap param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_251 & ~_T_1029) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_251 & ~_T_1033) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe contains invalid mask (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_251 & ~_T_1033) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_251 & ~_T_1037) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe is corrupt (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_251 & ~_T_1037) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_265 & ~reset) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Get type which is unexpected using diplomatic parameters (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_265 & ~reset) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_265 & ~_T_1019) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries unmanaged address (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_265 & ~_T_1019) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_265 & ~_T_1022) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries source that is not first source (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_265 & ~_T_1022) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_265 & ~_T_1025) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_265 & ~_T_1025) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_265 & ~_T_1102) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries invalid param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_265 & ~_T_1102) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_265 & ~_T_1033) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get contains invalid mask (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_265 & ~_T_1033) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_265 & ~_T_1037) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get is corrupt (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_265 & ~_T_1037) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_279 & ~reset) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries PutFull type which is unexpected using diplomatic parameters (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_279 & ~reset) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_279 & ~_T_1019) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries unmanaged address (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_279 & ~_T_1019) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_279 & ~_T_1022) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries source that is not first source (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_279 & ~_T_1022) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_279 & ~_T_1025) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_279 & ~_T_1025) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_279 & ~_T_1102) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries invalid param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_279 & ~_T_1102) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_279 & ~_T_1033) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull contains invalid mask (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_279 & ~_T_1033) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_291 & ~reset) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_291 & ~reset) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_291 & ~_T_1019) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries unmanaged address (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_291 & ~_T_1019) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_291 & ~_T_1022) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries source that is not first source (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_291 & ~_T_1022) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_291 & ~_T_1025) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_291 & ~_T_1025) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_291 & ~_T_1102) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries invalid param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_291 & ~_T_1102) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_291 & ~_T_1250) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial contains invalid mask (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_291 & ~_T_1250) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_303 & ~reset) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Arithmetic type unsupported by master (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_303 & ~reset) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_303 & ~_T_1019) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic carries unmanaged address (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_303 & ~_T_1019) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_303 & ~_T_1022) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic carries source that is not first source (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_303 & ~_T_1022) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_303 & ~_T_1025) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_303 & ~_T_1025) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_303 & ~_T_1033) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic contains invalid mask (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_303 & ~_T_1033) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_313 & ~reset) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Logical type unsupported by client (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_313 & ~reset) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_313 & ~_T_1019) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical carries unmanaged address (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_313 & ~_T_1019) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_313 & ~_T_1022) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical carries source that is not first source (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_313 & ~_T_1022) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_313 & ~_T_1025) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_313 & ~_T_1025) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_313 & ~_T_1033) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical contains invalid mask (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_313 & ~_T_1033) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_323 & ~reset) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Hint type unsupported by client (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_323 & ~reset) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_323 & ~_T_1019) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint carries unmanaged address (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_323 & ~_T_1019) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_323 & ~_T_1022) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint carries source that is not first source (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_323 & ~_T_1022) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_323 & ~_T_1025) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_323 & ~_T_1025) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_323 & ~_T_1033) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint contains invalid mask (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_323 & ~_T_1033) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_323 & ~_T_1037) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint is corrupt (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_323 & ~_T_1037) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_335 & ~_T_1485) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries unmanaged address (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_335 & ~_T_1485) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_335 & ~_T_1488) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_335 & ~_T_1488) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_335 & ~_T_1492) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck smaller than a beat (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_335 & ~_T_1492) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_335 & ~_T_1495) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_335 & ~_T_1495) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_335 & ~_T_1499) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries invalid report param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_335 & ~_T_1499) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_345 & ~_T_1485) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries unmanaged address (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_345 & ~_T_1485) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_345 & ~_T_1488) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_345 & ~_T_1488) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_345 & ~_T_1492) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData smaller than a beat (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_345 & ~_T_1492) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_345 & ~_T_1495) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_345 & ~_T_1495) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_345 & ~_T_1499) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries invalid report param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_345 & ~_T_1499) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_355 & ~_T_1583) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release type unsupported by manager (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_355 & ~_T_1583) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_355 & ~_T_1640) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_355 & ~_T_1640) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_355 & ~_T_1488) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_355 & ~_T_1488) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_355 & ~_T_1492) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release smaller than a beat (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_355 & ~_T_1492) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_355 & ~_T_1495) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_355 & ~_T_1495) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_355 & ~_T_1499) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release carries invalid report param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_355 & ~_T_1499) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_367 & ~_T_1583) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries ReleaseData type unsupported by manager (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_367 & ~_T_1583) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_367 & ~_T_1640) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_367 & ~_T_1640) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_367 & ~_T_1488) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_367 & ~_T_1488) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_367 & ~_T_1492) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData smaller than a beat (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_367 & ~_T_1492) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_367 & ~_T_1495) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_367 & ~_T_1495) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_367 & ~_T_1499) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData carries invalid report param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_367 & ~_T_1499) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_379 & ~_T_1485) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries unmanaged address (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_379 & ~_T_1485) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_379 & ~_T_1488) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_379 & ~_T_1488) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_379 & ~_T_1495) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_379 & ~_T_1495) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_379 & ~_T_1805) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries invalid param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_379 & ~_T_1805) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_387 & ~_T_1485) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries unmanaged address (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_387 & ~_T_1485) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_387 & ~_T_1488) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_387 & ~_T_1488) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_387 & ~_T_1495) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_387 & ~_T_1495) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_387 & ~_T_1805) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries invalid param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_387 & ~_T_1805) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_395 & ~_T_1485) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries unmanaged address (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_395 & ~_T_1485) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_395 & ~_T_1488) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_395 & ~_T_1488) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_395 & ~_T_1495) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_395 & ~_T_1495) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_395 & ~_T_1805) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries invalid param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_395 & ~_T_1805) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1847 & ~_T_1850) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel opcode changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1847 & ~_T_1850) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1847 & ~_T_1854) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel param changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1847 & ~_T_1854) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1847 & ~_T_1858) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel size changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1847 & ~_T_1858) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1847 & ~_T_1862) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel source changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1847 & ~_T_1862) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1847 & ~_T_1866) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel address changed with multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1847 & ~_T_1866) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1871 & ~_T_1874) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel opcode changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1871 & ~_T_1874) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1871 & ~_T_1878) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel param changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1871 & ~_T_1878) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1871 & ~_T_1882) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel size changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1871 & ~_T_1882) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1871 & ~_T_1886) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel source changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1871 & ~_T_1886) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1871 & ~_T_1890) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel sink changed with multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1871 & ~_T_1890) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1871 & ~_T_1894) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel denied changed with multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1871 & ~_T_1894) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1899 & ~_T_1902) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel opcode changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1899 & ~_T_1902) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1899 & ~_T_1906) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel param changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1899 & ~_T_1906) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1899 & ~_T_1910) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel size changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1899 & ~_T_1910) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1899 & ~_T_1914) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel source changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1899 & ~_T_1914) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1899 & ~_T_1918) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel addresss changed with multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1899 & ~_T_1918) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1923 & ~_T_1926) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel opcode changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1923 & ~_T_1926) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1923 & ~_T_1930) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel param changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1923 & ~_T_1930) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1923 & ~_T_1934) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel size changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1923 & ~_T_1934) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1923 & ~_T_1938) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel source changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1923 & ~_T_1938) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1923 & ~_T_1942) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel address changed with multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1923 & ~_T_1942) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1949 & ~_T_1955) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel re-used a source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1949 & ~_T_1955) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1960 & ~_T_1974) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel acknowledged for nothing inflight (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1960 & ~_T_1974) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_403 & ~_T_1980) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel contains improper opcode response (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_403 & ~_T_1980) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_403 & ~_T_1984) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel contains improper response size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_403 & ~_T_1984) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_408 & ~_T_1992) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel contains improper opcode response (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_408 & ~_T_1992) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_408 & ~_T_1996) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel contains improper response size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_408 & ~_T_1996) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2004 & ~_T_2008) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2004 & ~_T_2008) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_2015) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' and 'D' concurrent, despite minlatency 3 (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_2015) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_2024) begin
          $fwrite(32'h80000002,"Assertion failed: TileLink timeout expired (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_2024) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2039 & ~_T_2044) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel re-used a source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2039 & ~_T_2044) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2048 & ~_T_2060) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel acknowledged for nothing inflight (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2048 & ~_T_2060) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_415 & ~_T_2064) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel contains improper response size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_415 & ~_T_2064) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_418 & ~_T_2068) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel contains improper response size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_418 & ~_T_2068) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2075 & ~_T_2079) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2075 & ~_T_2079) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2081 & ~_T_2084) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' and 'D' concurrent, despite minlatency 3 (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2081 & ~_T_2084) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_2093) begin
          $fwrite(32'h80000002,"Assertion failed: TileLink timeout expired (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_2093) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2104 & ~_T_2109) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel re-used a sink ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2104 & ~_T_2109) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2111 & ~_T_2118) begin
          $fwrite(32'h80000002,"Assertion failed: 'E' channel acknowledged for nothing inflight (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2111 & ~_T_2118) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    if (metaReset) begin
      TLMonitor_23_metaAssert <= 1'h0;
    end else begin
      TLMonitor_23_metaAssert <= TLMonitor_23_metaAssert | TLMonitor_23_or0;
    end
  end
endmodule
module TLMonitor_24(
  input         clock,
  input         reset,
  input         io_in_a_ready,
  input         io_in_a_valid,
  input  [31:0] io_in_a_bits_address,
  input         io_in_d_valid,
  input  [2:0]  io_in_d_bits_opcode,
  input  [1:0]  io_in_d_bits_param,
  input  [3:0]  io_in_d_bits_size,
  input  [1:0]  io_in_d_bits_sink,
  input         io_in_d_bits_denied,
  input         io_in_d_bits_corrupt,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11]
  wire [31:0] plusarg_reader_1_out; // @[PlusArg.scala 80:11]
  wire [31:0] _is_aligned_T; // @[Edges.scala 20:16]
  wire  is_aligned; // @[Edges.scala 20:24]
  wire [32:0] _T_7; // @[Parameters.scala 137:49]
  wire [32:0] _T_26; // @[Parameters.scala 137:52]
  wire  _T_27; // @[Parameters.scala 137:67]
  wire [31:0] _T_28; // @[Parameters.scala 137:31]
  wire [32:0] _T_29; // @[Parameters.scala 137:49]
  wire [32:0] _T_31; // @[Parameters.scala 137:52]
  wire  _T_32; // @[Parameters.scala 137:67]
  wire [31:0] _T_33; // @[Parameters.scala 137:31]
  wire [32:0] _T_34; // @[Parameters.scala 137:49]
  wire [32:0] _T_36; // @[Parameters.scala 137:52]
  wire  _T_37; // @[Parameters.scala 137:67]
  wire [31:0] _T_38; // @[Parameters.scala 137:31]
  wire [32:0] _T_39; // @[Parameters.scala 137:49]
  wire [32:0] _T_41; // @[Parameters.scala 137:52]
  wire  _T_42; // @[Parameters.scala 137:67]
  wire [31:0] _T_43; // @[Parameters.scala 137:31]
  wire [32:0] _T_44; // @[Parameters.scala 137:49]
  wire [32:0] _T_46; // @[Parameters.scala 137:52]
  wire  _T_47; // @[Parameters.scala 137:67]
  wire [31:0] _T_48; // @[Parameters.scala 137:31]
  wire [32:0] _T_49; // @[Parameters.scala 137:49]
  wire [32:0] _T_51; // @[Parameters.scala 137:52]
  wire  _T_52; // @[Parameters.scala 137:67]
  wire [31:0] _T_63; // @[Parameters.scala 137:31]
  wire [32:0] _T_64; // @[Parameters.scala 137:49]
  wire [32:0] _T_66; // @[Parameters.scala 137:52]
  wire  _T_67; // @[Parameters.scala 137:67]
  wire  _T_134; // @[Monitor.scala 42:11]
  wire  _T_341; // @[Parameters.scala 671:42]
  wire  _T_342; // @[Parameters.scala 671:42]
  wire  _T_343; // @[Parameters.scala 671:42]
  wire  _T_344; // @[Parameters.scala 671:42]
  wire  _T_345; // @[Parameters.scala 671:42]
  wire  _T_348; // @[Parameters.scala 672:30]
  wire  _T_350; // @[Monitor.scala 42:11]
  wire  _T_766; // @[Bundles.scala 42:24]
  wire  _T_768; // @[Monitor.scala 49:11]
  wire  _T_770; // @[Monitor.scala 310:25]
  wire  _T_774; // @[Monitor.scala 312:27]
  wire  _T_776; // @[Monitor.scala 49:11]
  wire  _T_778; // @[Monitor.scala 313:28]
  wire  _T_780; // @[Monitor.scala 49:11]
  wire  _T_784; // @[Monitor.scala 49:11]
  wire  _T_788; // @[Monitor.scala 49:11]
  wire  _T_790; // @[Monitor.scala 318:25]
  wire  _T_801; // @[Bundles.scala 102:26]
  wire  _T_803; // @[Monitor.scala 49:11]
  wire  _T_805; // @[Monitor.scala 323:28]
  wire  _T_807; // @[Monitor.scala 49:11]
  wire  _T_818; // @[Monitor.scala 328:25]
  wire  _T_838; // @[Monitor.scala 334:30]
  wire  _T_840; // @[Monitor.scala 49:11]
  wire  _T_847; // @[Monitor.scala 338:25]
  wire  _T_864; // @[Monitor.scala 346:25]
  wire  _T_882; // @[Monitor.scala 354:25]
  wire  a_first_done; // @[Decoupled.scala 40:37]
  reg [8:0] a_first_counter; // @[Edges.scala 228:27]
  reg [31:0] _RAND_0;
  wire [8:0] a_first_counter1; // @[Edges.scala 229:28]
  wire  a_first; // @[Edges.scala 230:25]
  reg [31:0] address; // @[Monitor.scala 388:22]
  reg [31:0] _RAND_1;
  wire  _T_912; // @[Monitor.scala 389:19]
  wire  _T_929; // @[Monitor.scala 394:32]
  wire  _T_931; // @[Monitor.scala 42:11]
  wire  _T_934; // @[Monitor.scala 396:20]
  wire [26:0] _d_first_beats1_decode_T_1; // @[package.scala 234:77]
  wire [8:0] d_first_beats1_decode; // @[Edges.scala 219:59]
  wire  d_first_beats1_opdata; // @[Edges.scala 105:36]
  reg [8:0] d_first_counter; // @[Edges.scala 228:27]
  reg [31:0] _RAND_2;
  wire [8:0] d_first_counter1; // @[Edges.scala 229:28]
  wire  d_first; // @[Edges.scala 230:25]
  reg [2:0] opcode_1; // @[Monitor.scala 535:22]
  reg [31:0] _RAND_3;
  reg [1:0] param_1; // @[Monitor.scala 536:22]
  reg [31:0] _RAND_4;
  reg [3:0] size_1; // @[Monitor.scala 537:22]
  reg [31:0] _RAND_5;
  reg [1:0] sink; // @[Monitor.scala 539:22]
  reg [31:0] _RAND_6;
  reg  denied; // @[Monitor.scala 540:22]
  reg [31:0] _RAND_7;
  wire  _T_936; // @[Monitor.scala 541:19]
  wire  _T_937; // @[Monitor.scala 542:29]
  wire  _T_939; // @[Monitor.scala 49:11]
  wire  _T_941; // @[Monitor.scala 543:29]
  wire  _T_943; // @[Monitor.scala 49:11]
  wire  _T_945; // @[Monitor.scala 544:29]
  wire  _T_947; // @[Monitor.scala 49:11]
  wire  _T_953; // @[Monitor.scala 546:29]
  wire  _T_955; // @[Monitor.scala 49:11]
  wire  _T_957; // @[Monitor.scala 547:29]
  wire  _T_959; // @[Monitor.scala 49:11]
  wire  _T_962; // @[Monitor.scala 549:20]
  reg  inflight; // @[Monitor.scala 611:27]
  reg [31:0] _RAND_8;
  reg [3:0] inflight_opcodes; // @[Monitor.scala 613:35]
  reg [31:0] _RAND_9;
  reg [7:0] inflight_sizes; // @[Monitor.scala 615:33]
  reg [31:0] _RAND_10;
  reg [8:0] a_first_counter_1; // @[Edges.scala 228:27]
  reg [31:0] _RAND_11;
  wire [8:0] a_first_counter1_1; // @[Edges.scala 229:28]
  wire  a_first_1; // @[Edges.scala 230:25]
  reg [8:0] d_first_counter_1; // @[Edges.scala 228:27]
  reg [31:0] _RAND_12;
  wire [8:0] d_first_counter1_1; // @[Edges.scala 229:28]
  wire  d_first_1; // @[Edges.scala 230:25]
  wire [15:0] _a_opcode_lookup_T_5; // @[Monitor.scala 609:57]
  wire [15:0] _GEN_71; // @[Monitor.scala 634:97]
  wire [15:0] _a_opcode_lookup_T_6; // @[Monitor.scala 634:97]
  wire [15:0] _a_opcode_lookup_T_7; // @[Monitor.scala 634:152]
  wire [15:0] _a_size_lookup_T_5; // @[Monitor.scala 609:57]
  wire [15:0] _GEN_73; // @[Monitor.scala 638:91]
  wire [15:0] _a_size_lookup_T_6; // @[Monitor.scala 638:91]
  wire [15:0] _a_size_lookup_T_7; // @[Monitor.scala 638:144]
  wire  _T_963; // @[Monitor.scala 648:26]
  wire [1:0] _GEN_15; // @[Monitor.scala 648:71]
  wire  _T_966; // @[Monitor.scala 652:27]
  wire [3:0] a_opcodes_set_interm; // @[Monitor.scala 652:72]
  wire [18:0] _a_opcodes_set_T_1; // @[Monitor.scala 656:54]
  wire [4:0] a_sizes_set_interm; // @[Monitor.scala 652:72]
  wire [19:0] _a_sizes_set_T_1; // @[Monitor.scala 657:52]
  wire  _T_972; // @[Monitor.scala 42:11]
  wire [1:0] _GEN_16; // @[Monitor.scala 652:72]
  wire [18:0] _GEN_19; // @[Monitor.scala 652:72]
  wire [19:0] _GEN_20; // @[Monitor.scala 652:72]
  wire  _T_974; // @[Monitor.scala 671:26]
  wire  _T_977; // @[Monitor.scala 671:71]
  wire [1:0] _GEN_21; // @[Monitor.scala 671:90]
  wire [30:0] _d_opcodes_clr_T_5; // @[Monitor.scala 677:76]
  wire [30:0] _d_sizes_clr_T_5; // @[Monitor.scala 678:74]
  wire [30:0] _GEN_23; // @[Monitor.scala 675:91]
  wire [30:0] _GEN_24; // @[Monitor.scala 675:91]
  wire  _T_989; // @[Monitor.scala 682:49]
  wire  _T_991; // @[Monitor.scala 49:11]
  wire  _T_995; // @[Monitor.scala 685:77]
  wire  _T_997; // @[Monitor.scala 49:11]
  wire  _T_999; // @[Monitor.scala 687:36]
  wire  _T_1001; // @[Monitor.scala 49:11]
  wire [3:0] a_opcode_lookup; // @[Monitor.scala 634:21]
  wire [2:0] _GEN_43; // @[Monitor.scala 689:38]
  wire [2:0] _GEN_44; // @[Monitor.scala 689:38]
  wire [2:0] _GEN_45; // @[Monitor.scala 689:38]
  wire [2:0] _GEN_46; // @[Monitor.scala 689:38]
  wire [2:0] _GEN_47; // @[Monitor.scala 689:38]
  wire [2:0] _GEN_48; // @[Monitor.scala 689:38]
  wire  _T_1004; // @[Monitor.scala 689:38]
  wire [2:0] _GEN_55; // @[Monitor.scala 690:38]
  wire [2:0] _GEN_56; // @[Monitor.scala 690:38]
  wire  _T_1006; // @[Monitor.scala 690:38]
  wire  _T_1007; // @[Monitor.scala 689:72]
  wire  _T_1009; // @[Monitor.scala 49:11]
  wire [7:0] a_size_lookup; // @[Monitor.scala 638:19]
  wire [7:0] _GEN_75; // @[Monitor.scala 691:36]
  wire  _T_1011; // @[Monitor.scala 691:36]
  wire  _T_1013; // @[Monitor.scala 49:11]
  wire  _T_1016; // @[Monitor.scala 694:36]
  wire  _T_1017; // @[Monitor.scala 694:47]
  wire  _T_1021; // @[Monitor.scala 694:116]
  wire  _T_1025; // @[Monitor.scala 49:11]
  wire  a_set_wo_ready; // @[Monitor.scala 649:22]
  wire  d_clr_wo_ready; // @[Monitor.scala 672:22]
  wire  _T_1027; // @[Monitor.scala 699:29]
  wire  _T_1028; // @[Monitor.scala 699:67]
  wire  _T_1030; // @[Monitor.scala 699:48]
  wire  _T_1032; // @[Monitor.scala 49:11]
  wire  a_set; // @[Monitor.scala 653:28]
  wire  _inflight_T; // @[Monitor.scala 702:27]
  wire  _inflight_T_2; // @[Monitor.scala 702:36]
  wire [3:0] a_opcodes_set; // @[Monitor.scala 656:28]
  wire [3:0] _inflight_opcodes_T; // @[Monitor.scala 703:43]
  wire [3:0] d_opcodes_clr; // @[Monitor.scala 677:21]
  wire [3:0] _inflight_opcodes_T_2; // @[Monitor.scala 703:60]
  wire [7:0] a_sizes_set; // @[Monitor.scala 657:28]
  wire [7:0] _inflight_sizes_T; // @[Monitor.scala 704:39]
  wire [7:0] d_sizes_clr; // @[Monitor.scala 678:21]
  wire [7:0] _inflight_sizes_T_2; // @[Monitor.scala 704:54]
  reg [31:0] watchdog; // @[Monitor.scala 706:27]
  reg [31:0] _RAND_13;
  wire  _T_1034; // @[Monitor.scala 709:26]
  wire  _T_1036; // @[Monitor.scala 709:39]
  wire  _T_1037; // @[Monitor.scala 709:30]
  wire  _T_1038; // @[Monitor.scala 709:59]
  wire  _T_1039; // @[Monitor.scala 709:47]
  wire  _T_1041; // @[Monitor.scala 42:11]
  wire [31:0] _watchdog_T_1; // @[Monitor.scala 711:26]
  wire  _T_1045; // @[Monitor.scala 712:27]
  reg  inflight_1; // @[Monitor.scala 723:35]
  reg [31:0] _RAND_14;
  reg [7:0] inflight_sizes_1; // @[Monitor.scala 725:35]
  reg [31:0] _RAND_15;
  reg [8:0] d_first_counter_2; // @[Edges.scala 228:27]
  reg [31:0] _RAND_16;
  wire [8:0] d_first_counter1_2; // @[Edges.scala 229:28]
  wire  d_first_2; // @[Edges.scala 230:25]
  wire [15:0] _GEN_78; // @[Monitor.scala 747:93]
  wire [15:0] _c_size_lookup_T_6; // @[Monitor.scala 747:93]
  wire [15:0] _c_size_lookup_T_7; // @[Monitor.scala 747:146]
  wire  _T_1063; // @[Monitor.scala 779:26]
  wire  _T_1065; // @[Monitor.scala 779:71]
  wire [1:0] _GEN_66; // @[Monitor.scala 779:89]
  wire [30:0] _GEN_69; // @[Monitor.scala 783:90]
  wire  _T_1077; // @[Monitor.scala 49:11]
  wire [7:0] c_size_lookup; // @[Monitor.scala 747:21]
  wire  _T_1083; // @[Monitor.scala 795:36]
  wire  _T_1085; // @[Monitor.scala 49:11]
  wire  _T_1098; // @[Monitor.scala 804:28]
  wire  d_clr_wo_ready_1; // @[Monitor.scala 780:22]
  wire  _T_1101; // @[Monitor.scala 49:11]
  wire  _inflight_T_5; // @[Monitor.scala 809:44]
  wire [7:0] d_sizes_clr_1; // @[Monitor.scala 786:21]
  wire [7:0] _inflight_sizes_T_5; // @[Monitor.scala 811:56]
  reg [31:0] watchdog_1; // @[Monitor.scala 813:27]
  reg [31:0] _RAND_17;
  wire  _T_1103; // @[Monitor.scala 816:26]
  wire  _T_1105; // @[Monitor.scala 816:39]
  wire  _T_1106; // @[Monitor.scala 816:30]
  wire  _T_1107; // @[Monitor.scala 816:59]
  wire  _T_1108; // @[Monitor.scala 816:47]
  wire  _T_1110; // @[Monitor.scala 42:11]
  wire [31:0] _watchdog_T_3; // @[Monitor.scala 818:26]
  wire  _GEN_81; // @[Monitor.scala 49:11]
  wire  _GEN_89; // @[Monitor.scala 49:11]
  wire  _GEN_97; // @[Monitor.scala 49:11]
  wire  _GEN_105; // @[Monitor.scala 49:11]
  wire  _GEN_109; // @[Monitor.scala 49:11]
  wire  _GEN_113; // @[Monitor.scala 49:11]
  wire  _GEN_117; // @[Monitor.scala 49:11]
  wire  _GEN_122; // @[Monitor.scala 49:11]
  wire [29:0] TLMonitor_24_covSum;
  wire  stopEn0;
  wire  stopEn1;
  wire  stopEn2;
  wire  stopEn3;
  wire  stopEn4;
  wire  stopEn5;
  wire  stopEn6;
  wire  stopEn7;
  wire  stopEn8;
  wire  stopEn9;
  wire  stopEn10;
  wire  stopEn11;
  wire  stopEn12;
  wire  stopEn13;
  wire  stopEn14;
  wire  stopEn15;
  wire  stopEn16;
  wire  stopEn17;
  wire  stopEn18;
  wire  stopEn19;
  wire  stopEn20;
  wire  stopEn21;
  wire  stopEn22;
  wire  stopEn23;
  wire  stopEn24;
  wire  stopEn25;
  wire  stopEn26;
  wire  stopEn27;
  wire  stopEn28;
  wire  stopEn29;
  wire  stopEn30;
  wire  stopEn31;
  wire  stopEn32;
  wire  stopEn33;
  wire  stopEn34;
  wire  stopEn35;
  wire  stopEn36;
  wire  stopEn37;
  wire  stopEn38;
  wire  stopEn39;
  wire  plusarg_reader_metaAssert_wire;
  wire  plusarg_reader_1_metaAssert_wire;
  wire  TLMonitor_24_or15;
  wire  TLMonitor_24_or34;
  wire  TLMonitor_24_or16;
  wire  TLMonitor_24_or7;
  wire  TLMonitor_24_or17;
  wire  TLMonitor_24_or38;
  wire  TLMonitor_24_or18;
  wire  TLMonitor_24_or8;
  wire  TLMonitor_24_or3;
  wire  TLMonitor_24_or19;
  wire  TLMonitor_24_or42;
  wire  TLMonitor_24_or20;
  wire  TLMonitor_24_or9;
  wire  TLMonitor_24_or44;
  wire  TLMonitor_24_or21;
  wire  TLMonitor_24_or46;
  wire  TLMonitor_24_or22;
  wire  TLMonitor_24_or10;
  wire  TLMonitor_24_or4;
  wire  TLMonitor_24_or1;
  wire  TLMonitor_24_or23;
  wire  TLMonitor_24_or50;
  wire  TLMonitor_24_or24;
  wire  TLMonitor_24_or11;
  wire  TLMonitor_24_or25;
  wire  TLMonitor_24_or54;
  wire  TLMonitor_24_or26;
  wire  TLMonitor_24_or12;
  wire  TLMonitor_24_or5;
  wire  TLMonitor_24_or27;
  wire  TLMonitor_24_or58;
  wire  TLMonitor_24_or28;
  wire  TLMonitor_24_or13;
  wire  TLMonitor_24_or60;
  wire  TLMonitor_24_or29;
  wire  TLMonitor_24_or62;
  wire  TLMonitor_24_or30;
  wire  TLMonitor_24_or14;
  wire  TLMonitor_24_or6;
  wire  TLMonitor_24_or2;
  wire  TLMonitor_24_or0;
  reg  TLMonitor_24_metaAssert;
  reg [31:0] _RAND_18;
/*  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_out)
  );
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 ( // @[PlusArg.scala 80:11]
    .out(plusarg_reader_1_out)
  );*/
  assign _is_aligned_T = io_in_a_bits_address & 32'h3f; // @[Edges.scala 20:16]
  assign is_aligned = _is_aligned_T == 32'h0; // @[Edges.scala 20:24]
  assign _T_7 = {1'b0,$signed(io_in_a_bits_address)}; // @[Parameters.scala 137:49]
  assign _T_26 = $signed(_T_7) & -33'sh1000; // @[Parameters.scala 137:52]
  assign _T_27 = $signed(_T_26) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_28 = io_in_a_bits_address ^ 32'h3000; // @[Parameters.scala 137:31]
  assign _T_29 = {1'b0,$signed(_T_28)}; // @[Parameters.scala 137:49]
  assign _T_31 = $signed(_T_29) & -33'sh1000; // @[Parameters.scala 137:52]
  assign _T_32 = $signed(_T_31) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_33 = io_in_a_bits_address ^ 32'h10000; // @[Parameters.scala 137:31]
  assign _T_34 = {1'b0,$signed(_T_33)}; // @[Parameters.scala 137:49]
  assign _T_36 = $signed(_T_34) & -33'sh10000; // @[Parameters.scala 137:52]
  assign _T_37 = $signed(_T_36) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_38 = io_in_a_bits_address ^ 32'h2000000; // @[Parameters.scala 137:31]
  assign _T_39 = {1'b0,$signed(_T_38)}; // @[Parameters.scala 137:49]
  assign _T_41 = $signed(_T_39) & -33'sh10000; // @[Parameters.scala 137:52]
  assign _T_42 = $signed(_T_41) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_43 = io_in_a_bits_address ^ 32'hc000000; // @[Parameters.scala 137:31]
  assign _T_44 = {1'b0,$signed(_T_43)}; // @[Parameters.scala 137:49]
  assign _T_46 = $signed(_T_44) & -33'sh4000000; // @[Parameters.scala 137:52]
  assign _T_47 = $signed(_T_46) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_48 = io_in_a_bits_address ^ 32'h60000000; // @[Parameters.scala 137:31]
  assign _T_49 = {1'b0,$signed(_T_48)}; // @[Parameters.scala 137:49]
  assign _T_51 = $signed(_T_49) & -33'sh20000000; // @[Parameters.scala 137:52]
  assign _T_52 = $signed(_T_51) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_63 = io_in_a_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31]
  assign _T_64 = {1'b0,$signed(_T_63)}; // @[Parameters.scala 137:49]
  assign _T_66 = $signed(_T_64) & -33'sh10000000; // @[Parameters.scala 137:52]
  assign _T_67 = $signed(_T_66) == 33'sh0; // @[Parameters.scala 137:67]
  assign _T_134 = is_aligned | reset; // @[Monitor.scala 42:11]
  assign _T_341 = _T_27 | _T_37; // @[Parameters.scala 671:42]
  assign _T_342 = _T_341 | _T_42; // @[Parameters.scala 671:42]
  assign _T_343 = _T_342 | _T_47; // @[Parameters.scala 671:42]
  assign _T_344 = _T_343 | _T_52; // @[Parameters.scala 671:42]
  assign _T_345 = _T_344 | _T_67; // @[Parameters.scala 671:42]
  assign _T_348 = _T_32 | _T_345; // @[Parameters.scala 672:30]
  assign _T_350 = _T_348 | reset; // @[Monitor.scala 42:11]
  assign _T_766 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 42:24]
  assign _T_768 = _T_766 | reset; // @[Monitor.scala 49:11]
  assign _T_770 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25]
  assign _T_774 = io_in_d_bits_size >= 4'h3; // @[Monitor.scala 312:27]
  assign _T_776 = _T_774 | reset; // @[Monitor.scala 49:11]
  assign _T_778 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 313:28]
  assign _T_780 = _T_778 | reset; // @[Monitor.scala 49:11]
  assign _T_784 = ~io_in_d_bits_corrupt | reset; // @[Monitor.scala 49:11]
  assign _T_788 = ~io_in_d_bits_denied | reset; // @[Monitor.scala 49:11]
  assign _T_790 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25]
  assign _T_801 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 102:26]
  assign _T_803 = _T_801 | reset; // @[Monitor.scala 49:11]
  assign _T_805 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 323:28]
  assign _T_807 = _T_805 | reset; // @[Monitor.scala 49:11]
  assign _T_818 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25]
  assign _T_838 = ~io_in_d_bits_denied | io_in_d_bits_corrupt; // @[Monitor.scala 334:30]
  assign _T_840 = _T_838 | reset; // @[Monitor.scala 49:11]
  assign _T_847 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25]
  assign _T_864 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25]
  assign _T_882 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25]
  assign a_first_done = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37]
  assign a_first_counter1 = a_first_counter - 9'h1; // @[Edges.scala 229:28]
  assign a_first = a_first_counter == 9'h0; // @[Edges.scala 230:25]
  assign _T_912 = io_in_a_valid & ~a_first; // @[Monitor.scala 389:19]
  assign _T_929 = io_in_a_bits_address == address; // @[Monitor.scala 394:32]
  assign _T_931 = _T_929 | reset; // @[Monitor.scala 42:11]
  assign _T_934 = a_first_done & a_first; // @[Monitor.scala 396:20]
  assign _d_first_beats1_decode_T_1 = 27'hfff << io_in_d_bits_size; // @[package.scala 234:77]
  assign d_first_beats1_decode = ~_d_first_beats1_decode_T_1[11:3]; // @[Edges.scala 219:59]
  assign d_first_beats1_opdata = io_in_d_bits_opcode[0]; // @[Edges.scala 105:36]
  assign d_first_counter1 = d_first_counter - 9'h1; // @[Edges.scala 229:28]
  assign d_first = d_first_counter == 9'h0; // @[Edges.scala 230:25]
  assign _T_936 = io_in_d_valid & ~d_first; // @[Monitor.scala 541:19]
  assign _T_937 = io_in_d_bits_opcode == opcode_1; // @[Monitor.scala 542:29]
  assign _T_939 = _T_937 | reset; // @[Monitor.scala 49:11]
  assign _T_941 = io_in_d_bits_param == param_1; // @[Monitor.scala 543:29]
  assign _T_943 = _T_941 | reset; // @[Monitor.scala 49:11]
  assign _T_945 = io_in_d_bits_size == size_1; // @[Monitor.scala 544:29]
  assign _T_947 = _T_945 | reset; // @[Monitor.scala 49:11]
  assign _T_953 = io_in_d_bits_sink == sink; // @[Monitor.scala 546:29]
  assign _T_955 = _T_953 | reset; // @[Monitor.scala 49:11]
  assign _T_957 = io_in_d_bits_denied == denied; // @[Monitor.scala 547:29]
  assign _T_959 = _T_957 | reset; // @[Monitor.scala 49:11]
  assign _T_962 = io_in_d_valid & d_first; // @[Monitor.scala 549:20]
  assign a_first_counter1_1 = a_first_counter_1 - 9'h1; // @[Edges.scala 229:28]
  assign a_first_1 = a_first_counter_1 == 9'h0; // @[Edges.scala 230:25]
  assign d_first_counter1_1 = d_first_counter_1 - 9'h1; // @[Edges.scala 229:28]
  assign d_first_1 = d_first_counter_1 == 9'h0; // @[Edges.scala 230:25]
  assign _a_opcode_lookup_T_5 = 16'h10 - 16'h1; // @[Monitor.scala 609:57]
  assign _GEN_71 = {{12'd0}, inflight_opcodes}; // @[Monitor.scala 634:97]
  assign _a_opcode_lookup_T_6 = _GEN_71 & _a_opcode_lookup_T_5; // @[Monitor.scala 634:97]
  assign _a_opcode_lookup_T_7 = {{1'd0}, _a_opcode_lookup_T_6[15:1]}; // @[Monitor.scala 634:152]
  assign _a_size_lookup_T_5 = 16'h100 - 16'h1; // @[Monitor.scala 609:57]
  assign _GEN_73 = {{8'd0}, inflight_sizes}; // @[Monitor.scala 638:91]
  assign _a_size_lookup_T_6 = _GEN_73 & _a_size_lookup_T_5; // @[Monitor.scala 638:91]
  assign _a_size_lookup_T_7 = {{1'd0}, _a_size_lookup_T_6[15:1]}; // @[Monitor.scala 638:144]
  assign _T_963 = io_in_a_valid & a_first_1; // @[Monitor.scala 648:26]
  assign _GEN_15 = _T_963 ? 2'h1 : 2'h0; // @[Monitor.scala 648:71]
  assign _T_966 = a_first_done & a_first_1; // @[Monitor.scala 652:27]
  assign a_opcodes_set_interm = _T_966 ? 4'h9 : 4'h0; // @[Monitor.scala 652:72]
  assign _a_opcodes_set_T_1 = {{15'd0}, a_opcodes_set_interm}; // @[Monitor.scala 656:54]
  assign a_sizes_set_interm = _T_966 ? 5'hd : 5'h0; // @[Monitor.scala 652:72]
  assign _a_sizes_set_T_1 = {{15'd0}, a_sizes_set_interm}; // @[Monitor.scala 657:52]
  assign _T_972 = ~inflight | reset; // @[Monitor.scala 42:11]
  assign _GEN_16 = _T_966 ? 2'h1 : 2'h0; // @[Monitor.scala 652:72]
  assign _GEN_19 = _T_966 ? _a_opcodes_set_T_1 : 19'h0; // @[Monitor.scala 652:72]
  assign _GEN_20 = _T_966 ? _a_sizes_set_T_1 : 20'h0; // @[Monitor.scala 652:72]
  assign _T_974 = io_in_d_valid & d_first_1; // @[Monitor.scala 671:26]
  assign _T_977 = _T_974 & ~_T_770; // @[Monitor.scala 671:71]
  assign _GEN_21 = _T_977 ? 2'h1 : 2'h0; // @[Monitor.scala 671:90]
  assign _d_opcodes_clr_T_5 = {{15'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 677:76]
  assign _d_sizes_clr_T_5 = {{15'd0}, _a_size_lookup_T_5}; // @[Monitor.scala 678:74]
  assign _GEN_23 = _T_977 ? _d_opcodes_clr_T_5 : 31'h0; // @[Monitor.scala 675:91]
  assign _GEN_24 = _T_977 ? _d_sizes_clr_T_5 : 31'h0; // @[Monitor.scala 675:91]
  assign _T_989 = inflight | _T_963; // @[Monitor.scala 682:49]
  assign _T_991 = _T_989 | reset; // @[Monitor.scala 49:11]
  assign _T_995 = _T_864 | _T_864; // @[Monitor.scala 685:77]
  assign _T_997 = _T_995 | reset; // @[Monitor.scala 49:11]
  assign _T_999 = 4'h6 == io_in_d_bits_size; // @[Monitor.scala 687:36]
  assign _T_1001 = _T_999 | reset; // @[Monitor.scala 49:11]
  assign a_opcode_lookup = _a_opcode_lookup_T_7[3:0]; // @[Monitor.scala 634:21]
  assign _GEN_43 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 689:38]
  assign _GEN_44 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43; // @[Monitor.scala 689:38]
  assign _GEN_45 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44; // @[Monitor.scala 689:38]
  assign _GEN_46 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45; // @[Monitor.scala 689:38]
  assign _GEN_47 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46; // @[Monitor.scala 689:38]
  assign _GEN_48 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47; // @[Monitor.scala 689:38]
  assign _T_1004 = io_in_d_bits_opcode == _GEN_48; // @[Monitor.scala 689:38]
  assign _GEN_55 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46; // @[Monitor.scala 690:38]
  assign _GEN_56 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55; // @[Monitor.scala 690:38]
  assign _T_1006 = io_in_d_bits_opcode == _GEN_56; // @[Monitor.scala 690:38]
  assign _T_1007 = _T_1004 | _T_1006; // @[Monitor.scala 689:72]
  assign _T_1009 = _T_1007 | reset; // @[Monitor.scala 49:11]
  assign a_size_lookup = _a_size_lookup_T_7[7:0]; // @[Monitor.scala 638:19]
  assign _GEN_75 = {{4'd0}, io_in_d_bits_size}; // @[Monitor.scala 691:36]
  assign _T_1011 = _GEN_75 == a_size_lookup; // @[Monitor.scala 691:36]
  assign _T_1013 = _T_1011 | reset; // @[Monitor.scala 49:11]
  assign _T_1016 = _T_974 & a_first_1; // @[Monitor.scala 694:36]
  assign _T_1017 = _T_1016 & io_in_a_valid; // @[Monitor.scala 694:47]
  assign _T_1021 = _T_1017 & ~_T_770; // @[Monitor.scala 694:116]
  assign _T_1025 = io_in_a_ready | reset; // @[Monitor.scala 49:11]
  assign a_set_wo_ready = _GEN_15[0]; // @[Monitor.scala 649:22]
  assign d_clr_wo_ready = _GEN_21[0]; // @[Monitor.scala 672:22]
  assign _T_1027 = a_set_wo_ready != d_clr_wo_ready; // @[Monitor.scala 699:29]
  assign _T_1028 = |a_set_wo_ready; // @[Monitor.scala 699:67]
  assign _T_1030 = _T_1027 | ~_T_1028; // @[Monitor.scala 699:48]
  assign _T_1032 = _T_1030 | reset; // @[Monitor.scala 49:11]
  assign a_set = _GEN_16[0]; // @[Monitor.scala 653:28]
  assign _inflight_T = inflight | a_set; // @[Monitor.scala 702:27]
  assign _inflight_T_2 = _inflight_T & ~d_clr_wo_ready; // @[Monitor.scala 702:36]
  assign a_opcodes_set = _GEN_19[3:0]; // @[Monitor.scala 656:28]
  assign _inflight_opcodes_T = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 703:43]
  assign d_opcodes_clr = _GEN_23[3:0]; // @[Monitor.scala 677:21]
  assign _inflight_opcodes_T_2 = _inflight_opcodes_T & ~d_opcodes_clr; // @[Monitor.scala 703:60]
  assign a_sizes_set = _GEN_20[7:0]; // @[Monitor.scala 657:28]
  assign _inflight_sizes_T = inflight_sizes | a_sizes_set; // @[Monitor.scala 704:39]
  assign d_sizes_clr = _GEN_24[7:0]; // @[Monitor.scala 678:21]
  assign _inflight_sizes_T_2 = _inflight_sizes_T & ~d_sizes_clr; // @[Monitor.scala 704:54]
  assign _T_1034 = |inflight; // @[Monitor.scala 709:26]
  assign _T_1036 = plusarg_reader_out == 32'h0; // @[Monitor.scala 709:39]
  assign _T_1037 = ~_T_1034 | _T_1036; // @[Monitor.scala 709:30]
  assign _T_1038 = watchdog < plusarg_reader_out; // @[Monitor.scala 709:59]
  assign _T_1039 = _T_1037 | _T_1038; // @[Monitor.scala 709:47]
  assign _T_1041 = _T_1039 | reset; // @[Monitor.scala 42:11]
  assign _watchdog_T_1 = watchdog + 32'h1; // @[Monitor.scala 711:26]
  assign _T_1045 = a_first_done | io_in_d_valid; // @[Monitor.scala 712:27]
  assign d_first_counter1_2 = d_first_counter_2 - 9'h1; // @[Edges.scala 229:28]
  assign d_first_2 = d_first_counter_2 == 9'h0; // @[Edges.scala 230:25]
  assign _GEN_78 = {{8'd0}, inflight_sizes_1}; // @[Monitor.scala 747:93]
  assign _c_size_lookup_T_6 = _GEN_78 & _a_size_lookup_T_5; // @[Monitor.scala 747:93]
  assign _c_size_lookup_T_7 = {{1'd0}, _c_size_lookup_T_6[15:1]}; // @[Monitor.scala 747:146]
  assign _T_1063 = io_in_d_valid & d_first_2; // @[Monitor.scala 779:26]
  assign _T_1065 = _T_1063 & _T_770; // @[Monitor.scala 779:71]
  assign _GEN_66 = _T_1065 ? 2'h1 : 2'h0; // @[Monitor.scala 779:89]
  assign _GEN_69 = _T_1065 ? _d_sizes_clr_T_5 : 31'h0; // @[Monitor.scala 783:90]
  assign _T_1077 = inflight_1 | reset; // @[Monitor.scala 49:11]
  assign c_size_lookup = _c_size_lookup_T_7[7:0]; // @[Monitor.scala 747:21]
  assign _T_1083 = _GEN_75 == c_size_lookup; // @[Monitor.scala 795:36]
  assign _T_1085 = _T_1083 | reset; // @[Monitor.scala 49:11]
  assign _T_1098 = |1'h0; // @[Monitor.scala 804:28]
  assign d_clr_wo_ready_1 = _GEN_66[0]; // @[Monitor.scala 780:22]
  assign _T_1101 = d_clr_wo_ready_1 | reset; // @[Monitor.scala 49:11]
  assign _inflight_T_5 = inflight_1 & ~d_clr_wo_ready_1; // @[Monitor.scala 809:44]
  assign d_sizes_clr_1 = _GEN_69[7:0]; // @[Monitor.scala 786:21]
  assign _inflight_sizes_T_5 = inflight_sizes_1 & ~d_sizes_clr_1; // @[Monitor.scala 811:56]
  assign _T_1103 = |inflight_1; // @[Monitor.scala 816:26]
  assign _T_1105 = plusarg_reader_1_out == 32'h0; // @[Monitor.scala 816:39]
  assign _T_1106 = ~_T_1103 | _T_1105; // @[Monitor.scala 816:30]
  assign _T_1107 = watchdog_1 < plusarg_reader_1_out; // @[Monitor.scala 816:59]
  assign _T_1108 = _T_1106 | _T_1107; // @[Monitor.scala 816:47]
  assign _T_1110 = _T_1108 | reset; // @[Monitor.scala 42:11]
  assign _watchdog_T_3 = watchdog_1 + 32'h1; // @[Monitor.scala 818:26]
  assign _GEN_81 = io_in_d_valid & _T_770; // @[Monitor.scala 49:11]
  assign _GEN_89 = io_in_d_valid & _T_790; // @[Monitor.scala 49:11]
  assign _GEN_97 = io_in_d_valid & _T_818; // @[Monitor.scala 49:11]
  assign _GEN_105 = io_in_d_valid & _T_847; // @[Monitor.scala 49:11]
  assign _GEN_109 = io_in_d_valid & _T_864; // @[Monitor.scala 49:11]
  assign _GEN_113 = io_in_d_valid & _T_882; // @[Monitor.scala 49:11]
  assign _GEN_117 = _T_977 & _T_963; // @[Monitor.scala 49:11]
  assign _GEN_122 = _T_977 & ~_T_963; // @[Monitor.scala 49:11]
  assign TLMonitor_24_covSum = 30'h0;
  assign io_covSum = TLMonitor_24_covSum;
  assign stopEn0 = io_in_a_valid & ~_T_350;
  assign stopEn1 = io_in_a_valid & ~_T_134;
  assign stopEn2 = io_in_d_valid & ~_T_768;
  assign stopEn3 = _GEN_81 & ~_T_776;
  assign stopEn4 = _GEN_81 & ~_T_780;
  assign stopEn5 = _GEN_81 & ~_T_784;
  assign stopEn6 = _GEN_81 & ~_T_788;
  assign stopEn7 = _GEN_89 & ~_T_776;
  assign stopEn8 = _GEN_89 & ~_T_803;
  assign stopEn9 = _GEN_89 & ~_T_807;
  assign stopEn10 = _GEN_89 & ~_T_784;
  assign stopEn11 = _GEN_97 & ~_T_776;
  assign stopEn12 = _GEN_97 & ~_T_803;
  assign stopEn13 = _GEN_97 & ~_T_807;
  assign stopEn14 = _GEN_97 & ~_T_840;
  assign stopEn15 = _GEN_105 & ~_T_780;
  assign stopEn16 = _GEN_105 & ~_T_784;
  assign stopEn17 = _GEN_109 & ~_T_780;
  assign stopEn18 = _GEN_109 & ~_T_840;
  assign stopEn19 = _GEN_113 & ~_T_780;
  assign stopEn20 = _GEN_113 & ~_T_784;
  assign stopEn21 = _T_912 & ~_T_931;
  assign stopEn22 = _T_936 & ~_T_939;
  assign stopEn23 = _T_936 & ~_T_943;
  assign stopEn24 = _T_936 & ~_T_947;
  assign stopEn25 = _T_936 & ~_T_955;
  assign stopEn26 = _T_936 & ~_T_959;
  assign stopEn27 = _T_966 & ~_T_972;
  assign stopEn28 = _T_977 & ~_T_991;
  assign stopEn29 = _GEN_117 & ~_T_997;
  assign stopEn30 = _GEN_117 & ~_T_1001;
  assign stopEn31 = _GEN_122 & ~_T_1009;
  assign stopEn32 = _GEN_122 & ~_T_1013;
  assign stopEn33 = _T_1021 & ~_T_1025;
  assign stopEn34 = ~_T_1032;
  assign stopEn35 = ~_T_1041;
  assign stopEn36 = _T_1065 & ~_T_1077;
  assign stopEn37 = _T_1065 & ~_T_1085;
  assign stopEn38 = _T_1098 & ~_T_1101;
  assign stopEn39 = ~_T_1110;
//  assign plusarg_reader_metaAssert_wire = plusarg_reader_metaAssert;
//  assign plusarg_reader_1_metaAssert_wire = plusarg_reader_1_metaAssert;
  assign TLMonitor_24_or15 = stopEn0 | stopEn1;
  assign TLMonitor_24_or34 = stopEn3 | stopEn4;
  assign TLMonitor_24_or16 = stopEn2 | TLMonitor_24_or34;
  assign TLMonitor_24_or7 = TLMonitor_24_or15 | TLMonitor_24_or16;
  assign TLMonitor_24_or17 = stopEn5 | stopEn6;
  assign TLMonitor_24_or38 = stopEn8 | stopEn9;
  assign TLMonitor_24_or18 = stopEn7 | TLMonitor_24_or38;
  assign TLMonitor_24_or8 = TLMonitor_24_or17 | TLMonitor_24_or18;
  assign TLMonitor_24_or3 = TLMonitor_24_or7 | TLMonitor_24_or8;
  assign TLMonitor_24_or19 = stopEn10 | stopEn11;
  assign TLMonitor_24_or42 = stopEn13 | stopEn14;
  assign TLMonitor_24_or20 = stopEn12 | TLMonitor_24_or42;
  assign TLMonitor_24_or9 = TLMonitor_24_or19 | TLMonitor_24_or20;
  assign TLMonitor_24_or44 = stopEn16 | stopEn17;
  assign TLMonitor_24_or21 = stopEn15 | TLMonitor_24_or44;
  assign TLMonitor_24_or46 = stopEn19 | stopEn20;
  assign TLMonitor_24_or22 = stopEn18 | TLMonitor_24_or46;
  assign TLMonitor_24_or10 = TLMonitor_24_or21 | TLMonitor_24_or22;
  assign TLMonitor_24_or4 = TLMonitor_24_or9 | TLMonitor_24_or10;
  assign TLMonitor_24_or1 = TLMonitor_24_or3 | TLMonitor_24_or4;
  assign TLMonitor_24_or23 = stopEn21 | stopEn22;
  assign TLMonitor_24_or50 = stopEn24 | stopEn25;
  assign TLMonitor_24_or24 = stopEn23 | TLMonitor_24_or50;
  assign TLMonitor_24_or11 = TLMonitor_24_or23 | TLMonitor_24_or24;
  assign TLMonitor_24_or25 = stopEn26 | stopEn27;
  assign TLMonitor_24_or54 = stopEn29 | stopEn30;
  assign TLMonitor_24_or26 = stopEn28 | TLMonitor_24_or54;
  assign TLMonitor_24_or12 = TLMonitor_24_or25 | TLMonitor_24_or26;
  assign TLMonitor_24_or5 = TLMonitor_24_or11 | TLMonitor_24_or12;
  assign TLMonitor_24_or27 = stopEn31 | stopEn32;
  assign TLMonitor_24_or58 = stopEn34 | stopEn35;
  assign TLMonitor_24_or28 = stopEn33 | TLMonitor_24_or58;
  assign TLMonitor_24_or13 = TLMonitor_24_or27 | TLMonitor_24_or28;
  assign TLMonitor_24_or60 = stopEn37 | stopEn38;
  assign TLMonitor_24_or29 = stopEn36 | TLMonitor_24_or60;
  assign TLMonitor_24_or62 = plusarg_reader_metaAssert_wire | plusarg_reader_1_metaAssert_wire;
  assign TLMonitor_24_or30 = stopEn39 | TLMonitor_24_or62;
  assign TLMonitor_24_or14 = TLMonitor_24_or29 | TLMonitor_24_or30;
  assign TLMonitor_24_or6 = TLMonitor_24_or13 | TLMonitor_24_or14;
  assign TLMonitor_24_or2 = TLMonitor_24_or5 | TLMonitor_24_or6;
  assign TLMonitor_24_or0 = TLMonitor_24_or1 | TLMonitor_24_or2;
  assign metaAssert = TLMonitor_24_metaAssert;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  address = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  d_first_counter = _RAND_2[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  opcode_1 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  param_1 = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  size_1 = _RAND_5[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  sink = _RAND_6[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  denied = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  inflight = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  inflight_opcodes = _RAND_9[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  inflight_sizes = _RAND_10[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  a_first_counter_1 = _RAND_11[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  d_first_counter_1 = _RAND_12[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  watchdog = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  inflight_1 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  inflight_sizes_1 = _RAND_15[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  d_first_counter_2 = _RAND_16[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  watchdog_1 = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  TLMonitor_24_metaAssert = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      a_first_counter <= 9'h0;
    end else if (reset) begin
      a_first_counter <= 9'h0;
    end else if (a_first_done) begin
      if (a_first) begin
        a_first_counter <= 9'h0;
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (metaReset) begin
      address <= 32'h0;
    end else if (_T_934) begin
      address <= io_in_a_bits_address;
    end
    if (metaReset) begin
      d_first_counter <= 9'h0;
    end else if (reset) begin
      d_first_counter <= 9'h0;
    end else if (io_in_d_valid) begin
      if (d_first) begin
        if (d_first_beats1_opdata) begin
          d_first_counter <= d_first_beats1_decode;
        end else begin
          d_first_counter <= 9'h0;
        end
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    if (metaReset) begin
      opcode_1 <= 3'h0;
    end else if (_T_962) begin
      opcode_1 <= io_in_d_bits_opcode;
    end
    if (metaReset) begin
      param_1 <= 2'h0;
    end else if (_T_962) begin
      param_1 <= io_in_d_bits_param;
    end
    if (metaReset) begin
      size_1 <= 4'h0;
    end else if (_T_962) begin
      size_1 <= io_in_d_bits_size;
    end
    if (metaReset) begin
      sink <= 2'h0;
    end else if (_T_962) begin
      sink <= io_in_d_bits_sink;
    end
    if (metaReset) begin
      denied <= 1'h0;
    end else if (_T_962) begin
      denied <= io_in_d_bits_denied;
    end
    if (metaReset) begin
      inflight <= 1'h0;
    end else if (reset) begin
      inflight <= 1'h0;
    end else begin
      inflight <= _inflight_T_2;
    end
    if (metaReset) begin
      inflight_opcodes <= 4'h0;
    end else if (reset) begin
      inflight_opcodes <= 4'h0;
    end else begin
      inflight_opcodes <= _inflight_opcodes_T_2;
    end
    if (metaReset) begin
      inflight_sizes <= 8'h0;
    end else if (reset) begin
      inflight_sizes <= 8'h0;
    end else begin
      inflight_sizes <= _inflight_sizes_T_2;
    end
    if (metaReset) begin
      a_first_counter_1 <= 9'h0;
    end else if (reset) begin
      a_first_counter_1 <= 9'h0;
    end else if (a_first_done) begin
      if (a_first_1) begin
        a_first_counter_1 <= 9'h0;
      end else begin
        a_first_counter_1 <= a_first_counter1_1;
      end
    end
    if (metaReset) begin
      d_first_counter_1 <= 9'h0;
    end else if (reset) begin
      d_first_counter_1 <= 9'h0;
    end else if (io_in_d_valid) begin
      if (d_first_1) begin
        if (d_first_beats1_opdata) begin
          d_first_counter_1 <= d_first_beats1_decode;
        end else begin
          d_first_counter_1 <= 9'h0;
        end
      end else begin
        d_first_counter_1 <= d_first_counter1_1;
      end
    end
    if (metaReset) begin
      watchdog <= 32'h0;
    end else if (reset) begin
      watchdog <= 32'h0;
    end else if (_T_1045) begin
      watchdog <= 32'h0;
    end else begin
      watchdog <= _watchdog_T_1;
    end
    if (metaReset) begin
      inflight_1 <= 1'h0;
    end else if (reset) begin
      inflight_1 <= 1'h0;
    end else begin
      inflight_1 <= _inflight_T_5;
    end
    if (metaReset) begin
      inflight_sizes_1 <= 8'h0;
    end else if (reset) begin
      inflight_sizes_1 <= 8'h0;
    end else begin
      inflight_sizes_1 <= _inflight_sizes_T_5;
    end
    if (metaReset) begin
      d_first_counter_2 <= 9'h0;
    end else if (reset) begin
      d_first_counter_2 <= 9'h0;
    end else if (io_in_d_valid) begin
      if (d_first_2) begin
        if (d_first_beats1_opdata) begin
          d_first_counter_2 <= d_first_beats1_decode;
        end else begin
          d_first_counter_2 <= 9'h0;
        end
      end else begin
        d_first_counter_2 <= d_first_counter1_2;
      end
    end
    if (metaReset) begin
      watchdog_1 <= 32'h0;
    end else if (reset) begin
      watchdog_1 <= 32'h0;
    end else if (io_in_d_valid) begin
      watchdog_1 <= 32'h0;
    end else begin
      watchdog_1 <= _watchdog_T_3;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & ~_T_350) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at Frontend.scala:351:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & ~_T_350) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & ~_T_134) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get address not aligned to size (connected at Frontend.scala:351:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_a_valid & ~_T_134) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & ~_T_768) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel has invalid opcode (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & ~_T_768) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_81 & ~_T_776) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_81 & ~_T_776) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_81 & ~_T_780) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_81 & ~_T_780) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_81 & ~_T_784) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is corrupt (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_81 & ~_T_784) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_81 & ~_T_788) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is denied (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_81 & ~_T_788) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_89 & ~_T_776) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant smaller than a beat (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_89 & ~_T_776) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_89 & ~_T_803) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid cap param (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_89 & ~_T_803) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_89 & ~_T_807) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries toN param (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_89 & ~_T_807) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_89 & ~_T_784) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is corrupt (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_89 & ~_T_784) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_97 & ~_T_776) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData smaller than a beat (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_97 & ~_T_776) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_97 & ~_T_803) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid cap param (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_97 & ~_T_803) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_97 & ~_T_807) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries toN param (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_97 & ~_T_807) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_97 & ~_T_840) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_97 & ~_T_840) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & ~_T_780) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid param (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & ~_T_780) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & ~_T_784) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is corrupt (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & ~_T_784) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_109 & ~_T_780) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid param (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & ~_T_780) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_109 & ~_T_840) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & ~_T_840) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_113 & ~_T_780) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid param (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_113 & ~_T_780) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_113 & ~_T_784) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is corrupt (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_113 & ~_T_784) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_912 & ~_T_931) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel address changed with multibeat operation (connected at Frontend.scala:351:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_912 & ~_T_931) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_936 & ~_T_939) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel opcode changed within multibeat operation (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_936 & ~_T_939) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_936 & ~_T_943) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel param changed within multibeat operation (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_936 & ~_T_943) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_936 & ~_T_947) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel size changed within multibeat operation (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_936 & ~_T_947) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_936 & ~_T_955) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel sink changed with multibeat operation (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_936 & ~_T_955) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_936 & ~_T_959) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel denied changed with multibeat operation (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_936 & ~_T_959) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_966 & ~_T_972) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel re-used a source ID (connected at Frontend.scala:351:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_966 & ~_T_972) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_977 & ~_T_991) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel acknowledged for nothing inflight (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_977 & ~_T_991) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_117 & ~_T_997) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel contains improper opcode response (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_117 & ~_T_997) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_117 & ~_T_1001) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel contains improper response size (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_117 & ~_T_1001) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_122 & ~_T_1009) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel contains improper opcode response (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_122 & ~_T_1009) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_122 & ~_T_1013) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel contains improper response size (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_122 & ~_T_1013) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1021 & ~_T_1025) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1021 & ~_T_1025) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_1032) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' and 'D' concurrent, despite minlatency 3 (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_1032) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_1041) begin
          $fwrite(32'h80000002,"Assertion failed: TileLink timeout expired (connected at Frontend.scala:351:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_1041) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1065 & ~_T_1077) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel acknowledged for nothing inflight (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1065 & ~_T_1077) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1065 & ~_T_1085) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel contains improper response size (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1065 & ~_T_1085) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1098 & ~_T_1101) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' and 'D' concurrent, despite minlatency 3 (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1098 & ~_T_1101) begin
          $fatal; // @[Monitor.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_1110) begin
          $fwrite(32'h80000002,"Assertion failed: TileLink timeout expired (connected at Frontend.scala:351:21)\n    at Monitor.scala:42 assert(cond, message)\n"); // @[Monitor.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_1110) begin
          $fatal; // @[Monitor.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    if (metaReset) begin
      TLMonitor_24_metaAssert <= 1'h0;
    end else begin
      TLMonitor_24_metaAssert <= TLMonitor_24_metaAssert | TLMonitor_24_or0;
    end
  end
endmodule
module TLB(
  input         clock,
  input         reset,
  output        io_req_ready,
  input         io_req_valid,
  input  [39:0] io_req_bits_vaddr,
  input         io_req_bits_passthrough,
  input  [1:0]  io_req_bits_size,
  input  [4:0]  io_req_bits_cmd,
  output        io_resp_miss,
  output [31:0] io_resp_paddr,
  output        io_resp_pf_ld,
  output        io_resp_pf_st,
  output        io_resp_ae_ld,
  output        io_resp_ae_st,
  output        io_resp_ma_ld,
  output        io_resp_ma_st,
  output        io_resp_cacheable,
  input         io_sfence_valid,
  input         io_sfence_bits_rs1,
  input         io_sfence_bits_rs2,
  input  [38:0] io_sfence_bits_addr,
  input         io_ptw_req_ready,
  output        io_ptw_req_valid,
  output [26:0] io_ptw_req_bits_bits_addr,
  input         io_ptw_resp_valid,
  input         io_ptw_resp_bits_ae,
  input  [53:0] io_ptw_resp_bits_pte_ppn,
  input         io_ptw_resp_bits_pte_d,
  input         io_ptw_resp_bits_pte_a,
  input         io_ptw_resp_bits_pte_g,
  input         io_ptw_resp_bits_pte_u,
  input         io_ptw_resp_bits_pte_x,
  input         io_ptw_resp_bits_pte_w,
  input         io_ptw_resp_bits_pte_r,
  input         io_ptw_resp_bits_pte_v,
  input  [1:0]  io_ptw_resp_bits_level,
  input         io_ptw_resp_bits_homogeneous,
  input  [3:0]  io_ptw_ptbr_mode,
  input         io_ptw_status_debug,
  input  [1:0]  io_ptw_status_dprv,
  input         io_ptw_status_mxr,
  input         io_ptw_status_sum,
  input         io_ptw_pmp_0_cfg_l,
  input  [1:0]  io_ptw_pmp_0_cfg_a,
  input         io_ptw_pmp_0_cfg_x,
  input         io_ptw_pmp_0_cfg_w,
  input         io_ptw_pmp_0_cfg_r,
  input  [29:0] io_ptw_pmp_0_addr,
  input  [31:0] io_ptw_pmp_0_mask,
  input         io_ptw_pmp_1_cfg_l,
  input  [1:0]  io_ptw_pmp_1_cfg_a,
  input         io_ptw_pmp_1_cfg_x,
  input         io_ptw_pmp_1_cfg_w,
  input         io_ptw_pmp_1_cfg_r,
  input  [29:0] io_ptw_pmp_1_addr,
  input  [31:0] io_ptw_pmp_1_mask,
  input         io_ptw_pmp_2_cfg_l,
  input  [1:0]  io_ptw_pmp_2_cfg_a,
  input         io_ptw_pmp_2_cfg_x,
  input         io_ptw_pmp_2_cfg_w,
  input         io_ptw_pmp_2_cfg_r,
  input  [29:0] io_ptw_pmp_2_addr,
  input  [31:0] io_ptw_pmp_2_mask,
  input         io_ptw_pmp_3_cfg_l,
  input  [1:0]  io_ptw_pmp_3_cfg_a,
  input         io_ptw_pmp_3_cfg_x,
  input         io_ptw_pmp_3_cfg_w,
  input         io_ptw_pmp_3_cfg_r,
  input  [29:0] io_ptw_pmp_3_addr,
  input  [31:0] io_ptw_pmp_3_mask,
  input         io_ptw_pmp_4_cfg_l,
  input  [1:0]  io_ptw_pmp_4_cfg_a,
  input         io_ptw_pmp_4_cfg_x,
  input         io_ptw_pmp_4_cfg_w,
  input         io_ptw_pmp_4_cfg_r,
  input  [29:0] io_ptw_pmp_4_addr,
  input  [31:0] io_ptw_pmp_4_mask,
  input         io_ptw_pmp_5_cfg_l,
  input  [1:0]  io_ptw_pmp_5_cfg_a,
  input         io_ptw_pmp_5_cfg_x,
  input         io_ptw_pmp_5_cfg_w,
  input         io_ptw_pmp_5_cfg_r,
  input  [29:0] io_ptw_pmp_5_addr,
  input  [31:0] io_ptw_pmp_5_mask,
  input         io_ptw_pmp_6_cfg_l,
  input  [1:0]  io_ptw_pmp_6_cfg_a,
  input         io_ptw_pmp_6_cfg_x,
  input         io_ptw_pmp_6_cfg_w,
  input         io_ptw_pmp_6_cfg_r,
  input  [29:0] io_ptw_pmp_6_addr,
  input  [31:0] io_ptw_pmp_6_mask,
  input         io_ptw_pmp_7_cfg_l,
  input  [1:0]  io_ptw_pmp_7_cfg_a,
  input         io_ptw_pmp_7_cfg_x,
  input         io_ptw_pmp_7_cfg_w,
  input         io_ptw_pmp_7_cfg_r,
  input  [29:0] io_ptw_pmp_7_addr,
  input  [31:0] io_ptw_pmp_7_mask,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  wire [19:0] mpu_ppn_barrier_io_x_ppn; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_x_u; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_x_ae; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_x_sw; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_x_sx; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_x_sr; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_x_pw; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_x_px; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_x_pr; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_x_ppp; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_x_pal; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_x_paa; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_x_eff; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_x_c; // @[package.scala 258:25]
  wire [19:0] mpu_ppn_barrier_io_y_ppn; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_y_u; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_y_ae; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_y_sw; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_y_sx; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_y_sr; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_y_pw; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_y_px; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_y_pr; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_y_ppp; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_y_pal; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_y_paa; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_y_eff; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_y_c; // @[package.scala 258:25]
  wire [29:0] mpu_ppn_barrier_io_covSum; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_metaAssert; // @[package.scala 258:25]
  wire [1:0] pmp_io_prv; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_0_cfg_l; // @[TLB.scala 192:19]
  wire [1:0] pmp_io_pmp_0_cfg_a; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_0_cfg_x; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_0_cfg_w; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_0_cfg_r; // @[TLB.scala 192:19]
  wire [29:0] pmp_io_pmp_0_addr; // @[TLB.scala 192:19]
  wire [31:0] pmp_io_pmp_0_mask; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_1_cfg_l; // @[TLB.scala 192:19]
  wire [1:0] pmp_io_pmp_1_cfg_a; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_1_cfg_x; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_1_cfg_w; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_1_cfg_r; // @[TLB.scala 192:19]
  wire [29:0] pmp_io_pmp_1_addr; // @[TLB.scala 192:19]
  wire [31:0] pmp_io_pmp_1_mask; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_2_cfg_l; // @[TLB.scala 192:19]
  wire [1:0] pmp_io_pmp_2_cfg_a; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_2_cfg_x; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_2_cfg_w; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_2_cfg_r; // @[TLB.scala 192:19]
  wire [29:0] pmp_io_pmp_2_addr; // @[TLB.scala 192:19]
  wire [31:0] pmp_io_pmp_2_mask; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_3_cfg_l; // @[TLB.scala 192:19]
  wire [1:0] pmp_io_pmp_3_cfg_a; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_3_cfg_x; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_3_cfg_w; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_3_cfg_r; // @[TLB.scala 192:19]
  wire [29:0] pmp_io_pmp_3_addr; // @[TLB.scala 192:19]
  wire [31:0] pmp_io_pmp_3_mask; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_4_cfg_l; // @[TLB.scala 192:19]
  wire [1:0] pmp_io_pmp_4_cfg_a; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_4_cfg_x; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_4_cfg_w; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_4_cfg_r; // @[TLB.scala 192:19]
  wire [29:0] pmp_io_pmp_4_addr; // @[TLB.scala 192:19]
  wire [31:0] pmp_io_pmp_4_mask; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_5_cfg_l; // @[TLB.scala 192:19]
  wire [1:0] pmp_io_pmp_5_cfg_a; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_5_cfg_x; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_5_cfg_w; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_5_cfg_r; // @[TLB.scala 192:19]
  wire [29:0] pmp_io_pmp_5_addr; // @[TLB.scala 192:19]
  wire [31:0] pmp_io_pmp_5_mask; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_6_cfg_l; // @[TLB.scala 192:19]
  wire [1:0] pmp_io_pmp_6_cfg_a; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_6_cfg_x; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_6_cfg_w; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_6_cfg_r; // @[TLB.scala 192:19]
  wire [29:0] pmp_io_pmp_6_addr; // @[TLB.scala 192:19]
  wire [31:0] pmp_io_pmp_6_mask; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_7_cfg_l; // @[TLB.scala 192:19]
  wire [1:0] pmp_io_pmp_7_cfg_a; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_7_cfg_x; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_7_cfg_w; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_7_cfg_r; // @[TLB.scala 192:19]
  wire [29:0] pmp_io_pmp_7_addr; // @[TLB.scala 192:19]
  wire [31:0] pmp_io_pmp_7_mask; // @[TLB.scala 192:19]
  wire [31:0] pmp_io_addr; // @[TLB.scala 192:19]
  wire [1:0] pmp_io_size; // @[TLB.scala 192:19]
  wire  pmp_io_r; // @[TLB.scala 192:19]
  wire  pmp_io_w; // @[TLB.scala 192:19]
  wire  pmp_io_x; // @[TLB.scala 192:19]
  wire [29:0] pmp_io_covSum; // @[TLB.scala 192:19]
  wire  pmp_metaAssert; // @[TLB.scala 192:19]
  wire [19:0] entries_barrier_io_x_ppn; // @[package.scala 258:25]
  wire  entries_barrier_io_x_u; // @[package.scala 258:25]
  wire  entries_barrier_io_x_ae; // @[package.scala 258:25]
  wire  entries_barrier_io_x_sw; // @[package.scala 258:25]
  wire  entries_barrier_io_x_sx; // @[package.scala 258:25]
  wire  entries_barrier_io_x_sr; // @[package.scala 258:25]
  wire  entries_barrier_io_x_pw; // @[package.scala 258:25]
  wire  entries_barrier_io_x_px; // @[package.scala 258:25]
  wire  entries_barrier_io_x_pr; // @[package.scala 258:25]
  wire  entries_barrier_io_x_ppp; // @[package.scala 258:25]
  wire  entries_barrier_io_x_pal; // @[package.scala 258:25]
  wire  entries_barrier_io_x_paa; // @[package.scala 258:25]
  wire  entries_barrier_io_x_eff; // @[package.scala 258:25]
  wire  entries_barrier_io_x_c; // @[package.scala 258:25]
  wire [19:0] entries_barrier_io_y_ppn; // @[package.scala 258:25]
  wire  entries_barrier_io_y_u; // @[package.scala 258:25]
  wire  entries_barrier_io_y_ae; // @[package.scala 258:25]
  wire  entries_barrier_io_y_sw; // @[package.scala 258:25]
  wire  entries_barrier_io_y_sx; // @[package.scala 258:25]
  wire  entries_barrier_io_y_sr; // @[package.scala 258:25]
  wire  entries_barrier_io_y_pw; // @[package.scala 258:25]
  wire  entries_barrier_io_y_px; // @[package.scala 258:25]
  wire  entries_barrier_io_y_pr; // @[package.scala 258:25]
  wire  entries_barrier_io_y_ppp; // @[package.scala 258:25]
  wire  entries_barrier_io_y_pal; // @[package.scala 258:25]
  wire  entries_barrier_io_y_paa; // @[package.scala 258:25]
  wire  entries_barrier_io_y_eff; // @[package.scala 258:25]
  wire  entries_barrier_io_y_c; // @[package.scala 258:25]
  wire [29:0] entries_barrier_io_covSum; // @[package.scala 258:25]
  wire  entries_barrier_metaAssert; // @[package.scala 258:25]
  wire [19:0] entries_barrier_1_io_x_ppn; // @[package.scala 258:25]
  wire  entries_barrier_1_io_x_u; // @[package.scala 258:25]
  wire  entries_barrier_1_io_x_ae; // @[package.scala 258:25]
  wire  entries_barrier_1_io_x_sw; // @[package.scala 258:25]
  wire  entries_barrier_1_io_x_sx; // @[package.scala 258:25]
  wire  entries_barrier_1_io_x_sr; // @[package.scala 258:25]
  wire  entries_barrier_1_io_x_pw; // @[package.scala 258:25]
  wire  entries_barrier_1_io_x_px; // @[package.scala 258:25]
  wire  entries_barrier_1_io_x_pr; // @[package.scala 258:25]
  wire  entries_barrier_1_io_x_ppp; // @[package.scala 258:25]
  wire  entries_barrier_1_io_x_pal; // @[package.scala 258:25]
  wire  entries_barrier_1_io_x_paa; // @[package.scala 258:25]
  wire  entries_barrier_1_io_x_eff; // @[package.scala 258:25]
  wire  entries_barrier_1_io_x_c; // @[package.scala 258:25]
  wire [19:0] entries_barrier_1_io_y_ppn; // @[package.scala 258:25]
  wire  entries_barrier_1_io_y_u; // @[package.scala 258:25]
  wire  entries_barrier_1_io_y_ae; // @[package.scala 258:25]
  wire  entries_barrier_1_io_y_sw; // @[package.scala 258:25]
  wire  entries_barrier_1_io_y_sx; // @[package.scala 258:25]
  wire  entries_barrier_1_io_y_sr; // @[package.scala 258:25]
  wire  entries_barrier_1_io_y_pw; // @[package.scala 258:25]
  wire  entries_barrier_1_io_y_px; // @[package.scala 258:25]
  wire  entries_barrier_1_io_y_pr; // @[package.scala 258:25]
  wire  entries_barrier_1_io_y_ppp; // @[package.scala 258:25]
  wire  entries_barrier_1_io_y_pal; // @[package.scala 258:25]
  wire  entries_barrier_1_io_y_paa; // @[package.scala 258:25]
  wire  entries_barrier_1_io_y_eff; // @[package.scala 258:25]
  wire  entries_barrier_1_io_y_c; // @[package.scala 258:25]
  wire [29:0] entries_barrier_1_io_covSum; // @[package.scala 258:25]
  wire  entries_barrier_1_metaAssert; // @[package.scala 258:25]
  wire [19:0] entries_barrier_2_io_x_ppn; // @[package.scala 258:25]
  wire  entries_barrier_2_io_x_u; // @[package.scala 258:25]
  wire  entries_barrier_2_io_x_ae; // @[package.scala 258:25]
  wire  entries_barrier_2_io_x_sw; // @[package.scala 258:25]
  wire  entries_barrier_2_io_x_sx; // @[package.scala 258:25]
  wire  entries_barrier_2_io_x_sr; // @[package.scala 258:25]
  wire  entries_barrier_2_io_x_pw; // @[package.scala 258:25]
  wire  entries_barrier_2_io_x_px; // @[package.scala 258:25]
  wire  entries_barrier_2_io_x_pr; // @[package.scala 258:25]
  wire  entries_barrier_2_io_x_ppp; // @[package.scala 258:25]
  wire  entries_barrier_2_io_x_pal; // @[package.scala 258:25]
  wire  entries_barrier_2_io_x_paa; // @[package.scala 258:25]
  wire  entries_barrier_2_io_x_eff; // @[package.scala 258:25]
  wire  entries_barrier_2_io_x_c; // @[package.scala 258:25]
  wire [19:0] entries_barrier_2_io_y_ppn; // @[package.scala 258:25]
  wire  entries_barrier_2_io_y_u; // @[package.scala 258:25]
  wire  entries_barrier_2_io_y_ae; // @[package.scala 258:25]
  wire  entries_barrier_2_io_y_sw; // @[package.scala 258:25]
  wire  entries_barrier_2_io_y_sx; // @[package.scala 258:25]
  wire  entries_barrier_2_io_y_sr; // @[package.scala 258:25]
  wire  entries_barrier_2_io_y_pw; // @[package.scala 258:25]
  wire  entries_barrier_2_io_y_px; // @[package.scala 258:25]
  wire  entries_barrier_2_io_y_pr; // @[package.scala 258:25]
  wire  entries_barrier_2_io_y_ppp; // @[package.scala 258:25]
  wire  entries_barrier_2_io_y_pal; // @[package.scala 258:25]
  wire  entries_barrier_2_io_y_paa; // @[package.scala 258:25]
  wire  entries_barrier_2_io_y_eff; // @[package.scala 258:25]
  wire  entries_barrier_2_io_y_c; // @[package.scala 258:25]
  wire [29:0] entries_barrier_2_io_covSum; // @[package.scala 258:25]
  wire  entries_barrier_2_metaAssert; // @[package.scala 258:25]
  wire [19:0] entries_barrier_3_io_x_ppn; // @[package.scala 258:25]
  wire  entries_barrier_3_io_x_u; // @[package.scala 258:25]
  wire  entries_barrier_3_io_x_ae; // @[package.scala 258:25]
  wire  entries_barrier_3_io_x_sw; // @[package.scala 258:25]
  wire  entries_barrier_3_io_x_sx; // @[package.scala 258:25]
  wire  entries_barrier_3_io_x_sr; // @[package.scala 258:25]
  wire  entries_barrier_3_io_x_pw; // @[package.scala 258:25]
  wire  entries_barrier_3_io_x_px; // @[package.scala 258:25]
  wire  entries_barrier_3_io_x_pr; // @[package.scala 258:25]
  wire  entries_barrier_3_io_x_ppp; // @[package.scala 258:25]
  wire  entries_barrier_3_io_x_pal; // @[package.scala 258:25]
  wire  entries_barrier_3_io_x_paa; // @[package.scala 258:25]
  wire  entries_barrier_3_io_x_eff; // @[package.scala 258:25]
  wire  entries_barrier_3_io_x_c; // @[package.scala 258:25]
  wire [19:0] entries_barrier_3_io_y_ppn; // @[package.scala 258:25]
  wire  entries_barrier_3_io_y_u; // @[package.scala 258:25]
  wire  entries_barrier_3_io_y_ae; // @[package.scala 258:25]
  wire  entries_barrier_3_io_y_sw; // @[package.scala 258:25]
  wire  entries_barrier_3_io_y_sx; // @[package.scala 258:25]
  wire  entries_barrier_3_io_y_sr; // @[package.scala 258:25]
  wire  entries_barrier_3_io_y_pw; // @[package.scala 258:25]
  wire  entries_barrier_3_io_y_px; // @[package.scala 258:25]
  wire  entries_barrier_3_io_y_pr; // @[package.scala 258:25]
  wire  entries_barrier_3_io_y_ppp; // @[package.scala 258:25]
  wire  entries_barrier_3_io_y_pal; // @[package.scala 258:25]
  wire  entries_barrier_3_io_y_paa; // @[package.scala 258:25]
  wire  entries_barrier_3_io_y_eff; // @[package.scala 258:25]
  wire  entries_barrier_3_io_y_c; // @[package.scala 258:25]
  wire [29:0] entries_barrier_3_io_covSum; // @[package.scala 258:25]
  wire  entries_barrier_3_metaAssert; // @[package.scala 258:25]
  wire [19:0] entries_barrier_4_io_x_ppn; // @[package.scala 258:25]
  wire  entries_barrier_4_io_x_u; // @[package.scala 258:25]
  wire  entries_barrier_4_io_x_ae; // @[package.scala 258:25]
  wire  entries_barrier_4_io_x_sw; // @[package.scala 258:25]
  wire  entries_barrier_4_io_x_sx; // @[package.scala 258:25]
  wire  entries_barrier_4_io_x_sr; // @[package.scala 258:25]
  wire  entries_barrier_4_io_x_pw; // @[package.scala 258:25]
  wire  entries_barrier_4_io_x_px; // @[package.scala 258:25]
  wire  entries_barrier_4_io_x_pr; // @[package.scala 258:25]
  wire  entries_barrier_4_io_x_ppp; // @[package.scala 258:25]
  wire  entries_barrier_4_io_x_pal; // @[package.scala 258:25]
  wire  entries_barrier_4_io_x_paa; // @[package.scala 258:25]
  wire  entries_barrier_4_io_x_eff; // @[package.scala 258:25]
  wire  entries_barrier_4_io_x_c; // @[package.scala 258:25]
  wire [19:0] entries_barrier_4_io_y_ppn; // @[package.scala 258:25]
  wire  entries_barrier_4_io_y_u; // @[package.scala 258:25]
  wire  entries_barrier_4_io_y_ae; // @[package.scala 258:25]
  wire  entries_barrier_4_io_y_sw; // @[package.scala 258:25]
  wire  entries_barrier_4_io_y_sx; // @[package.scala 258:25]
  wire  entries_barrier_4_io_y_sr; // @[package.scala 258:25]
  wire  entries_barrier_4_io_y_pw; // @[package.scala 258:25]
  wire  entries_barrier_4_io_y_px; // @[package.scala 258:25]
  wire  entries_barrier_4_io_y_pr; // @[package.scala 258:25]
  wire  entries_barrier_4_io_y_ppp; // @[package.scala 258:25]
  wire  entries_barrier_4_io_y_pal; // @[package.scala 258:25]
  wire  entries_barrier_4_io_y_paa; // @[package.scala 258:25]
  wire  entries_barrier_4_io_y_eff; // @[package.scala 258:25]
  wire  entries_barrier_4_io_y_c; // @[package.scala 258:25]
  wire [29:0] entries_barrier_4_io_covSum; // @[package.scala 258:25]
  wire  entries_barrier_4_metaAssert; // @[package.scala 258:25]
  wire [19:0] entries_barrier_5_io_x_ppn; // @[package.scala 258:25]
  wire  entries_barrier_5_io_x_u; // @[package.scala 258:25]
  wire  entries_barrier_5_io_x_ae; // @[package.scala 258:25]
  wire  entries_barrier_5_io_x_sw; // @[package.scala 258:25]
  wire  entries_barrier_5_io_x_sx; // @[package.scala 258:25]
  wire  entries_barrier_5_io_x_sr; // @[package.scala 258:25]
  wire  entries_barrier_5_io_x_pw; // @[package.scala 258:25]
  wire  entries_barrier_5_io_x_px; // @[package.scala 258:25]
  wire  entries_barrier_5_io_x_pr; // @[package.scala 258:25]
  wire  entries_barrier_5_io_x_ppp; // @[package.scala 258:25]
  wire  entries_barrier_5_io_x_pal; // @[package.scala 258:25]
  wire  entries_barrier_5_io_x_paa; // @[package.scala 258:25]
  wire  entries_barrier_5_io_x_eff; // @[package.scala 258:25]
  wire  entries_barrier_5_io_x_c; // @[package.scala 258:25]
  wire [19:0] entries_barrier_5_io_y_ppn; // @[package.scala 258:25]
  wire  entries_barrier_5_io_y_u; // @[package.scala 258:25]
  wire  entries_barrier_5_io_y_ae; // @[package.scala 258:25]
  wire  entries_barrier_5_io_y_sw; // @[package.scala 258:25]
  wire  entries_barrier_5_io_y_sx; // @[package.scala 258:25]
  wire  entries_barrier_5_io_y_sr; // @[package.scala 258:25]
  wire  entries_barrier_5_io_y_pw; // @[package.scala 258:25]
  wire  entries_barrier_5_io_y_px; // @[package.scala 258:25]
  wire  entries_barrier_5_io_y_pr; // @[package.scala 258:25]
  wire  entries_barrier_5_io_y_ppp; // @[package.scala 258:25]
  wire  entries_barrier_5_io_y_pal; // @[package.scala 258:25]
  wire  entries_barrier_5_io_y_paa; // @[package.scala 258:25]
  wire  entries_barrier_5_io_y_eff; // @[package.scala 258:25]
  wire  entries_barrier_5_io_y_c; // @[package.scala 258:25]
  wire [29:0] entries_barrier_5_io_covSum; // @[package.scala 258:25]
  wire  entries_barrier_5_metaAssert; // @[package.scala 258:25]
  wire [19:0] entries_barrier_6_io_x_ppn; // @[package.scala 258:25]
  wire  entries_barrier_6_io_x_u; // @[package.scala 258:25]
  wire  entries_barrier_6_io_x_ae; // @[package.scala 258:25]
  wire  entries_barrier_6_io_x_sw; // @[package.scala 258:25]
  wire  entries_barrier_6_io_x_sx; // @[package.scala 258:25]
  wire  entries_barrier_6_io_x_sr; // @[package.scala 258:25]
  wire  entries_barrier_6_io_x_pw; // @[package.scala 258:25]
  wire  entries_barrier_6_io_x_px; // @[package.scala 258:25]
  wire  entries_barrier_6_io_x_pr; // @[package.scala 258:25]
  wire  entries_barrier_6_io_x_ppp; // @[package.scala 258:25]
  wire  entries_barrier_6_io_x_pal; // @[package.scala 258:25]
  wire  entries_barrier_6_io_x_paa; // @[package.scala 258:25]
  wire  entries_barrier_6_io_x_eff; // @[package.scala 258:25]
  wire  entries_barrier_6_io_x_c; // @[package.scala 258:25]
  wire [19:0] entries_barrier_6_io_y_ppn; // @[package.scala 258:25]
  wire  entries_barrier_6_io_y_u; // @[package.scala 258:25]
  wire  entries_barrier_6_io_y_ae; // @[package.scala 258:25]
  wire  entries_barrier_6_io_y_sw; // @[package.scala 258:25]
  wire  entries_barrier_6_io_y_sx; // @[package.scala 258:25]
  wire  entries_barrier_6_io_y_sr; // @[package.scala 258:25]
  wire  entries_barrier_6_io_y_pw; // @[package.scala 258:25]
  wire  entries_barrier_6_io_y_px; // @[package.scala 258:25]
  wire  entries_barrier_6_io_y_pr; // @[package.scala 258:25]
  wire  entries_barrier_6_io_y_ppp; // @[package.scala 258:25]
  wire  entries_barrier_6_io_y_pal; // @[package.scala 258:25]
  wire  entries_barrier_6_io_y_paa; // @[package.scala 258:25]
  wire  entries_barrier_6_io_y_eff; // @[package.scala 258:25]
  wire  entries_barrier_6_io_y_c; // @[package.scala 258:25]
  wire [29:0] entries_barrier_6_io_covSum; // @[package.scala 258:25]
  wire  entries_barrier_6_metaAssert; // @[package.scala 258:25]
  wire [19:0] entries_barrier_7_io_x_ppn; // @[package.scala 258:25]
  wire  entries_barrier_7_io_x_u; // @[package.scala 258:25]
  wire  entries_barrier_7_io_x_ae; // @[package.scala 258:25]
  wire  entries_barrier_7_io_x_sw; // @[package.scala 258:25]
  wire  entries_barrier_7_io_x_sx; // @[package.scala 258:25]
  wire  entries_barrier_7_io_x_sr; // @[package.scala 258:25]
  wire  entries_barrier_7_io_x_pw; // @[package.scala 258:25]
  wire  entries_barrier_7_io_x_px; // @[package.scala 258:25]
  wire  entries_barrier_7_io_x_pr; // @[package.scala 258:25]
  wire  entries_barrier_7_io_x_ppp; // @[package.scala 258:25]
  wire  entries_barrier_7_io_x_pal; // @[package.scala 258:25]
  wire  entries_barrier_7_io_x_paa; // @[package.scala 258:25]
  wire  entries_barrier_7_io_x_eff; // @[package.scala 258:25]
  wire  entries_barrier_7_io_x_c; // @[package.scala 258:25]
  wire [19:0] entries_barrier_7_io_y_ppn; // @[package.scala 258:25]
  wire  entries_barrier_7_io_y_u; // @[package.scala 258:25]
  wire  entries_barrier_7_io_y_ae; // @[package.scala 258:25]
  wire  entries_barrier_7_io_y_sw; // @[package.scala 258:25]
  wire  entries_barrier_7_io_y_sx; // @[package.scala 258:25]
  wire  entries_barrier_7_io_y_sr; // @[package.scala 258:25]
  wire  entries_barrier_7_io_y_pw; // @[package.scala 258:25]
  wire  entries_barrier_7_io_y_px; // @[package.scala 258:25]
  wire  entries_barrier_7_io_y_pr; // @[package.scala 258:25]
  wire  entries_barrier_7_io_y_ppp; // @[package.scala 258:25]
  wire  entries_barrier_7_io_y_pal; // @[package.scala 258:25]
  wire  entries_barrier_7_io_y_paa; // @[package.scala 258:25]
  wire  entries_barrier_7_io_y_eff; // @[package.scala 258:25]
  wire  entries_barrier_7_io_y_c; // @[package.scala 258:25]
  wire [29:0] entries_barrier_7_io_covSum; // @[package.scala 258:25]
  wire  entries_barrier_7_metaAssert; // @[package.scala 258:25]
  wire [19:0] entries_barrier_8_io_x_ppn; // @[package.scala 258:25]
  wire  entries_barrier_8_io_x_u; // @[package.scala 258:25]
  wire  entries_barrier_8_io_x_ae; // @[package.scala 258:25]
  wire  entries_barrier_8_io_x_sw; // @[package.scala 258:25]
  wire  entries_barrier_8_io_x_sx; // @[package.scala 258:25]
  wire  entries_barrier_8_io_x_sr; // @[package.scala 258:25]
  wire  entries_barrier_8_io_x_pw; // @[package.scala 258:25]
  wire  entries_barrier_8_io_x_px; // @[package.scala 258:25]
  wire  entries_barrier_8_io_x_pr; // @[package.scala 258:25]
  wire  entries_barrier_8_io_x_ppp; // @[package.scala 258:25]
  wire  entries_barrier_8_io_x_pal; // @[package.scala 258:25]
  wire  entries_barrier_8_io_x_paa; // @[package.scala 258:25]
  wire  entries_barrier_8_io_x_eff; // @[package.scala 258:25]
  wire  entries_barrier_8_io_x_c; // @[package.scala 258:25]
  wire [19:0] entries_barrier_8_io_y_ppn; // @[package.scala 258:25]
  wire  entries_barrier_8_io_y_u; // @[package.scala 258:25]
  wire  entries_barrier_8_io_y_ae; // @[package.scala 258:25]
  wire  entries_barrier_8_io_y_sw; // @[package.scala 258:25]
  wire  entries_barrier_8_io_y_sx; // @[package.scala 258:25]
  wire  entries_barrier_8_io_y_sr; // @[package.scala 258:25]
  wire  entries_barrier_8_io_y_pw; // @[package.scala 258:25]
  wire  entries_barrier_8_io_y_px; // @[package.scala 258:25]
  wire  entries_barrier_8_io_y_pr; // @[package.scala 258:25]
  wire  entries_barrier_8_io_y_ppp; // @[package.scala 258:25]
  wire  entries_barrier_8_io_y_pal; // @[package.scala 258:25]
  wire  entries_barrier_8_io_y_paa; // @[package.scala 258:25]
  wire  entries_barrier_8_io_y_eff; // @[package.scala 258:25]
  wire  entries_barrier_8_io_y_c; // @[package.scala 258:25]
  wire [29:0] entries_barrier_8_io_covSum; // @[package.scala 258:25]
  wire  entries_barrier_8_metaAssert; // @[package.scala 258:25]
  wire [19:0] entries_barrier_9_io_x_ppn; // @[package.scala 258:25]
  wire  entries_barrier_9_io_x_u; // @[package.scala 258:25]
  wire  entries_barrier_9_io_x_ae; // @[package.scala 258:25]
  wire  entries_barrier_9_io_x_sw; // @[package.scala 258:25]
  wire  entries_barrier_9_io_x_sx; // @[package.scala 258:25]
  wire  entries_barrier_9_io_x_sr; // @[package.scala 258:25]
  wire  entries_barrier_9_io_x_pw; // @[package.scala 258:25]
  wire  entries_barrier_9_io_x_px; // @[package.scala 258:25]
  wire  entries_barrier_9_io_x_pr; // @[package.scala 258:25]
  wire  entries_barrier_9_io_x_ppp; // @[package.scala 258:25]
  wire  entries_barrier_9_io_x_pal; // @[package.scala 258:25]
  wire  entries_barrier_9_io_x_paa; // @[package.scala 258:25]
  wire  entries_barrier_9_io_x_eff; // @[package.scala 258:25]
  wire  entries_barrier_9_io_x_c; // @[package.scala 258:25]
  wire [19:0] entries_barrier_9_io_y_ppn; // @[package.scala 258:25]
  wire  entries_barrier_9_io_y_u; // @[package.scala 258:25]
  wire  entries_barrier_9_io_y_ae; // @[package.scala 258:25]
  wire  entries_barrier_9_io_y_sw; // @[package.scala 258:25]
  wire  entries_barrier_9_io_y_sx; // @[package.scala 258:25]
  wire  entries_barrier_9_io_y_sr; // @[package.scala 258:25]
  wire  entries_barrier_9_io_y_pw; // @[package.scala 258:25]
  wire  entries_barrier_9_io_y_px; // @[package.scala 258:25]
  wire  entries_barrier_9_io_y_pr; // @[package.scala 258:25]
  wire  entries_barrier_9_io_y_ppp; // @[package.scala 258:25]
  wire  entries_barrier_9_io_y_pal; // @[package.scala 258:25]
  wire  entries_barrier_9_io_y_paa; // @[package.scala 258:25]
  wire  entries_barrier_9_io_y_eff; // @[package.scala 258:25]
  wire  entries_barrier_9_io_y_c; // @[package.scala 258:25]
  wire [29:0] entries_barrier_9_io_covSum; // @[package.scala 258:25]
  wire  entries_barrier_9_metaAssert; // @[package.scala 258:25]
  wire [19:0] entries_barrier_10_io_x_ppn; // @[package.scala 258:25]
  wire  entries_barrier_10_io_x_u; // @[package.scala 258:25]
  wire  entries_barrier_10_io_x_ae; // @[package.scala 258:25]
  wire  entries_barrier_10_io_x_sw; // @[package.scala 258:25]
  wire  entries_barrier_10_io_x_sx; // @[package.scala 258:25]
  wire  entries_barrier_10_io_x_sr; // @[package.scala 258:25]
  wire  entries_barrier_10_io_x_pw; // @[package.scala 258:25]
  wire  entries_barrier_10_io_x_px; // @[package.scala 258:25]
  wire  entries_barrier_10_io_x_pr; // @[package.scala 258:25]
  wire  entries_barrier_10_io_x_ppp; // @[package.scala 258:25]
  wire  entries_barrier_10_io_x_pal; // @[package.scala 258:25]
  wire  entries_barrier_10_io_x_paa; // @[package.scala 258:25]
  wire  entries_barrier_10_io_x_eff; // @[package.scala 258:25]
  wire  entries_barrier_10_io_x_c; // @[package.scala 258:25]
  wire [19:0] entries_barrier_10_io_y_ppn; // @[package.scala 258:25]
  wire  entries_barrier_10_io_y_u; // @[package.scala 258:25]
  wire  entries_barrier_10_io_y_ae; // @[package.scala 258:25]
  wire  entries_barrier_10_io_y_sw; // @[package.scala 258:25]
  wire  entries_barrier_10_io_y_sx; // @[package.scala 258:25]
  wire  entries_barrier_10_io_y_sr; // @[package.scala 258:25]
  wire  entries_barrier_10_io_y_pw; // @[package.scala 258:25]
  wire  entries_barrier_10_io_y_px; // @[package.scala 258:25]
  wire  entries_barrier_10_io_y_pr; // @[package.scala 258:25]
  wire  entries_barrier_10_io_y_ppp; // @[package.scala 258:25]
  wire  entries_barrier_10_io_y_pal; // @[package.scala 258:25]
  wire  entries_barrier_10_io_y_paa; // @[package.scala 258:25]
  wire  entries_barrier_10_io_y_eff; // @[package.scala 258:25]
  wire  entries_barrier_10_io_y_c; // @[package.scala 258:25]
  wire [29:0] entries_barrier_10_io_covSum; // @[package.scala 258:25]
  wire  entries_barrier_10_metaAssert; // @[package.scala 258:25]
  wire [19:0] entries_barrier_11_io_x_ppn; // @[package.scala 258:25]
  wire  entries_barrier_11_io_x_u; // @[package.scala 258:25]
  wire  entries_barrier_11_io_x_ae; // @[package.scala 258:25]
  wire  entries_barrier_11_io_x_sw; // @[package.scala 258:25]
  wire  entries_barrier_11_io_x_sx; // @[package.scala 258:25]
  wire  entries_barrier_11_io_x_sr; // @[package.scala 258:25]
  wire  entries_barrier_11_io_x_pw; // @[package.scala 258:25]
  wire  entries_barrier_11_io_x_px; // @[package.scala 258:25]
  wire  entries_barrier_11_io_x_pr; // @[package.scala 258:25]
  wire  entries_barrier_11_io_x_ppp; // @[package.scala 258:25]
  wire  entries_barrier_11_io_x_pal; // @[package.scala 258:25]
  wire  entries_barrier_11_io_x_paa; // @[package.scala 258:25]
  wire  entries_barrier_11_io_x_eff; // @[package.scala 258:25]
  wire  entries_barrier_11_io_x_c; // @[package.scala 258:25]
  wire [19:0] entries_barrier_11_io_y_ppn; // @[package.scala 258:25]
  wire  entries_barrier_11_io_y_u; // @[package.scala 258:25]
  wire  entries_barrier_11_io_y_ae; // @[package.scala 258:25]
  wire  entries_barrier_11_io_y_sw; // @[package.scala 258:25]
  wire  entries_barrier_11_io_y_sx; // @[package.scala 258:25]
  wire  entries_barrier_11_io_y_sr; // @[package.scala 258:25]
  wire  entries_barrier_11_io_y_pw; // @[package.scala 258:25]
  wire  entries_barrier_11_io_y_px; // @[package.scala 258:25]
  wire  entries_barrier_11_io_y_pr; // @[package.scala 258:25]
  wire  entries_barrier_11_io_y_ppp; // @[package.scala 258:25]
  wire  entries_barrier_11_io_y_pal; // @[package.scala 258:25]
  wire  entries_barrier_11_io_y_paa; // @[package.scala 258:25]
  wire  entries_barrier_11_io_y_eff; // @[package.scala 258:25]
  wire  entries_barrier_11_io_y_c; // @[package.scala 258:25]
  wire [29:0] entries_barrier_11_io_covSum; // @[package.scala 258:25]
  wire  entries_barrier_11_metaAssert; // @[package.scala 258:25]
  wire [19:0] entries_barrier_12_io_x_ppn; // @[package.scala 258:25]
  wire  entries_barrier_12_io_x_u; // @[package.scala 258:25]
  wire  entries_barrier_12_io_x_ae; // @[package.scala 258:25]
  wire  entries_barrier_12_io_x_sw; // @[package.scala 258:25]
  wire  entries_barrier_12_io_x_sx; // @[package.scala 258:25]
  wire  entries_barrier_12_io_x_sr; // @[package.scala 258:25]
  wire  entries_barrier_12_io_x_pw; // @[package.scala 258:25]
  wire  entries_barrier_12_io_x_px; // @[package.scala 258:25]
  wire  entries_barrier_12_io_x_pr; // @[package.scala 258:25]
  wire  entries_barrier_12_io_x_ppp; // @[package.scala 258:25]
  wire  entries_barrier_12_io_x_pal; // @[package.scala 258:25]
  wire  entries_barrier_12_io_x_paa; // @[package.scala 258:25]
  wire  entries_barrier_12_io_x_eff; // @[package.scala 258:25]
  wire  entries_barrier_12_io_x_c; // @[package.scala 258:25]
  wire [19:0] entries_barrier_12_io_y_ppn; // @[package.scala 258:25]
  wire  entries_barrier_12_io_y_u; // @[package.scala 258:25]
  wire  entries_barrier_12_io_y_ae; // @[package.scala 258:25]
  wire  entries_barrier_12_io_y_sw; // @[package.scala 258:25]
  wire  entries_barrier_12_io_y_sx; // @[package.scala 258:25]
  wire  entries_barrier_12_io_y_sr; // @[package.scala 258:25]
  wire  entries_barrier_12_io_y_pw; // @[package.scala 258:25]
  wire  entries_barrier_12_io_y_px; // @[package.scala 258:25]
  wire  entries_barrier_12_io_y_pr; // @[package.scala 258:25]
  wire  entries_barrier_12_io_y_ppp; // @[package.scala 258:25]
  wire  entries_barrier_12_io_y_pal; // @[package.scala 258:25]
  wire  entries_barrier_12_io_y_paa; // @[package.scala 258:25]
  wire  entries_barrier_12_io_y_eff; // @[package.scala 258:25]
  wire  entries_barrier_12_io_y_c; // @[package.scala 258:25]
  wire [29:0] entries_barrier_12_io_covSum; // @[package.scala 258:25]
  wire  entries_barrier_12_metaAssert; // @[package.scala 258:25]
  wire [26:0] vpn; // @[TLB.scala 162:30]
  reg [26:0] sectored_entries_0_0_tag; // @[TLB.scala 164:29]
  reg [31:0] _RAND_0;
  reg [34:0] sectored_entries_0_0_data_0; // @[TLB.scala 164:29]
  reg [63:0] _RAND_1;
  reg [34:0] sectored_entries_0_0_data_1; // @[TLB.scala 164:29]
  reg [63:0] _RAND_2;
  reg [34:0] sectored_entries_0_0_data_2; // @[TLB.scala 164:29]
  reg [63:0] _RAND_3;
  reg [34:0] sectored_entries_0_0_data_3; // @[TLB.scala 164:29]
  reg [63:0] _RAND_4;
  reg  sectored_entries_0_0_valid_0; // @[TLB.scala 164:29]
  reg [31:0] _RAND_5;
  reg  sectored_entries_0_0_valid_1; // @[TLB.scala 164:29]
  reg [31:0] _RAND_6;
  reg  sectored_entries_0_0_valid_2; // @[TLB.scala 164:29]
  reg [31:0] _RAND_7;
  reg  sectored_entries_0_0_valid_3; // @[TLB.scala 164:29]
  reg [31:0] _RAND_8;
  reg [26:0] sectored_entries_0_1_tag; // @[TLB.scala 164:29]
  reg [31:0] _RAND_9;
  reg [34:0] sectored_entries_0_1_data_0; // @[TLB.scala 164:29]
  reg [63:0] _RAND_10;
  reg [34:0] sectored_entries_0_1_data_1; // @[TLB.scala 164:29]
  reg [63:0] _RAND_11;
  reg [34:0] sectored_entries_0_1_data_2; // @[TLB.scala 164:29]
  reg [63:0] _RAND_12;
  reg [34:0] sectored_entries_0_1_data_3; // @[TLB.scala 164:29]
  reg [63:0] _RAND_13;
  reg  sectored_entries_0_1_valid_0; // @[TLB.scala 164:29]
  reg [31:0] _RAND_14;
  reg  sectored_entries_0_1_valid_1; // @[TLB.scala 164:29]
  reg [31:0] _RAND_15;
  reg  sectored_entries_0_1_valid_2; // @[TLB.scala 164:29]
  reg [31:0] _RAND_16;
  reg  sectored_entries_0_1_valid_3; // @[TLB.scala 164:29]
  reg [31:0] _RAND_17;
  reg [26:0] sectored_entries_0_2_tag; // @[TLB.scala 164:29]
  reg [31:0] _RAND_18;
  reg [34:0] sectored_entries_0_2_data_0; // @[TLB.scala 164:29]
  reg [63:0] _RAND_19;
  reg [34:0] sectored_entries_0_2_data_1; // @[TLB.scala 164:29]
  reg [63:0] _RAND_20;
  reg [34:0] sectored_entries_0_2_data_2; // @[TLB.scala 164:29]
  reg [63:0] _RAND_21;
  reg [34:0] sectored_entries_0_2_data_3; // @[TLB.scala 164:29]
  reg [63:0] _RAND_22;
  reg  sectored_entries_0_2_valid_0; // @[TLB.scala 164:29]
  reg [31:0] _RAND_23;
  reg  sectored_entries_0_2_valid_1; // @[TLB.scala 164:29]
  reg [31:0] _RAND_24;
  reg  sectored_entries_0_2_valid_2; // @[TLB.scala 164:29]
  reg [31:0] _RAND_25;
  reg  sectored_entries_0_2_valid_3; // @[TLB.scala 164:29]
  reg [31:0] _RAND_26;
  reg [26:0] sectored_entries_0_3_tag; // @[TLB.scala 164:29]
  reg [31:0] _RAND_27;
  reg [34:0] sectored_entries_0_3_data_0; // @[TLB.scala 164:29]
  reg [63:0] _RAND_28;
  reg [34:0] sectored_entries_0_3_data_1; // @[TLB.scala 164:29]
  reg [63:0] _RAND_29;
  reg [34:0] sectored_entries_0_3_data_2; // @[TLB.scala 164:29]
  reg [63:0] _RAND_30;
  reg [34:0] sectored_entries_0_3_data_3; // @[TLB.scala 164:29]
  reg [63:0] _RAND_31;
  reg  sectored_entries_0_3_valid_0; // @[TLB.scala 164:29]
  reg [31:0] _RAND_32;
  reg  sectored_entries_0_3_valid_1; // @[TLB.scala 164:29]
  reg [31:0] _RAND_33;
  reg  sectored_entries_0_3_valid_2; // @[TLB.scala 164:29]
  reg [31:0] _RAND_34;
  reg  sectored_entries_0_3_valid_3; // @[TLB.scala 164:29]
  reg [31:0] _RAND_35;
  reg [26:0] sectored_entries_0_4_tag; // @[TLB.scala 164:29]
  reg [31:0] _RAND_36;
  reg [34:0] sectored_entries_0_4_data_0; // @[TLB.scala 164:29]
  reg [63:0] _RAND_37;
  reg [34:0] sectored_entries_0_4_data_1; // @[TLB.scala 164:29]
  reg [63:0] _RAND_38;
  reg [34:0] sectored_entries_0_4_data_2; // @[TLB.scala 164:29]
  reg [63:0] _RAND_39;
  reg [34:0] sectored_entries_0_4_data_3; // @[TLB.scala 164:29]
  reg [63:0] _RAND_40;
  reg  sectored_entries_0_4_valid_0; // @[TLB.scala 164:29]
  reg [31:0] _RAND_41;
  reg  sectored_entries_0_4_valid_1; // @[TLB.scala 164:29]
  reg [31:0] _RAND_42;
  reg  sectored_entries_0_4_valid_2; // @[TLB.scala 164:29]
  reg [31:0] _RAND_43;
  reg  sectored_entries_0_4_valid_3; // @[TLB.scala 164:29]
  reg [31:0] _RAND_44;
  reg [26:0] sectored_entries_0_5_tag; // @[TLB.scala 164:29]
  reg [31:0] _RAND_45;
  reg [34:0] sectored_entries_0_5_data_0; // @[TLB.scala 164:29]
  reg [63:0] _RAND_46;
  reg [34:0] sectored_entries_0_5_data_1; // @[TLB.scala 164:29]
  reg [63:0] _RAND_47;
  reg [34:0] sectored_entries_0_5_data_2; // @[TLB.scala 164:29]
  reg [63:0] _RAND_48;
  reg [34:0] sectored_entries_0_5_data_3; // @[TLB.scala 164:29]
  reg [63:0] _RAND_49;
  reg  sectored_entries_0_5_valid_0; // @[TLB.scala 164:29]
  reg [31:0] _RAND_50;
  reg  sectored_entries_0_5_valid_1; // @[TLB.scala 164:29]
  reg [31:0] _RAND_51;
  reg  sectored_entries_0_5_valid_2; // @[TLB.scala 164:29]
  reg [31:0] _RAND_52;
  reg  sectored_entries_0_5_valid_3; // @[TLB.scala 164:29]
  reg [31:0] _RAND_53;
  reg [26:0] sectored_entries_0_6_tag; // @[TLB.scala 164:29]
  reg [31:0] _RAND_54;
  reg [34:0] sectored_entries_0_6_data_0; // @[TLB.scala 164:29]
  reg [63:0] _RAND_55;
  reg [34:0] sectored_entries_0_6_data_1; // @[TLB.scala 164:29]
  reg [63:0] _RAND_56;
  reg [34:0] sectored_entries_0_6_data_2; // @[TLB.scala 164:29]
  reg [63:0] _RAND_57;
  reg [34:0] sectored_entries_0_6_data_3; // @[TLB.scala 164:29]
  reg [63:0] _RAND_58;
  reg  sectored_entries_0_6_valid_0; // @[TLB.scala 164:29]
  reg [31:0] _RAND_59;
  reg  sectored_entries_0_6_valid_1; // @[TLB.scala 164:29]
  reg [31:0] _RAND_60;
  reg  sectored_entries_0_6_valid_2; // @[TLB.scala 164:29]
  reg [31:0] _RAND_61;
  reg  sectored_entries_0_6_valid_3; // @[TLB.scala 164:29]
  reg [31:0] _RAND_62;
  reg [26:0] sectored_entries_0_7_tag; // @[TLB.scala 164:29]
  reg [31:0] _RAND_63;
  reg [34:0] sectored_entries_0_7_data_0; // @[TLB.scala 164:29]
  reg [63:0] _RAND_64;
  reg [34:0] sectored_entries_0_7_data_1; // @[TLB.scala 164:29]
  reg [63:0] _RAND_65;
  reg [34:0] sectored_entries_0_7_data_2; // @[TLB.scala 164:29]
  reg [63:0] _RAND_66;
  reg [34:0] sectored_entries_0_7_data_3; // @[TLB.scala 164:29]
  reg [63:0] _RAND_67;
  reg  sectored_entries_0_7_valid_0; // @[TLB.scala 164:29]
  reg [31:0] _RAND_68;
  reg  sectored_entries_0_7_valid_1; // @[TLB.scala 164:29]
  reg [31:0] _RAND_69;
  reg  sectored_entries_0_7_valid_2; // @[TLB.scala 164:29]
  reg [31:0] _RAND_70;
  reg  sectored_entries_0_7_valid_3; // @[TLB.scala 164:29]
  reg [31:0] _RAND_71;
  reg [1:0] superpage_entries_0_level; // @[TLB.scala 165:30]
  reg [31:0] _RAND_72;
  reg [26:0] superpage_entries_0_tag; // @[TLB.scala 165:30]
  reg [31:0] _RAND_73;
  reg [34:0] superpage_entries_0_data_0; // @[TLB.scala 165:30]
  reg [63:0] _RAND_74;
  reg  superpage_entries_0_valid_0; // @[TLB.scala 165:30]
  reg [31:0] _RAND_75;
  reg [1:0] superpage_entries_1_level; // @[TLB.scala 165:30]
  reg [31:0] _RAND_76;
  reg [26:0] superpage_entries_1_tag; // @[TLB.scala 165:30]
  reg [31:0] _RAND_77;
  reg [34:0] superpage_entries_1_data_0; // @[TLB.scala 165:30]
  reg [63:0] _RAND_78;
  reg  superpage_entries_1_valid_0; // @[TLB.scala 165:30]
  reg [31:0] _RAND_79;
  reg [1:0] superpage_entries_2_level; // @[TLB.scala 165:30]
  reg [31:0] _RAND_80;
  reg [26:0] superpage_entries_2_tag; // @[TLB.scala 165:30]
  reg [31:0] _RAND_81;
  reg [34:0] superpage_entries_2_data_0; // @[TLB.scala 165:30]
  reg [63:0] _RAND_82;
  reg  superpage_entries_2_valid_0; // @[TLB.scala 165:30]
  reg [31:0] _RAND_83;
  reg [1:0] superpage_entries_3_level; // @[TLB.scala 165:30]
  reg [31:0] _RAND_84;
  reg [26:0] superpage_entries_3_tag; // @[TLB.scala 165:30]
  reg [31:0] _RAND_85;
  reg [34:0] superpage_entries_3_data_0; // @[TLB.scala 165:30]
  reg [63:0] _RAND_86;
  reg  superpage_entries_3_valid_0; // @[TLB.scala 165:30]
  reg [31:0] _RAND_87;
  reg [1:0] special_entry_level; // @[TLB.scala 166:56]
  reg [31:0] _RAND_88;
  reg [26:0] special_entry_tag; // @[TLB.scala 166:56]
  reg [31:0] _RAND_89;
  reg [34:0] special_entry_data_0; // @[TLB.scala 166:56]
  reg [63:0] _RAND_90;
  reg  special_entry_valid_0; // @[TLB.scala 166:56]
  reg [31:0] _RAND_91;
  reg [1:0] state; // @[TLB.scala 172:18]
  reg [31:0] _RAND_92;
  reg [26:0] r_refill_tag; // @[TLB.scala 173:25]
  reg [31:0] _RAND_93;
  reg [1:0] r_superpage_repl_addr; // @[TLB.scala 174:34]
  reg [31:0] _RAND_94;
  reg [2:0] r_sectored_repl_addr; // @[TLB.scala 175:33]
  reg [31:0] _RAND_95;
  reg [2:0] r_sectored_hit_addr; // @[TLB.scala 176:32]
  reg [31:0] _RAND_96;
  reg  r_sectored_hit; // @[TLB.scala 177:27]
  reg [31:0] _RAND_97;
  wire  priv_s; // @[TLB.scala 180:20]
  wire  priv_uses_vm; // @[TLB.scala 181:27]
  wire  _vm_enabled_T_2; // @[TLB.scala 182:83]
  wire  vm_enabled; // @[TLB.scala 182:99]
  wire [19:0] refill_ppn; // @[TLB.scala 185:44]
  wire  _invalidate_refill_T; // @[package.scala 15:47]
  wire  _invalidate_refill_T_1; // @[package.scala 15:47]
  wire  _invalidate_refill_T_2; // @[package.scala 72:59]
  wire  invalidate_refill; // @[TLB.scala 187:88]
  wire [1:0] mpu_ppn_hi; // @[TLB.scala 105:26]
  wire  mpu_ppn_ignore; // @[TLB.scala 107:28]
  wire [26:0] _mpu_ppn_T_17; // @[TLB.scala 108:28]
  wire [26:0] _GEN_919; // @[TLB.scala 108:47]
  wire [26:0] _mpu_ppn_T_18; // @[TLB.scala 108:47]
  wire [8:0] mpu_ppn_lo; // @[TLB.scala 108:58]
  wire  mpu_ppn_ignore_1; // @[TLB.scala 107:28]
  wire [26:0] _mpu_ppn_T_19; // @[TLB.scala 108:28]
  wire [26:0] _mpu_ppn_T_20; // @[TLB.scala 108:47]
  wire [8:0] mpu_ppn_lo_1; // @[TLB.scala 108:58]
  wire [19:0] _mpu_ppn_T_21; // @[Cat.scala 30:58]
  wire [27:0] _mpu_ppn_T_23; // @[TLB.scala 189:20]
  wire [27:0] mpu_ppn; // @[TLB.scala 188:20]
  wire [11:0] mpu_physaddr_lo; // @[TLB.scala 190:52]
  wire [39:0] mpu_physaddr; // @[Cat.scala 30:58]
  wire  _mpu_priv_T; // @[TLB.scala 191:56]
  wire [2:0] _mpu_priv_T_2; // @[Cat.scala 30:58]
  wire [2:0] mpu_priv; // @[TLB.scala 191:27]
  wire [39:0] _legal_address_T; // @[Parameters.scala 137:31]
  wire [40:0] _legal_address_T_1; // @[Parameters.scala 137:49]
  wire [40:0] _legal_address_T_3; // @[Parameters.scala 137:52]
  wire  _legal_address_T_4; // @[Parameters.scala 137:67]
  wire [39:0] _legal_address_T_5; // @[Parameters.scala 137:31]
  wire [40:0] _legal_address_T_6; // @[Parameters.scala 137:49]
  wire [40:0] _legal_address_T_8; // @[Parameters.scala 137:52]
  wire  _legal_address_T_9; // @[Parameters.scala 137:67]
  wire [39:0] _legal_address_T_10; // @[Parameters.scala 137:31]
  wire [40:0] _legal_address_T_11; // @[Parameters.scala 137:49]
  wire [40:0] _legal_address_T_13; // @[Parameters.scala 137:52]
  wire  _legal_address_T_14; // @[Parameters.scala 137:67]
  wire [40:0] _legal_address_T_16; // @[Parameters.scala 137:49]
  wire [40:0] _legal_address_T_18; // @[Parameters.scala 137:52]
  wire  _legal_address_T_19; // @[Parameters.scala 137:67]
  wire [39:0] _legal_address_T_20; // @[Parameters.scala 137:31]
  wire [40:0] _legal_address_T_21; // @[Parameters.scala 137:49]
  wire [40:0] _legal_address_T_23; // @[Parameters.scala 137:52]
  wire  _legal_address_T_24; // @[Parameters.scala 137:67]
  wire [39:0] _legal_address_T_25; // @[Parameters.scala 137:31]
  wire [40:0] _legal_address_T_26; // @[Parameters.scala 137:49]
  wire [40:0] _legal_address_T_28; // @[Parameters.scala 137:52]
  wire  _legal_address_T_29; // @[Parameters.scala 137:67]
  wire [39:0] _legal_address_T_30; // @[Parameters.scala 137:31]
  wire [40:0] _legal_address_T_31; // @[Parameters.scala 137:49]
  wire [40:0] _legal_address_T_33; // @[Parameters.scala 137:52]
  wire  _legal_address_T_34; // @[Parameters.scala 137:67]
  wire  _legal_address_T_35; // @[TLB.scala 197:67]
  wire  _legal_address_T_36; // @[TLB.scala 197:67]
  wire  _legal_address_T_37; // @[TLB.scala 197:67]
  wire  _legal_address_T_38; // @[TLB.scala 197:67]
  wire  _legal_address_T_39; // @[TLB.scala 197:67]
  wire  legal_address; // @[TLB.scala 197:67]
  wire [40:0] _cacheable_T_8; // @[Parameters.scala 137:52]
  wire  _cacheable_T_9; // @[Parameters.scala 137:67]
  wire  cacheable; // @[TLB.scala 199:19]
  wire [39:0] _homogeneous_T_54; // @[Parameters.scala 137:31]
  wire [40:0] _homogeneous_T_55; // @[Parameters.scala 137:49]
  wire [40:0] _homogeneous_T_57; // @[Parameters.scala 137:52]
  wire  _homogeneous_T_58; // @[Parameters.scala 137:67]
  wire [40:0] _homogeneous_T_71; // @[Parameters.scala 137:52]
  wire  _homogeneous_T_72; // @[Parameters.scala 137:67]
  wire  _homogeneous_T_79; // @[TLBPermissions.scala 83:66]
  wire  _deny_access_to_debug_T; // @[TLB.scala 202:39]
  wire  deny_access_to_debug; // @[TLB.scala 202:48]
  wire  _prot_r_T_7; // @[TLB.scala 203:41]
  wire  prot_r; // @[TLB.scala 203:66]
  wire [39:0] _prot_w_T_10; // @[Parameters.scala 137:31]
  wire [40:0] _prot_w_T_11; // @[Parameters.scala 137:49]
  wire [40:0] _prot_w_T_13; // @[Parameters.scala 137:52]
  wire  _prot_w_T_14; // @[Parameters.scala 137:67]
  wire [40:0] _prot_w_T_18; // @[Parameters.scala 137:52]
  wire  _prot_w_T_19; // @[Parameters.scala 137:67]
  wire  _prot_w_T_21; // @[Parameters.scala 615:89]
  wire  _prot_w_T_22; // @[Parameters.scala 615:89]
  wire  _prot_w_T_31; // @[TLB.scala 199:19]
  wire  _prot_w_T_33; // @[TLB.scala 204:45]
  wire  prot_w; // @[TLB.scala 204:70]
  wire  prot_al; // @[TLB.scala 199:19]
  wire [40:0] _prot_x_T_3; // @[Parameters.scala 137:52]
  wire  _prot_x_T_4; // @[Parameters.scala 137:67]
  wire  _prot_x_T_15; // @[Parameters.scala 615:89]
  wire  _prot_x_T_16; // @[Parameters.scala 615:89]
  wire  _prot_x_T_31; // @[TLB.scala 199:19]
  wire  _prot_x_T_33; // @[TLB.scala 208:40]
  wire  prot_x; // @[TLB.scala 208:65]
  wire [40:0] _prot_eff_T_20; // @[Parameters.scala 137:52]
  wire  _prot_eff_T_21; // @[Parameters.scala 137:67]
  wire [40:0] _prot_eff_T_25; // @[Parameters.scala 137:52]
  wire  _prot_eff_T_26; // @[Parameters.scala 137:67]
  wire  _prot_eff_T_37; // @[Parameters.scala 615:89]
  wire  _prot_eff_T_38; // @[Parameters.scala 615:89]
  wire  _prot_eff_T_39; // @[Parameters.scala 615:89]
  wire  prot_eff; // @[TLB.scala 199:19]
  wire  _sector_hits_T; // @[package.scala 72:59]
  wire  _sector_hits_T_1; // @[package.scala 72:59]
  wire  _sector_hits_T_2; // @[package.scala 72:59]
  wire [26:0] _sector_hits_T_3; // @[TLB.scala 88:41]
  wire  _sector_hits_T_5; // @[TLB.scala 88:66]
  wire  sector_hits_0; // @[TLB.scala 87:40]
  wire  _sector_hits_T_6; // @[package.scala 72:59]
  wire  _sector_hits_T_7; // @[package.scala 72:59]
  wire  _sector_hits_T_8; // @[package.scala 72:59]
  wire [26:0] _sector_hits_T_9; // @[TLB.scala 88:41]
  wire  _sector_hits_T_11; // @[TLB.scala 88:66]
  wire  sector_hits_1; // @[TLB.scala 87:40]
  wire  _sector_hits_T_12; // @[package.scala 72:59]
  wire  _sector_hits_T_13; // @[package.scala 72:59]
  wire  _sector_hits_T_14; // @[package.scala 72:59]
  wire [26:0] _sector_hits_T_15; // @[TLB.scala 88:41]
  wire  _sector_hits_T_17; // @[TLB.scala 88:66]
  wire  sector_hits_2; // @[TLB.scala 87:40]
  wire  _sector_hits_T_18; // @[package.scala 72:59]
  wire  _sector_hits_T_19; // @[package.scala 72:59]
  wire  _sector_hits_T_20; // @[package.scala 72:59]
  wire [26:0] _sector_hits_T_21; // @[TLB.scala 88:41]
  wire  _sector_hits_T_23; // @[TLB.scala 88:66]
  wire  sector_hits_3; // @[TLB.scala 87:40]
  wire  _sector_hits_T_24; // @[package.scala 72:59]
  wire  _sector_hits_T_25; // @[package.scala 72:59]
  wire  _sector_hits_T_26; // @[package.scala 72:59]
  wire [26:0] _sector_hits_T_27; // @[TLB.scala 88:41]
  wire  _sector_hits_T_29; // @[TLB.scala 88:66]
  wire  sector_hits_4; // @[TLB.scala 87:40]
  wire  _sector_hits_T_30; // @[package.scala 72:59]
  wire  _sector_hits_T_31; // @[package.scala 72:59]
  wire  _sector_hits_T_32; // @[package.scala 72:59]
  wire [26:0] _sector_hits_T_33; // @[TLB.scala 88:41]
  wire  _sector_hits_T_35; // @[TLB.scala 88:66]
  wire  sector_hits_5; // @[TLB.scala 87:40]
  wire  _sector_hits_T_36; // @[package.scala 72:59]
  wire  _sector_hits_T_37; // @[package.scala 72:59]
  wire  _sector_hits_T_38; // @[package.scala 72:59]
  wire [26:0] _sector_hits_T_39; // @[TLB.scala 88:41]
  wire  _sector_hits_T_41; // @[TLB.scala 88:66]
  wire  sector_hits_6; // @[TLB.scala 87:40]
  wire  _sector_hits_T_42; // @[package.scala 72:59]
  wire  _sector_hits_T_43; // @[package.scala 72:59]
  wire  _sector_hits_T_44; // @[package.scala 72:59]
  wire [26:0] _sector_hits_T_45; // @[TLB.scala 88:41]
  wire  _sector_hits_T_47; // @[TLB.scala 88:66]
  wire  sector_hits_7; // @[TLB.scala 87:40]
  wire  _superpage_hits_T_2; // @[TLB.scala 95:77]
  wire  _superpage_hits_T_4; // @[TLB.scala 95:29]
  wire  superpage_hits_ignore_1; // @[TLB.scala 94:28]
  wire  _superpage_hits_T_7; // @[TLB.scala 95:77]
  wire  _superpage_hits_T_8; // @[TLB.scala 95:40]
  wire  superpage_hits_0; // @[TLB.scala 95:29]
  wire  _superpage_hits_T_16; // @[TLB.scala 95:77]
  wire  _superpage_hits_T_18; // @[TLB.scala 95:29]
  wire  superpage_hits_ignore_4; // @[TLB.scala 94:28]
  wire  _superpage_hits_T_21; // @[TLB.scala 95:77]
  wire  _superpage_hits_T_22; // @[TLB.scala 95:40]
  wire  superpage_hits_1; // @[TLB.scala 95:29]
  wire  _superpage_hits_T_30; // @[TLB.scala 95:77]
  wire  _superpage_hits_T_32; // @[TLB.scala 95:29]
  wire  superpage_hits_ignore_7; // @[TLB.scala 94:28]
  wire  _superpage_hits_T_35; // @[TLB.scala 95:77]
  wire  _superpage_hits_T_36; // @[TLB.scala 95:40]
  wire  superpage_hits_2; // @[TLB.scala 95:29]
  wire  _superpage_hits_T_44; // @[TLB.scala 95:77]
  wire  _superpage_hits_T_46; // @[TLB.scala 95:29]
  wire  superpage_hits_ignore_10; // @[TLB.scala 94:28]
  wire  _superpage_hits_T_49; // @[TLB.scala 95:77]
  wire  _superpage_hits_T_50; // @[TLB.scala 95:40]
  wire  superpage_hits_3; // @[TLB.scala 95:29]
  wire [1:0] hitsVec_idx; // @[package.scala 154:13]
  wire  _GEN_1; // @[TLB.scala 100:18]
  wire  _GEN_2; // @[TLB.scala 100:18]
  wire  _GEN_3; // @[TLB.scala 100:18]
  wire  _hitsVec_T_3; // @[TLB.scala 100:18]
  wire  hitsVec_0; // @[TLB.scala 213:44]
  wire  _GEN_5; // @[TLB.scala 100:18]
  wire  _GEN_6; // @[TLB.scala 100:18]
  wire  _GEN_7; // @[TLB.scala 100:18]
  wire  _hitsVec_T_7; // @[TLB.scala 100:18]
  wire  hitsVec_1; // @[TLB.scala 213:44]
  wire  _GEN_9; // @[TLB.scala 100:18]
  wire  _GEN_10; // @[TLB.scala 100:18]
  wire  _GEN_11; // @[TLB.scala 100:18]
  wire  _hitsVec_T_11; // @[TLB.scala 100:18]
  wire  hitsVec_2; // @[TLB.scala 213:44]
  wire  _GEN_13; // @[TLB.scala 100:18]
  wire  _GEN_14; // @[TLB.scala 100:18]
  wire  _GEN_15; // @[TLB.scala 100:18]
  wire  _hitsVec_T_15; // @[TLB.scala 100:18]
  wire  hitsVec_3; // @[TLB.scala 213:44]
  wire  _GEN_17; // @[TLB.scala 100:18]
  wire  _GEN_18; // @[TLB.scala 100:18]
  wire  _GEN_19; // @[TLB.scala 100:18]
  wire  _hitsVec_T_19; // @[TLB.scala 100:18]
  wire  hitsVec_4; // @[TLB.scala 213:44]
  wire  _GEN_21; // @[TLB.scala 100:18]
  wire  _GEN_22; // @[TLB.scala 100:18]
  wire  _GEN_23; // @[TLB.scala 100:18]
  wire  _hitsVec_T_23; // @[TLB.scala 100:18]
  wire  hitsVec_5; // @[TLB.scala 213:44]
  wire  _GEN_25; // @[TLB.scala 100:18]
  wire  _GEN_26; // @[TLB.scala 100:18]
  wire  _GEN_27; // @[TLB.scala 100:18]
  wire  _hitsVec_T_27; // @[TLB.scala 100:18]
  wire  hitsVec_6; // @[TLB.scala 213:44]
  wire  _GEN_29; // @[TLB.scala 100:18]
  wire  _GEN_30; // @[TLB.scala 100:18]
  wire  _GEN_31; // @[TLB.scala 100:18]
  wire  _hitsVec_T_31; // @[TLB.scala 100:18]
  wire  hitsVec_7; // @[TLB.scala 213:44]
  wire  hitsVec_8; // @[TLB.scala 213:44]
  wire  hitsVec_9; // @[TLB.scala 213:44]
  wire  hitsVec_10; // @[TLB.scala 213:44]
  wire  hitsVec_11; // @[TLB.scala 213:44]
  wire  _hitsVec_T_94; // @[TLB.scala 95:77]
  wire  _hitsVec_T_96; // @[TLB.scala 95:29]
  wire  _hitsVec_T_99; // @[TLB.scala 95:77]
  wire  _hitsVec_T_100; // @[TLB.scala 95:40]
  wire  _hitsVec_T_101; // @[TLB.scala 95:29]
  wire  _hitsVec_T_104; // @[TLB.scala 95:77]
  wire  _hitsVec_T_105; // @[TLB.scala 95:40]
  wire  _hitsVec_T_106; // @[TLB.scala 95:29]
  wire  hitsVec_12; // @[TLB.scala 213:44]
  wire [5:0] real_hits_lo; // @[Cat.scala 30:58]
  wire [12:0] real_hits; // @[Cat.scala 30:58]
  wire  hits_hi; // @[TLB.scala 215:18]
  wire [13:0] hits; // @[Cat.scala 30:58]
  wire  newEntry_g; // @[TLB.scala 224:25]
  wire  _newEntry_sr_T_1; // @[PTW.scala 73:44]
  wire  _newEntry_sr_T_2; // @[PTW.scala 73:38]
  wire  _newEntry_sr_T_3; // @[PTW.scala 73:32]
  wire  _newEntry_sr_T_4; // @[PTW.scala 73:52]
  wire  newEntry_sr; // @[PTW.scala 77:35]
  wire  _newEntry_sw_T_5; // @[PTW.scala 78:35]
  wire  newEntry_sw; // @[PTW.scala 78:40]
  wire  newEntry_sx; // @[PTW.scala 79:35]
  wire [7:0] special_entry_data_0_lo; // @[TLB.scala 122:24]
  wire [34:0] _special_entry_data_0_T; // @[TLB.scala 122:24]
  wire  _GEN_32; // @[TLB.scala 241:34]
  wire  _T_2; // @[TLB.scala 243:40]
  wire  _T_3; // @[TLB.scala 244:82]
  wire  _GEN_35; // @[TLB.scala 244:89]
  wire  _T_4; // @[TLB.scala 244:82]
  wire  _GEN_39; // @[TLB.scala 244:89]
  wire  _T_5; // @[TLB.scala 244:82]
  wire  _GEN_43; // @[TLB.scala 244:89]
  wire  _T_6; // @[TLB.scala 244:82]
  wire  _GEN_47; // @[TLB.scala 244:89]
  wire [2:0] waddr; // @[TLB.scala 250:22]
  wire  _T_7; // @[TLB.scala 251:75]
  wire  _GEN_49; // @[TLB.scala 252:32]
  wire  _GEN_50; // @[TLB.scala 252:32]
  wire  _GEN_51; // @[TLB.scala 252:32]
  wire  _GEN_52; // @[TLB.scala 252:32]
  wire [1:0] idx; // @[package.scala 154:13]
  wire  _GEN_921; // @[TLB.scala 121:16]
  wire  _GEN_53; // @[TLB.scala 121:16]
  wire  _GEN_922; // @[TLB.scala 121:16]
  wire  _GEN_54; // @[TLB.scala 121:16]
  wire  _GEN_923; // @[TLB.scala 121:16]
  wire  _GEN_55; // @[TLB.scala 121:16]
  wire  _GEN_924; // @[TLB.scala 121:16]
  wire  _GEN_56; // @[TLB.scala 121:16]
  wire  _GEN_61; // @[TLB.scala 254:34]
  wire  _GEN_62; // @[TLB.scala 254:34]
  wire  _GEN_63; // @[TLB.scala 254:34]
  wire  _GEN_64; // @[TLB.scala 254:34]
  wire  _GEN_65; // @[TLB.scala 251:82]
  wire  _GEN_66; // @[TLB.scala 251:82]
  wire  _GEN_67; // @[TLB.scala 251:82]
  wire  _GEN_68; // @[TLB.scala 251:82]
  wire  _T_9; // @[TLB.scala 251:75]
  wire  _GEN_75; // @[TLB.scala 252:32]
  wire  _GEN_76; // @[TLB.scala 252:32]
  wire  _GEN_77; // @[TLB.scala 252:32]
  wire  _GEN_78; // @[TLB.scala 252:32]
  wire  _GEN_79; // @[TLB.scala 121:16]
  wire  _GEN_80; // @[TLB.scala 121:16]
  wire  _GEN_81; // @[TLB.scala 121:16]
  wire  _GEN_82; // @[TLB.scala 121:16]
  wire  _GEN_87; // @[TLB.scala 254:34]
  wire  _GEN_88; // @[TLB.scala 254:34]
  wire  _GEN_89; // @[TLB.scala 254:34]
  wire  _GEN_90; // @[TLB.scala 254:34]
  wire  _GEN_91; // @[TLB.scala 251:82]
  wire  _GEN_92; // @[TLB.scala 251:82]
  wire  _GEN_93; // @[TLB.scala 251:82]
  wire  _GEN_94; // @[TLB.scala 251:82]
  wire  _T_11; // @[TLB.scala 251:75]
  wire  _GEN_101; // @[TLB.scala 252:32]
  wire  _GEN_102; // @[TLB.scala 252:32]
  wire  _GEN_103; // @[TLB.scala 252:32]
  wire  _GEN_104; // @[TLB.scala 252:32]
  wire  _GEN_105; // @[TLB.scala 121:16]
  wire  _GEN_106; // @[TLB.scala 121:16]
  wire  _GEN_107; // @[TLB.scala 121:16]
  wire  _GEN_108; // @[TLB.scala 121:16]
  wire  _GEN_113; // @[TLB.scala 254:34]
  wire  _GEN_114; // @[TLB.scala 254:34]
  wire  _GEN_115; // @[TLB.scala 254:34]
  wire  _GEN_116; // @[TLB.scala 254:34]
  wire  _GEN_117; // @[TLB.scala 251:82]
  wire  _GEN_118; // @[TLB.scala 251:82]
  wire  _GEN_119; // @[TLB.scala 251:82]
  wire  _GEN_120; // @[TLB.scala 251:82]
  wire  _T_13; // @[TLB.scala 251:75]
  wire  _GEN_127; // @[TLB.scala 252:32]
  wire  _GEN_128; // @[TLB.scala 252:32]
  wire  _GEN_129; // @[TLB.scala 252:32]
  wire  _GEN_130; // @[TLB.scala 252:32]
  wire  _GEN_131; // @[TLB.scala 121:16]
  wire  _GEN_132; // @[TLB.scala 121:16]
  wire  _GEN_133; // @[TLB.scala 121:16]
  wire  _GEN_134; // @[TLB.scala 121:16]
  wire  _GEN_139; // @[TLB.scala 254:34]
  wire  _GEN_140; // @[TLB.scala 254:34]
  wire  _GEN_141; // @[TLB.scala 254:34]
  wire  _GEN_142; // @[TLB.scala 254:34]
  wire  _GEN_143; // @[TLB.scala 251:82]
  wire  _GEN_144; // @[TLB.scala 251:82]
  wire  _GEN_145; // @[TLB.scala 251:82]
  wire  _GEN_146; // @[TLB.scala 251:82]
  wire  _T_15; // @[TLB.scala 251:75]
  wire  _GEN_153; // @[TLB.scala 252:32]
  wire  _GEN_154; // @[TLB.scala 252:32]
  wire  _GEN_155; // @[TLB.scala 252:32]
  wire  _GEN_156; // @[TLB.scala 252:32]
  wire  _GEN_157; // @[TLB.scala 121:16]
  wire  _GEN_158; // @[TLB.scala 121:16]
  wire  _GEN_159; // @[TLB.scala 121:16]
  wire  _GEN_160; // @[TLB.scala 121:16]
  wire  _GEN_165; // @[TLB.scala 254:34]
  wire  _GEN_166; // @[TLB.scala 254:34]
  wire  _GEN_167; // @[TLB.scala 254:34]
  wire  _GEN_168; // @[TLB.scala 254:34]
  wire  _GEN_169; // @[TLB.scala 251:82]
  wire  _GEN_170; // @[TLB.scala 251:82]
  wire  _GEN_171; // @[TLB.scala 251:82]
  wire  _GEN_172; // @[TLB.scala 251:82]
  wire  _T_17; // @[TLB.scala 251:75]
  wire  _GEN_179; // @[TLB.scala 252:32]
  wire  _GEN_180; // @[TLB.scala 252:32]
  wire  _GEN_181; // @[TLB.scala 252:32]
  wire  _GEN_182; // @[TLB.scala 252:32]
  wire  _GEN_183; // @[TLB.scala 121:16]
  wire  _GEN_184; // @[TLB.scala 121:16]
  wire  _GEN_185; // @[TLB.scala 121:16]
  wire  _GEN_186; // @[TLB.scala 121:16]
  wire  _GEN_191; // @[TLB.scala 254:34]
  wire  _GEN_192; // @[TLB.scala 254:34]
  wire  _GEN_193; // @[TLB.scala 254:34]
  wire  _GEN_194; // @[TLB.scala 254:34]
  wire  _GEN_195; // @[TLB.scala 251:82]
  wire  _GEN_196; // @[TLB.scala 251:82]
  wire  _GEN_197; // @[TLB.scala 251:82]
  wire  _GEN_198; // @[TLB.scala 251:82]
  wire  _T_19; // @[TLB.scala 251:75]
  wire  _GEN_205; // @[TLB.scala 252:32]
  wire  _GEN_206; // @[TLB.scala 252:32]
  wire  _GEN_207; // @[TLB.scala 252:32]
  wire  _GEN_208; // @[TLB.scala 252:32]
  wire  _GEN_209; // @[TLB.scala 121:16]
  wire  _GEN_210; // @[TLB.scala 121:16]
  wire  _GEN_211; // @[TLB.scala 121:16]
  wire  _GEN_212; // @[TLB.scala 121:16]
  wire  _GEN_217; // @[TLB.scala 254:34]
  wire  _GEN_218; // @[TLB.scala 254:34]
  wire  _GEN_219; // @[TLB.scala 254:34]
  wire  _GEN_220; // @[TLB.scala 254:34]
  wire  _GEN_221; // @[TLB.scala 251:82]
  wire  _GEN_222; // @[TLB.scala 251:82]
  wire  _GEN_223; // @[TLB.scala 251:82]
  wire  _GEN_224; // @[TLB.scala 251:82]
  wire  _T_21; // @[TLB.scala 251:75]
  wire  _GEN_231; // @[TLB.scala 252:32]
  wire  _GEN_232; // @[TLB.scala 252:32]
  wire  _GEN_233; // @[TLB.scala 252:32]
  wire  _GEN_234; // @[TLB.scala 252:32]
  wire  _GEN_235; // @[TLB.scala 121:16]
  wire  _GEN_236; // @[TLB.scala 121:16]
  wire  _GEN_237; // @[TLB.scala 121:16]
  wire  _GEN_238; // @[TLB.scala 121:16]
  wire  _GEN_243; // @[TLB.scala 254:34]
  wire  _GEN_244; // @[TLB.scala 254:34]
  wire  _GEN_245; // @[TLB.scala 254:34]
  wire  _GEN_246; // @[TLB.scala 254:34]
  wire  _GEN_247; // @[TLB.scala 251:82]
  wire  _GEN_248; // @[TLB.scala 251:82]
  wire  _GEN_249; // @[TLB.scala 251:82]
  wire  _GEN_250; // @[TLB.scala 251:82]
  wire  _GEN_259; // @[TLB.scala 243:54]
  wire  _GEN_263; // @[TLB.scala 243:54]
  wire  _GEN_267; // @[TLB.scala 243:54]
  wire  _GEN_271; // @[TLB.scala 243:54]
  wire  _GEN_273; // @[TLB.scala 243:54]
  wire  _GEN_274; // @[TLB.scala 243:54]
  wire  _GEN_275; // @[TLB.scala 243:54]
  wire  _GEN_276; // @[TLB.scala 243:54]
  wire  _GEN_283; // @[TLB.scala 243:54]
  wire  _GEN_284; // @[TLB.scala 243:54]
  wire  _GEN_285; // @[TLB.scala 243:54]
  wire  _GEN_286; // @[TLB.scala 243:54]
  wire  _GEN_293; // @[TLB.scala 243:54]
  wire  _GEN_294; // @[TLB.scala 243:54]
  wire  _GEN_295; // @[TLB.scala 243:54]
  wire  _GEN_296; // @[TLB.scala 243:54]
  wire  _GEN_303; // @[TLB.scala 243:54]
  wire  _GEN_304; // @[TLB.scala 243:54]
  wire  _GEN_305; // @[TLB.scala 243:54]
  wire  _GEN_306; // @[TLB.scala 243:54]
  wire  _GEN_313; // @[TLB.scala 243:54]
  wire  _GEN_314; // @[TLB.scala 243:54]
  wire  _GEN_315; // @[TLB.scala 243:54]
  wire  _GEN_316; // @[TLB.scala 243:54]
  wire  _GEN_323; // @[TLB.scala 243:54]
  wire  _GEN_324; // @[TLB.scala 243:54]
  wire  _GEN_325; // @[TLB.scala 243:54]
  wire  _GEN_326; // @[TLB.scala 243:54]
  wire  _GEN_333; // @[TLB.scala 243:54]
  wire  _GEN_334; // @[TLB.scala 243:54]
  wire  _GEN_335; // @[TLB.scala 243:54]
  wire  _GEN_336; // @[TLB.scala 243:54]
  wire  _GEN_343; // @[TLB.scala 243:54]
  wire  _GEN_344; // @[TLB.scala 243:54]
  wire  _GEN_345; // @[TLB.scala 243:54]
  wire  _GEN_346; // @[TLB.scala 243:54]
  wire  _GEN_355; // @[TLB.scala 238:68]
  wire  _GEN_359; // @[TLB.scala 238:68]
  wire  _GEN_363; // @[TLB.scala 238:68]
  wire  _GEN_367; // @[TLB.scala 238:68]
  wire  _GEN_371; // @[TLB.scala 238:68]
  wire  _GEN_373; // @[TLB.scala 238:68]
  wire  _GEN_374; // @[TLB.scala 238:68]
  wire  _GEN_375; // @[TLB.scala 238:68]
  wire  _GEN_376; // @[TLB.scala 238:68]
  wire  _GEN_383; // @[TLB.scala 238:68]
  wire  _GEN_384; // @[TLB.scala 238:68]
  wire  _GEN_385; // @[TLB.scala 238:68]
  wire  _GEN_386; // @[TLB.scala 238:68]
  wire  _GEN_393; // @[TLB.scala 238:68]
  wire  _GEN_394; // @[TLB.scala 238:68]
  wire  _GEN_395; // @[TLB.scala 238:68]
  wire  _GEN_396; // @[TLB.scala 238:68]
  wire  _GEN_403; // @[TLB.scala 238:68]
  wire  _GEN_404; // @[TLB.scala 238:68]
  wire  _GEN_405; // @[TLB.scala 238:68]
  wire  _GEN_406; // @[TLB.scala 238:68]
  wire  _GEN_413; // @[TLB.scala 238:68]
  wire  _GEN_414; // @[TLB.scala 238:68]
  wire  _GEN_415; // @[TLB.scala 238:68]
  wire  _GEN_416; // @[TLB.scala 238:68]
  wire  _GEN_423; // @[TLB.scala 238:68]
  wire  _GEN_424; // @[TLB.scala 238:68]
  wire  _GEN_425; // @[TLB.scala 238:68]
  wire  _GEN_426; // @[TLB.scala 238:68]
  wire  _GEN_433; // @[TLB.scala 238:68]
  wire  _GEN_434; // @[TLB.scala 238:68]
  wire  _GEN_435; // @[TLB.scala 238:68]
  wire  _GEN_436; // @[TLB.scala 238:68]
  wire  _GEN_443; // @[TLB.scala 238:68]
  wire  _GEN_444; // @[TLB.scala 238:68]
  wire  _GEN_445; // @[TLB.scala 238:68]
  wire  _GEN_446; // @[TLB.scala 238:68]
  wire  _GEN_455; // @[TLB.scala 218:20]
  wire  _GEN_459; // @[TLB.scala 218:20]
  wire  _GEN_463; // @[TLB.scala 218:20]
  wire  _GEN_467; // @[TLB.scala 218:20]
  wire  _GEN_471; // @[TLB.scala 218:20]
  wire  _GEN_473; // @[TLB.scala 218:20]
  wire  _GEN_474; // @[TLB.scala 218:20]
  wire  _GEN_475; // @[TLB.scala 218:20]
  wire  _GEN_476; // @[TLB.scala 218:20]
  wire  _GEN_483; // @[TLB.scala 218:20]
  wire  _GEN_484; // @[TLB.scala 218:20]
  wire  _GEN_485; // @[TLB.scala 218:20]
  wire  _GEN_486; // @[TLB.scala 218:20]
  wire  _GEN_493; // @[TLB.scala 218:20]
  wire  _GEN_494; // @[TLB.scala 218:20]
  wire  _GEN_495; // @[TLB.scala 218:20]
  wire  _GEN_496; // @[TLB.scala 218:20]
  wire  _GEN_503; // @[TLB.scala 218:20]
  wire  _GEN_504; // @[TLB.scala 218:20]
  wire  _GEN_505; // @[TLB.scala 218:20]
  wire  _GEN_506; // @[TLB.scala 218:20]
  wire  _GEN_513; // @[TLB.scala 218:20]
  wire  _GEN_514; // @[TLB.scala 218:20]
  wire  _GEN_515; // @[TLB.scala 218:20]
  wire  _GEN_516; // @[TLB.scala 218:20]
  wire  _GEN_523; // @[TLB.scala 218:20]
  wire  _GEN_524; // @[TLB.scala 218:20]
  wire  _GEN_525; // @[TLB.scala 218:20]
  wire  _GEN_526; // @[TLB.scala 218:20]
  wire  _GEN_533; // @[TLB.scala 218:20]
  wire  _GEN_534; // @[TLB.scala 218:20]
  wire  _GEN_535; // @[TLB.scala 218:20]
  wire  _GEN_536; // @[TLB.scala 218:20]
  wire  _GEN_543; // @[TLB.scala 218:20]
  wire  _GEN_544; // @[TLB.scala 218:20]
  wire  _GEN_545; // @[TLB.scala 218:20]
  wire  _GEN_546; // @[TLB.scala 218:20]
  wire [34:0] _GEN_554;
  wire [34:0] _GEN_555;
  wire [34:0] _GEN_556;
  wire [34:0] _GEN_558;
  wire [34:0] _GEN_559;
  wire [34:0] _GEN_560;
  wire [34:0] _GEN_562;
  wire [34:0] _GEN_563;
  wire [34:0] _GEN_564;
  wire [34:0] _GEN_566;
  wire [34:0] _GEN_567;
  wire [34:0] _GEN_568;
  wire [34:0] _GEN_570;
  wire [34:0] _GEN_571;
  wire [34:0] _GEN_572;
  wire [34:0] _GEN_574;
  wire [34:0] _GEN_575;
  wire [34:0] _GEN_576;
  wire [34:0] _GEN_578;
  wire [34:0] _GEN_579;
  wire [34:0] _GEN_580;
  wire [34:0] _GEN_582;
  wire [34:0] _GEN_583;
  wire [34:0] _GEN_584;
  wire [1:0] ppn_hi; // @[TLB.scala 105:26]
  wire [26:0] _ppn_T_1; // @[TLB.scala 108:28]
  wire [26:0] _GEN_953; // @[TLB.scala 108:47]
  wire [26:0] _ppn_T_2; // @[TLB.scala 108:47]
  wire [8:0] ppn_lo; // @[TLB.scala 108:58]
  wire [26:0] _ppn_T_4; // @[TLB.scala 108:47]
  wire [8:0] ppn_lo_1; // @[TLB.scala 108:58]
  wire [19:0] _ppn_T_5; // @[Cat.scala 30:58]
  wire [1:0] ppn_hi_2; // @[TLB.scala 105:26]
  wire [26:0] _ppn_T_6; // @[TLB.scala 108:28]
  wire [26:0] _GEN_955; // @[TLB.scala 108:47]
  wire [26:0] _ppn_T_7; // @[TLB.scala 108:47]
  wire [8:0] ppn_lo_2; // @[TLB.scala 108:58]
  wire [26:0] _ppn_T_9; // @[TLB.scala 108:47]
  wire [8:0] ppn_lo_3; // @[TLB.scala 108:58]
  wire [19:0] _ppn_T_10; // @[Cat.scala 30:58]
  wire [1:0] ppn_hi_4; // @[TLB.scala 105:26]
  wire [26:0] _ppn_T_11; // @[TLB.scala 108:28]
  wire [26:0] _GEN_957; // @[TLB.scala 108:47]
  wire [26:0] _ppn_T_12; // @[TLB.scala 108:47]
  wire [8:0] ppn_lo_4; // @[TLB.scala 108:58]
  wire [26:0] _ppn_T_14; // @[TLB.scala 108:47]
  wire [8:0] ppn_lo_5; // @[TLB.scala 108:58]
  wire [19:0] _ppn_T_15; // @[Cat.scala 30:58]
  wire [1:0] ppn_hi_6; // @[TLB.scala 105:26]
  wire [26:0] _ppn_T_16; // @[TLB.scala 108:28]
  wire [26:0] _GEN_959; // @[TLB.scala 108:47]
  wire [26:0] _ppn_T_17; // @[TLB.scala 108:47]
  wire [8:0] ppn_lo_6; // @[TLB.scala 108:58]
  wire [26:0] _ppn_T_19; // @[TLB.scala 108:47]
  wire [8:0] ppn_lo_7; // @[TLB.scala 108:58]
  wire [19:0] _ppn_T_20; // @[Cat.scala 30:58]
  wire [1:0] ppn_hi_8; // @[TLB.scala 105:26]
  wire [26:0] _GEN_961; // @[TLB.scala 108:47]
  wire [26:0] _ppn_T_22; // @[TLB.scala 108:47]
  wire [8:0] ppn_lo_8; // @[TLB.scala 108:58]
  wire [26:0] _ppn_T_24; // @[TLB.scala 108:47]
  wire [8:0] ppn_lo_9; // @[TLB.scala 108:58]
  wire [19:0] _ppn_T_25; // @[Cat.scala 30:58]
  wire [19:0] _ppn_T_27; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_28; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_29; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_30; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_31; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_32; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_33; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_34; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_35; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_36; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_37; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_38; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_39; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_40; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_41; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_42; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_43; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_44; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_45; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_46; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_47; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_48; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_49; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_50; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_51; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_52; // @[Mux.scala 27:72]
  wire [19:0] ppn; // @[Mux.scala 27:72]
  wire [5:0] ptw_ae_array_lo; // @[Cat.scala 30:58]
  wire [13:0] ptw_ae_array; // @[Cat.scala 30:58]
  wire  _priv_rw_ok_T_1; // @[TLB.scala 265:32]
  wire [5:0] priv_rw_ok_lo; // @[Cat.scala 30:58]
  wire [12:0] _priv_rw_ok_T_2; // @[Cat.scala 30:58]
  wire [12:0] _priv_rw_ok_T_3; // @[TLB.scala 265:23]
  wire [12:0] _priv_rw_ok_T_6; // @[TLB.scala 265:89]
  wire [12:0] priv_rw_ok; // @[TLB.scala 265:84]
  wire [5:0] r_array_lo; // @[Cat.scala 30:58]
  wire [12:0] _r_array_T; // @[Cat.scala 30:58]
  wire [5:0] r_array_lo_1; // @[Cat.scala 30:58]
  wire [12:0] _r_array_T_1; // @[Cat.scala 30:58]
  wire [12:0] _r_array_T_2; // @[TLB.scala 267:73]
  wire [12:0] _r_array_T_3; // @[TLB.scala 267:68]
  wire [12:0] r_array_lo_2; // @[TLB.scala 267:40]
  wire [13:0] r_array; // @[Cat.scala 30:58]
  wire [5:0] w_array_lo; // @[Cat.scala 30:58]
  wire [12:0] _w_array_T; // @[Cat.scala 30:58]
  wire [12:0] w_array_lo_1; // @[TLB.scala 268:40]
  wire [13:0] w_array; // @[Cat.scala 30:58]
  wire [1:0] pr_array_hi; // @[Bitwise.scala 72:12]
  wire [5:0] pr_array_lo; // @[Cat.scala 30:58]
  wire [13:0] _pr_array_T_1; // @[Cat.scala 30:58]
  wire [13:0] pr_array; // @[TLB.scala 270:87]
  wire [1:0] pw_array_hi; // @[Bitwise.scala 72:12]
  wire [5:0] pw_array_lo; // @[Cat.scala 30:58]
  wire [13:0] _pw_array_T_1; // @[Cat.scala 30:58]
  wire [13:0] pw_array; // @[TLB.scala 271:87]
  wire [1:0] eff_array_hi; // @[Bitwise.scala 72:12]
  wire [5:0] eff_array_lo; // @[Cat.scala 30:58]
  wire [13:0] eff_array; // @[Cat.scala 30:58]
  wire [1:0] c_array_hi; // @[Bitwise.scala 72:12]
  wire [5:0] c_array_lo; // @[Cat.scala 30:58]
  wire [13:0] c_array; // @[Cat.scala 30:58]
  wire [1:0] ppp_array_hi; // @[Bitwise.scala 72:12]
  wire [5:0] ppp_array_lo; // @[Cat.scala 30:58]
  wire [13:0] ppp_array; // @[Cat.scala 30:58]
  wire [1:0] paa_array_hi; // @[Bitwise.scala 72:12]
  wire [5:0] paa_array_lo; // @[Cat.scala 30:58]
  wire [13:0] paa_array; // @[Cat.scala 30:58]
  wire [5:0] pal_array_lo; // @[Cat.scala 30:58]
  wire [13:0] pal_array; // @[Cat.scala 30:58]
  wire [13:0] ppp_array_if_cached; // @[TLB.scala 278:39]
  wire [13:0] paa_array_if_cached; // @[TLB.scala 279:39]
  wire [13:0] pal_array_if_cached; // @[TLB.scala 280:39]
  wire [3:0] _misaligned_T; // @[OneHot.scala 58:35]
  wire [3:0] _misaligned_T_2; // @[TLB.scala 283:69]
  wire [39:0] _GEN_963; // @[TLB.scala 283:39]
  wire [39:0] _misaligned_T_3; // @[TLB.scala 283:39]
  wire  misaligned; // @[TLB.scala 283:75]
  wire [39:0] bad_va_maskedVAddr; // @[TLB.scala 289:43]
  wire  _bad_va_T_1; // @[TLB.scala 290:61]
  wire  _bad_va_T_2; // @[TLB.scala 290:82]
  wire  _bad_va_T_3; // @[TLB.scala 290:67]
  wire  bad_va; // @[TLB.scala 284:117]
  wire  _cmd_lrsc_T; // @[package.scala 15:47]
  wire  _cmd_lrsc_T_1; // @[package.scala 15:47]
  wire  cmd_lrsc; // @[package.scala 72:59]
  wire  _cmd_amo_logical_T; // @[package.scala 15:47]
  wire  _cmd_amo_logical_T_1; // @[package.scala 15:47]
  wire  _cmd_amo_logical_T_2; // @[package.scala 15:47]
  wire  _cmd_amo_logical_T_3; // @[package.scala 15:47]
  wire  _cmd_amo_logical_T_4; // @[package.scala 72:59]
  wire  _cmd_amo_logical_T_5; // @[package.scala 72:59]
  wire  cmd_amo_logical; // @[package.scala 72:59]
  wire  _cmd_amo_arithmetic_T; // @[package.scala 15:47]
  wire  _cmd_amo_arithmetic_T_1; // @[package.scala 15:47]
  wire  _cmd_amo_arithmetic_T_2; // @[package.scala 15:47]
  wire  _cmd_amo_arithmetic_T_3; // @[package.scala 15:47]
  wire  _cmd_amo_arithmetic_T_4; // @[package.scala 15:47]
  wire  _cmd_amo_arithmetic_T_5; // @[package.scala 72:59]
  wire  _cmd_amo_arithmetic_T_6; // @[package.scala 72:59]
  wire  _cmd_amo_arithmetic_T_7; // @[package.scala 72:59]
  wire  cmd_amo_arithmetic; // @[package.scala 72:59]
  wire  cmd_put_partial; // @[TLB.scala 297:41]
  wire  _cmd_read_T; // @[Consts.scala 81:31]
  wire  _cmd_read_T_2; // @[Consts.scala 81:41]
  wire  _cmd_read_T_4; // @[Consts.scala 81:58]
  wire  _cmd_read_T_21; // @[Consts.scala 79:44]
  wire  cmd_read; // @[Consts.scala 81:75]
  wire  _cmd_write_T; // @[Consts.scala 82:32]
  wire  _cmd_write_T_2; // @[Consts.scala 82:42]
  wire  _cmd_write_T_4; // @[Consts.scala 82:59]
  wire  cmd_write; // @[Consts.scala 82:76]
  wire  _cmd_write_perms_T; // @[package.scala 15:47]
  wire  _cmd_write_perms_T_1; // @[package.scala 15:47]
  wire  _cmd_write_perms_T_2; // @[package.scala 72:59]
  wire  cmd_write_perms; // @[TLB.scala 300:35]
  wire [13:0] _ae_array_T; // @[TLB.scala 305:8]
  wire [13:0] _ae_array_T_2; // @[TLB.scala 306:8]
  wire [13:0] ae_array; // @[TLB.scala 305:37]
  wire [13:0] _ae_ld_array_T_1; // @[TLB.scala 307:44]
  wire [13:0] ae_ld_array; // @[TLB.scala 307:24]
  wire [13:0] _ae_st_array_T_1; // @[TLB.scala 309:35]
  wire [13:0] _ae_st_array_T_2; // @[TLB.scala 309:8]
  wire [13:0] _ae_st_array_T_4; // @[TLB.scala 310:8]
  wire [13:0] _ae_st_array_T_5; // @[TLB.scala 309:53]
  wire [13:0] _ae_st_array_T_7; // @[TLB.scala 311:8]
  wire [13:0] _ae_st_array_T_8; // @[TLB.scala 310:53]
  wire [13:0] _ae_st_array_T_10; // @[TLB.scala 312:8]
  wire [13:0] ae_st_array; // @[TLB.scala 311:53]
  wire  _ma_ld_array_T; // @[TLB.scala 318:36]
  wire [13:0] ma_ld_array; // @[TLB.scala 318:24]
  wire  _ma_st_array_T; // @[TLB.scala 319:36]
  wire [13:0] ma_st_array; // @[TLB.scala 319:24]
  wire [13:0] _pf_ld_array_T; // @[TLB.scala 320:45]
  wire [13:0] pf_ld_array; // @[TLB.scala 320:24]
  wire [13:0] _pf_st_array_T; // @[TLB.scala 321:52]
  wire [13:0] pf_st_array; // @[TLB.scala 321:24]
  wire  tlb_hit; // @[TLB.scala 324:27]
  wire  _tlb_miss_T_1; // @[TLB.scala 325:29]
  wire  tlb_miss; // @[TLB.scala 325:40]
  reg [6:0] state_vec_0; // @[Replacement.scala 305:17]
  reg [31:0] _RAND_98;
  reg [2:0] state_reg_1; // @[Replacement.scala 168:70]
  reg [31:0] _RAND_99;
  wire  _T_23; // @[TLB.scala 329:22]
  wire  _T_24; // @[package.scala 72:59]
  wire  _T_25; // @[package.scala 72:59]
  wire  _T_26; // @[package.scala 72:59]
  wire  _T_27; // @[package.scala 72:59]
  wire  _T_28; // @[package.scala 72:59]
  wire  _T_29; // @[package.scala 72:59]
  wire  _T_30; // @[package.scala 72:59]
  wire [7:0] _T_31; // @[Cat.scala 30:58]
  wire [3:0] hi_1; // @[OneHot.scala 30:18]
  wire [3:0] lo_1; // @[OneHot.scala 31:18]
  wire  hi_2; // @[OneHot.scala 32:14]
  wire [3:0] _T_32; // @[OneHot.scala 32:28]
  wire [1:0] hi_3; // @[OneHot.scala 30:18]
  wire [1:0] lo_2; // @[OneHot.scala 31:18]
  wire  hi_4; // @[OneHot.scala 32:14]
  wire [1:0] _T_33; // @[OneHot.scala 32:28]
  wire  lo_3; // @[CircuitMath.scala 30:8]
  wire [2:0] state_vec_0_touch_way_sized; // @[Cat.scala 30:58]
  wire  state_vec_0_hi_hi; // @[Replacement.scala 196:33]
  wire [2:0] state_vec_0_left_subtree_state; // @[package.scala 154:13]
  wire [2:0] state_vec_0_right_subtree_state; // @[Replacement.scala 198:38]
  wire  state_vec_0_hi_hi_1; // @[Replacement.scala 196:33]
  wire  state_vec_0_left_subtree_state_1; // @[package.scala 154:13]
  wire  state_vec_0_right_subtree_state_1; // @[Replacement.scala 198:38]
  wire  state_vec_0_hi_lo; // @[Replacement.scala 203:16]
  wire  state_vec_0_lo; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_0_T_7; // @[Cat.scala 30:58]
  wire [2:0] state_vec_0_hi_lo_1; // @[Replacement.scala 203:16]
  wire  state_vec_0_left_subtree_state_2; // @[package.scala 154:13]
  wire  state_vec_0_right_subtree_state_2; // @[Replacement.scala 198:38]
  wire  state_vec_0_hi_lo_2; // @[Replacement.scala 203:16]
  wire  state_vec_0_lo_1; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_0_T_15; // @[Cat.scala 30:58]
  wire [2:0] state_vec_0_lo_2; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_0_T_16; // @[Cat.scala 30:58]
  wire  _T_35; // @[package.scala 72:59]
  wire  _T_36; // @[package.scala 72:59]
  wire  _T_37; // @[package.scala 72:59]
  wire [3:0] _T_38; // @[Cat.scala 30:58]
  wire [1:0] hi_6; // @[OneHot.scala 30:18]
  wire [1:0] lo_6; // @[OneHot.scala 31:18]
  wire  hi_7; // @[OneHot.scala 32:14]
  wire [1:0] _T_39; // @[OneHot.scala 32:28]
  wire  lo_7; // @[CircuitMath.scala 30:8]
  wire [1:0] state_reg_touch_way_sized; // @[Cat.scala 30:58]
  wire  state_reg_hi_hi; // @[Replacement.scala 196:33]
  wire  state_reg_left_subtree_state; // @[package.scala 154:13]
  wire  state_reg_right_subtree_state; // @[Replacement.scala 198:38]
  wire  state_reg_hi_lo; // @[Replacement.scala 203:16]
  wire  state_reg_lo; // @[Replacement.scala 206:16]
  wire [2:0] _state_reg_T_6; // @[Cat.scala 30:58]
  wire  multipleHits_leftOne; // @[Misc.scala 180:37]
  wire  multipleHits_leftOne_1; // @[Misc.scala 180:37]
  wire  multipleHits_rightOne; // @[Misc.scala 181:39]
  wire  multipleHits_rightOne_1; // @[Misc.scala 182:16]
  wire  multipleHits_rightTwo; // @[Misc.scala 182:61]
  wire  multipleHits_leftOne_2; // @[Misc.scala 182:16]
  wire  _multipleHits_T_9; // @[Misc.scala 182:61]
  wire  multipleHits_leftTwo; // @[Misc.scala 182:49]
  wire  multipleHits_leftOne_3; // @[Misc.scala 180:37]
  wire  multipleHits_leftOne_4; // @[Misc.scala 180:37]
  wire  multipleHits_rightOne_2; // @[Misc.scala 181:39]
  wire  multipleHits_rightOne_3; // @[Misc.scala 182:16]
  wire  multipleHits_rightTwo_1; // @[Misc.scala 182:61]
  wire  multipleHits_rightOne_4; // @[Misc.scala 182:16]
  wire  _multipleHits_T_18; // @[Misc.scala 182:61]
  wire  multipleHits_rightTwo_2; // @[Misc.scala 182:49]
  wire  multipleHits_leftOne_5; // @[Misc.scala 182:16]
  wire  _multipleHits_T_19; // @[Misc.scala 182:37]
  wire  _multipleHits_T_20; // @[Misc.scala 182:61]
  wire  multipleHits_leftTwo_1; // @[Misc.scala 182:49]
  wire  multipleHits_leftOne_6; // @[Misc.scala 180:37]
  wire  multipleHits_leftOne_7; // @[Misc.scala 180:37]
  wire  multipleHits_rightOne_5; // @[Misc.scala 181:39]
  wire  multipleHits_rightOne_6; // @[Misc.scala 182:16]
  wire  multipleHits_rightTwo_3; // @[Misc.scala 182:61]
  wire  multipleHits_leftOne_8; // @[Misc.scala 182:16]
  wire  _multipleHits_T_30; // @[Misc.scala 182:61]
  wire  multipleHits_leftTwo_2; // @[Misc.scala 182:49]
  wire  multipleHits_leftOne_9; // @[Misc.scala 180:37]
  wire  multipleHits_rightOne_7; // @[Misc.scala 181:39]
  wire  multipleHits_leftOne_10; // @[Misc.scala 182:16]
  wire  multipleHits_leftTwo_3; // @[Misc.scala 182:61]
  wire  multipleHits_leftOne_11; // @[Misc.scala 180:37]
  wire  multipleHits_rightOne_8; // @[Misc.scala 181:39]
  wire  multipleHits_rightOne_9; // @[Misc.scala 182:16]
  wire  multipleHits_rightTwo_4; // @[Misc.scala 182:61]
  wire  multipleHits_rightOne_10; // @[Misc.scala 182:16]
  wire  _multipleHits_T_42; // @[Misc.scala 182:37]
  wire  _multipleHits_T_43; // @[Misc.scala 182:61]
  wire  multipleHits_rightTwo_5; // @[Misc.scala 182:49]
  wire  multipleHits_rightOne_11; // @[Misc.scala 182:16]
  wire  _multipleHits_T_44; // @[Misc.scala 182:37]
  wire  _multipleHits_T_45; // @[Misc.scala 182:61]
  wire  multipleHits_rightTwo_6; // @[Misc.scala 182:49]
  wire  _multipleHits_T_47; // @[Misc.scala 182:37]
  wire  _multipleHits_T_48; // @[Misc.scala 182:61]
  wire  multipleHits; // @[Misc.scala 182:49]
  wire  _io_resp_pf_ld_T; // @[TLB.scala 342:28]
  wire [13:0] _io_resp_pf_ld_T_1; // @[TLB.scala 342:57]
  wire  _io_resp_pf_ld_T_2; // @[TLB.scala 342:65]
  wire  _io_resp_pf_st_T; // @[TLB.scala 343:28]
  wire [13:0] _io_resp_pf_st_T_1; // @[TLB.scala 343:64]
  wire  _io_resp_pf_st_T_2; // @[TLB.scala 343:72]
  wire [13:0] _io_resp_ae_ld_T; // @[TLB.scala 345:33]
  wire [13:0] _io_resp_ae_st_T; // @[TLB.scala 346:33]
  wire [13:0] _io_resp_ma_ld_T; // @[TLB.scala 348:33]
  wire [13:0] _io_resp_ma_st_T; // @[TLB.scala 349:33]
  wire [13:0] _io_resp_cacheable_T; // @[TLB.scala 351:33]
  wire  _io_resp_miss_T; // @[TLB.scala 354:29]
  wire  _T_41; // @[Decoupled.scala 40:37]
  wire  _T_42; // @[TLB.scala 363:25]
  wire  r_superpage_repl_addr_hi; // @[Replacement.scala 243:38]
  wire  r_superpage_repl_addr_lo; // @[Replacement.scala 250:16]
  wire [1:0] _r_superpage_repl_addr_T_2; // @[Cat.scala 30:58]
  wire [3:0] r_superpage_repl_addr_valids; // @[Cat.scala 30:58]
  wire  _r_superpage_repl_addr_T_3; // @[TLB.scala 411:16]
  wire  _r_superpage_repl_addr_T_5; // @[OneHot.scala 47:40]
  wire  _r_superpage_repl_addr_T_6; // @[OneHot.scala 47:40]
  wire  _r_superpage_repl_addr_T_7; // @[OneHot.scala 47:40]
  wire  r_sectored_repl_addr_hi; // @[Replacement.scala 243:38]
  wire  r_sectored_repl_addr_hi_1; // @[Replacement.scala 243:38]
  wire  r_sectored_repl_addr_lo; // @[Replacement.scala 250:16]
  wire [1:0] _r_sectored_repl_addr_T_2; // @[Cat.scala 30:58]
  wire  r_sectored_repl_addr_hi_2; // @[Replacement.scala 243:38]
  wire  r_sectored_repl_addr_lo_1; // @[Replacement.scala 250:16]
  wire [1:0] _r_sectored_repl_addr_T_5; // @[Cat.scala 30:58]
  wire [1:0] r_sectored_repl_addr_lo_2; // @[Replacement.scala 250:16]
  wire [2:0] _r_sectored_repl_addr_T_6; // @[Cat.scala 30:58]
  wire [7:0] r_sectored_repl_addr_valids; // @[Cat.scala 30:58]
  wire  _r_sectored_repl_addr_T_7; // @[TLB.scala 411:16]
  wire  _r_sectored_repl_addr_T_9; // @[OneHot.scala 47:40]
  wire  _r_sectored_repl_addr_T_10; // @[OneHot.scala 47:40]
  wire  _r_sectored_repl_addr_T_11; // @[OneHot.scala 47:40]
  wire  _r_sectored_repl_addr_T_12; // @[OneHot.scala 47:40]
  wire  _r_sectored_repl_addr_T_13; // @[OneHot.scala 47:40]
  wire  _r_sectored_repl_addr_T_14; // @[OneHot.scala 47:40]
  wire  _r_sectored_repl_addr_T_15; // @[OneHot.scala 47:40]
  wire  _T_44; // @[TLB.scala 377:17]
  wire  _T_45; // @[TLB.scala 377:28]
  wire  _T_48; // @[TLB.scala 385:72]
  wire  _T_49; // @[TLB.scala 385:34]
  wire  _T_51; // @[TLB.scala 385:13]
  wire  _T_59; // @[TLB.scala 134:61]
  wire  _GEN_617; // @[TLB.scala 142:19]
  wire  _GEN_618; // @[TLB.scala 142:19]
  wire  _GEN_619; // @[TLB.scala 142:19]
  wire  _GEN_620; // @[TLB.scala 142:19]
  wire  _GEN_621; // @[TLB.scala 388:40]
  wire  _GEN_622; // @[TLB.scala 388:40]
  wire  _GEN_623; // @[TLB.scala 388:40]
  wire  _GEN_624; // @[TLB.scala 388:40]
  wire  _T_198; // @[TLB.scala 134:61]
  wire  _GEN_645; // @[TLB.scala 142:19]
  wire  _GEN_646; // @[TLB.scala 142:19]
  wire  _GEN_647; // @[TLB.scala 142:19]
  wire  _GEN_648; // @[TLB.scala 142:19]
  wire  _GEN_649; // @[TLB.scala 388:40]
  wire  _GEN_650; // @[TLB.scala 388:40]
  wire  _GEN_651; // @[TLB.scala 388:40]
  wire  _GEN_652; // @[TLB.scala 388:40]
  wire  _T_337; // @[TLB.scala 134:61]
  wire  _GEN_673; // @[TLB.scala 142:19]
  wire  _GEN_674; // @[TLB.scala 142:19]
  wire  _GEN_675; // @[TLB.scala 142:19]
  wire  _GEN_676; // @[TLB.scala 142:19]
  wire  _GEN_677; // @[TLB.scala 388:40]
  wire  _GEN_678; // @[TLB.scala 388:40]
  wire  _GEN_679; // @[TLB.scala 388:40]
  wire  _GEN_680; // @[TLB.scala 388:40]
  wire  _T_476; // @[TLB.scala 134:61]
  wire  _GEN_701; // @[TLB.scala 142:19]
  wire  _GEN_702; // @[TLB.scala 142:19]
  wire  _GEN_703; // @[TLB.scala 142:19]
  wire  _GEN_704; // @[TLB.scala 142:19]
  wire  _GEN_705; // @[TLB.scala 388:40]
  wire  _GEN_706; // @[TLB.scala 388:40]
  wire  _GEN_707; // @[TLB.scala 388:40]
  wire  _GEN_708; // @[TLB.scala 388:40]
  wire  _T_615; // @[TLB.scala 134:61]
  wire  _GEN_729; // @[TLB.scala 142:19]
  wire  _GEN_730; // @[TLB.scala 142:19]
  wire  _GEN_731; // @[TLB.scala 142:19]
  wire  _GEN_732; // @[TLB.scala 142:19]
  wire  _GEN_733; // @[TLB.scala 388:40]
  wire  _GEN_734; // @[TLB.scala 388:40]
  wire  _GEN_735; // @[TLB.scala 388:40]
  wire  _GEN_736; // @[TLB.scala 388:40]
  wire  _T_754; // @[TLB.scala 134:61]
  wire  _GEN_757; // @[TLB.scala 142:19]
  wire  _GEN_758; // @[TLB.scala 142:19]
  wire  _GEN_759; // @[TLB.scala 142:19]
  wire  _GEN_760; // @[TLB.scala 142:19]
  wire  _GEN_761; // @[TLB.scala 388:40]
  wire  _GEN_762; // @[TLB.scala 388:40]
  wire  _GEN_763; // @[TLB.scala 388:40]
  wire  _GEN_764; // @[TLB.scala 388:40]
  wire  _T_893; // @[TLB.scala 134:61]
  wire  _GEN_785; // @[TLB.scala 142:19]
  wire  _GEN_786; // @[TLB.scala 142:19]
  wire  _GEN_787; // @[TLB.scala 142:19]
  wire  _GEN_788; // @[TLB.scala 142:19]
  wire  _GEN_789; // @[TLB.scala 388:40]
  wire  _GEN_790; // @[TLB.scala 388:40]
  wire  _GEN_791; // @[TLB.scala 388:40]
  wire  _GEN_792; // @[TLB.scala 388:40]
  wire  _T_1032; // @[TLB.scala 134:61]
  wire  _GEN_813; // @[TLB.scala 142:19]
  wire  _GEN_814; // @[TLB.scala 142:19]
  wire  _GEN_815; // @[TLB.scala 142:19]
  wire  _GEN_816; // @[TLB.scala 142:19]
  wire  _GEN_817; // @[TLB.scala 388:40]
  wire  _GEN_818; // @[TLB.scala 388:40]
  wire  _GEN_819; // @[TLB.scala 388:40]
  wire  _GEN_820; // @[TLB.scala 388:40]
  wire  _GEN_826; // @[TLB.scala 142:19]
  wire  _GEN_827; // @[TLB.scala 388:40]
  wire  _GEN_830; // @[TLB.scala 142:19]
  wire  _GEN_831; // @[TLB.scala 388:40]
  wire  _GEN_834; // @[TLB.scala 142:19]
  wire  _GEN_835; // @[TLB.scala 388:40]
  wire  _GEN_838; // @[TLB.scala 142:19]
  wire  _GEN_839; // @[TLB.scala 388:40]
  wire  _GEN_842; // @[TLB.scala 142:19]
  wire  _GEN_843; // @[TLB.scala 388:40]
  wire  _T_1326; // @[TLB.scala 392:24]
  reg [19:0] TLB_state; // @[Register tracking TLB state]
  reg [31:0] _RAND_100;
  reg  TLB_cov [0:1048575]; // @[Coverage map for TLB]
  reg [31:0] _RAND_101;
  wire  TLB_cov_read_data; // @[Coverage map for TLB]
  wire [19:0] TLB_cov_read_addr; // @[Coverage map for TLB]
  wire  TLB_cov_write_data; // @[Coverage map for TLB]
  wire [19:0] TLB_cov_write_addr; // @[Coverage map for TLB]
  wire  TLB_cov_write_mask; // @[Coverage map for TLB]
  wire  TLB_cov_write_en; // @[Coverage map for TLB]
  reg [29:0] TLB_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_102;
  wire  mux_cond_0;
  wire  mux_cond_1;
  wire  mux_cond_2;
  wire  mux_cond_3;
  wire  mux_cond_4;
  wire  mux_cond_5;
  wire  mux_cond_6;
  wire  mux_cond_7;
  wire  mux_cond_8;
  wire  mux_cond_9;
  wire  mux_cond_10;
  wire  mux_cond_11;
  wire  mux_cond_12;
  wire  mux_cond_13;
  wire  mux_cond_14;
  wire  mux_cond_15;
  wire  mux_cond_16;
  wire  mux_cond_17;
  wire  mux_cond_18;
  wire  mux_cond_19;
  wire  mux_cond_20;
  wire  mux_cond_21;
  wire  mux_cond_22;
  wire  mux_cond_23;
  wire  mux_cond_24;
  wire  mux_cond_25;
  wire  mux_cond_26;
  wire  mux_cond_27;
  wire  mux_cond_28;
  wire  mux_cond_29;
  wire  mux_cond_30;
  wire  mux_cond_31;
  wire  mux_cond_32;
  wire  mux_cond_33;
  wire  mux_cond_34;
  wire  mux_cond_35;
  wire  mux_cond_36;
  wire  mux_cond_37;
  wire  mux_cond_38;
  wire  mux_cond_39;
  wire  mux_cond_40;
  wire  mux_cond_41;
  wire  mux_cond_42;
  wire  mux_cond_43;
  wire  mux_cond_44;
  wire  mux_cond_45;
  wire  mux_cond_46;
  wire  mux_cond_47;
  wire  mux_cond_48;
  wire  mux_cond_49;
  wire  mux_cond_50;
  wire  mux_cond_51;
  wire  mux_cond_52;
  wire  mux_cond_53;
  wire  mux_cond_54;
  wire  mux_cond_55;
  wire  mux_cond_56;
  wire  mux_cond_57;
  wire  mux_cond_58;
  wire  mux_cond_59;
  wire  mux_cond_60;
  wire  mux_cond_61;
  wire  mux_cond_62;
  wire  mux_cond_63;
  wire  mux_cond_64;
  wire  mux_cond_65;
  wire  mux_cond_66;
  wire  mux_cond_67;
  wire  mux_cond_68;
  wire  r_sectored_hit_shl;
  wire [19:0] r_sectored_hit_pad;
  wire [9:0] r_sectored_repl_addr_shl;
  wire [19:0] r_sectored_repl_addr_pad;
  wire [19:0] r_superpage_repl_addr_shl;
  wire [19:0] r_superpage_repl_addr_pad;
  wire [7:0] special_entry_valid_0_shl;
  wire [19:0] special_entry_valid_0_pad;
  wire [19:0] special_entry_level_shl;
  wire [19:0] special_entry_level_pad;
  wire [7:0] state_shl;
  wire [19:0] state_pad;
  wire [14:0] r_sectored_hit_addr_shl;
  wire [19:0] r_sectored_hit_addr_pad;
  wire [5:0] mux_cond_0_shl;
  wire [19:0] mux_cond_0_pad;
  wire [11:0] mux_cond_1_shl;
  wire [19:0] mux_cond_1_pad;
  wire [2:0] mux_cond_2_shl;
  wire [19:0] mux_cond_2_pad;
  wire [12:0] mux_cond_3_shl;
  wire [19:0] mux_cond_3_pad;
  wire [11:0] mux_cond_4_shl;
  wire [19:0] mux_cond_4_pad;
  wire [1:0] mux_cond_5_shl;
  wire [19:0] mux_cond_5_pad;
  wire [13:0] mux_cond_6_shl;
  wire [19:0] mux_cond_6_pad;
  wire [6:0] mux_cond_7_shl;
  wire [19:0] mux_cond_7_pad;
  wire [4:0] mux_cond_8_shl;
  wire [19:0] mux_cond_8_pad;
  wire [17:0] mux_cond_9_shl;
  wire [19:0] mux_cond_9_pad;
  wire [5:0] mux_cond_10_shl;
  wire [19:0] mux_cond_10_pad;
  wire [9:0] mux_cond_11_shl;
  wire [19:0] mux_cond_11_pad;
  wire [1:0] mux_cond_12_shl;
  wire [19:0] mux_cond_12_pad;
  wire [9:0] mux_cond_13_shl;
  wire [19:0] mux_cond_13_pad;
  wire [12:0] mux_cond_14_shl;
  wire [19:0] mux_cond_14_pad;
  wire [7:0] mux_cond_15_shl;
  wire [19:0] mux_cond_15_pad;
  wire [6:0] mux_cond_16_shl;
  wire [19:0] mux_cond_16_pad;
  wire [7:0] mux_cond_17_shl;
  wire [19:0] mux_cond_17_pad;
  wire [16:0] mux_cond_18_shl;
  wire [19:0] mux_cond_18_pad;
  wire [8:0] mux_cond_19_shl;
  wire [19:0] mux_cond_19_pad;
  wire [1:0] mux_cond_20_shl;
  wire [19:0] mux_cond_20_pad;
  wire [5:0] mux_cond_21_shl;
  wire [19:0] mux_cond_21_pad;
  wire [11:0] mux_cond_22_shl;
  wire [19:0] mux_cond_22_pad;
  wire [2:0] mux_cond_23_shl;
  wire [19:0] mux_cond_23_pad;
  wire [14:0] mux_cond_24_shl;
  wire [19:0] mux_cond_24_pad;
  wire [3:0] mux_cond_25_shl;
  wire [19:0] mux_cond_25_pad;
  wire [11:0] mux_cond_26_shl;
  wire [19:0] mux_cond_26_pad;
  wire  mux_cond_27_shl;
  wire [19:0] mux_cond_27_pad;
  wire [18:0] mux_cond_28_shl;
  wire [19:0] mux_cond_28_pad;
  wire [14:0] mux_cond_29_shl;
  wire [19:0] mux_cond_29_pad;
  wire [8:0] mux_cond_30_shl;
  wire [19:0] mux_cond_30_pad;
  wire [3:0] mux_cond_31_shl;
  wire [19:0] mux_cond_31_pad;
  wire [2:0] mux_cond_32_shl;
  wire [19:0] mux_cond_32_pad;
  wire  mux_cond_33_shl;
  wire [19:0] mux_cond_33_pad;
  wire [7:0] mux_cond_34_shl;
  wire [19:0] mux_cond_34_pad;
  wire [4:0] mux_cond_35_shl;
  wire [19:0] mux_cond_35_pad;
  wire [3:0] mux_cond_36_shl;
  wire [19:0] mux_cond_36_pad;
  wire [4:0] mux_cond_37_shl;
  wire [19:0] mux_cond_37_pad;
  wire [12:0] mux_cond_38_shl;
  wire [19:0] mux_cond_38_pad;
  wire [9:0] mux_cond_39_shl;
  wire [19:0] mux_cond_39_pad;
  wire  mux_cond_40_shl;
  wire [19:0] mux_cond_40_pad;
  wire [16:0] mux_cond_41_shl;
  wire [19:0] mux_cond_41_pad;
  wire [4:0] mux_cond_42_shl;
  wire [19:0] mux_cond_42_pad;
  wire [18:0] mux_cond_43_shl;
  wire [19:0] mux_cond_43_pad;
  wire [8:0] mux_cond_44_shl;
  wire [19:0] mux_cond_44_pad;
  wire [17:0] mux_cond_45_shl;
  wire [19:0] mux_cond_45_pad;
  wire [5:0] mux_cond_46_shl;
  wire [19:0] mux_cond_46_pad;
  wire [8:0] mux_cond_47_shl;
  wire [19:0] mux_cond_47_pad;
  wire [7:0] mux_cond_48_shl;
  wire [19:0] mux_cond_48_pad;
  wire [16:0] mux_cond_49_shl;
  wire [19:0] mux_cond_49_pad;
  wire [8:0] mux_cond_50_shl;
  wire [19:0] mux_cond_50_pad;
  wire [4:0] mux_cond_51_shl;
  wire [19:0] mux_cond_51_pad;
  wire [3:0] mux_cond_52_shl;
  wire [19:0] mux_cond_52_pad;
  wire [6:0] mux_cond_53_shl;
  wire [19:0] mux_cond_53_pad;
  wire [18:0] mux_cond_54_shl;
  wire [19:0] mux_cond_54_pad;
  wire [15:0] mux_cond_55_shl;
  wire [19:0] mux_cond_55_pad;
  wire [16:0] mux_cond_56_shl;
  wire [19:0] mux_cond_56_pad;
  wire [7:0] mux_cond_57_shl;
  wire [19:0] mux_cond_57_pad;
  wire [11:0] mux_cond_58_shl;
  wire [19:0] mux_cond_58_pad;
  wire [14:0] mux_cond_59_shl;
  wire [19:0] mux_cond_59_pad;
  wire [13:0] mux_cond_60_shl;
  wire [19:0] mux_cond_60_pad;
  wire [8:0] mux_cond_61_shl;
  wire [19:0] mux_cond_61_pad;
  wire [7:0] mux_cond_62_shl;
  wire [19:0] mux_cond_62_pad;
  wire [6:0] mux_cond_63_shl;
  wire [19:0] mux_cond_63_pad;
  wire [19:0] mux_cond_64_shl;
  wire [19:0] mux_cond_64_pad;
  wire [11:0] mux_cond_65_shl;
  wire [19:0] mux_cond_65_pad;
  wire [6:0] mux_cond_66_shl;
  wire [19:0] mux_cond_66_pad;
  wire [10:0] mux_cond_67_shl;
  wire [19:0] mux_cond_67_pad;
  wire [13:0] mux_cond_68_shl;
  wire [19:0] mux_cond_68_pad;
  wire [16:0] sectored_entries_0_0_valid_3_shl;
  wire [19:0] sectored_entries_0_0_valid_3_pad;
  wire [8:0] sectored_entries_0_0_valid_2_shl;
  wire [19:0] sectored_entries_0_0_valid_2_pad;
  wire [8:0] sectored_entries_0_2_valid_0_shl;
  wire [19:0] sectored_entries_0_2_valid_0_pad;
  wire [8:0] sectored_entries_0_3_valid_0_shl;
  wire [19:0] sectored_entries_0_3_valid_0_pad;
  wire [1:0] superpage_entries_2_level_shl;
  wire [19:0] superpage_entries_2_level_pad;
  wire  sectored_entries_0_7_valid_1_shl;
  wire [19:0] sectored_entries_0_7_valid_1_pad;
  wire [8:0] sectored_entries_0_4_valid_0_shl;
  wire [19:0] sectored_entries_0_4_valid_0_pad;
  wire [16:0] sectored_entries_0_1_valid_3_shl;
  wire [19:0] sectored_entries_0_1_valid_3_pad;
  wire  sectored_entries_0_1_valid_1_shl;
  wire [19:0] sectored_entries_0_1_valid_1_pad;
  wire [16:0] sectored_entries_0_2_valid_3_shl;
  wire [19:0] sectored_entries_0_2_valid_3_pad;
  wire  sectored_entries_0_2_valid_1_shl;
  wire [19:0] sectored_entries_0_2_valid_1_pad;
  wire [11:0] superpage_entries_1_valid_0_shl;
  wire [19:0] superpage_entries_1_valid_0_pad;
  wire [8:0] sectored_entries_0_7_valid_0_shl;
  wire [19:0] sectored_entries_0_7_valid_0_pad;
  wire [11:0] superpage_entries_3_valid_0_shl;
  wire [19:0] superpage_entries_3_valid_0_pad;
  wire [16:0] sectored_entries_0_5_valid_3_shl;
  wire [19:0] sectored_entries_0_5_valid_3_pad;
  wire  sectored_entries_0_5_valid_1_shl;
  wire [19:0] sectored_entries_0_5_valid_1_pad;
  wire [16:0] sectored_entries_0_4_valid_3_shl;
  wire [19:0] sectored_entries_0_4_valid_3_pad;
  wire [8:0] sectored_entries_0_5_valid_2_shl;
  wire [19:0] sectored_entries_0_5_valid_2_pad;
  wire [8:0] sectored_entries_0_1_valid_2_shl;
  wire [19:0] sectored_entries_0_1_valid_2_pad;
  wire  sectored_entries_0_3_valid_1_shl;
  wire [19:0] sectored_entries_0_3_valid_1_pad;
  wire [8:0] sectored_entries_0_1_valid_0_shl;
  wire [19:0] sectored_entries_0_1_valid_0_pad;
  wire [8:0] sectored_entries_0_4_valid_2_shl;
  wire [19:0] sectored_entries_0_4_valid_2_pad;
  wire  sectored_entries_0_4_valid_1_shl;
  wire [19:0] sectored_entries_0_4_valid_1_pad;
  wire [1:0] superpage_entries_3_level_shl;
  wire [19:0] superpage_entries_3_level_pad;
  wire  sectored_entries_0_0_valid_1_shl;
  wire [19:0] sectored_entries_0_0_valid_1_pad;
  wire [8:0] sectored_entries_0_3_valid_2_shl;
  wire [19:0] sectored_entries_0_3_valid_2_pad;
  wire  sectored_entries_0_6_valid_1_shl;
  wire [19:0] sectored_entries_0_6_valid_1_pad;
  wire [16:0] sectored_entries_0_7_valid_3_shl;
  wire [19:0] sectored_entries_0_7_valid_3_pad;
  wire [16:0] sectored_entries_0_3_valid_3_shl;
  wire [19:0] sectored_entries_0_3_valid_3_pad;
  wire [8:0] sectored_entries_0_0_valid_0_shl;
  wire [19:0] sectored_entries_0_0_valid_0_pad;
  wire [11:0] superpage_entries_0_valid_0_shl;
  wire [19:0] superpage_entries_0_valid_0_pad;
  wire [8:0] sectored_entries_0_2_valid_2_shl;
  wire [19:0] sectored_entries_0_2_valid_2_pad;
  wire [8:0] sectored_entries_0_6_valid_2_shl;
  wire [19:0] sectored_entries_0_6_valid_2_pad;
  wire [11:0] superpage_entries_2_valid_0_shl;
  wire [19:0] superpage_entries_2_valid_0_pad;
  wire [16:0] sectored_entries_0_6_valid_3_shl;
  wire [19:0] sectored_entries_0_6_valid_3_pad;
  wire [8:0] sectored_entries_0_6_valid_0_shl;
  wire [19:0] sectored_entries_0_6_valid_0_pad;
  wire [8:0] sectored_entries_0_7_valid_2_shl;
  wire [19:0] sectored_entries_0_7_valid_2_pad;
  wire [1:0] superpage_entries_0_level_shl;
  wire [19:0] superpage_entries_0_level_pad;
  wire [1:0] superpage_entries_1_level_shl;
  wire [19:0] superpage_entries_1_level_pad;
  wire [8:0] sectored_entries_0_5_valid_0_shl;
  wire [19:0] sectored_entries_0_5_valid_0_pad;
  wire [19:0] TLB_xor64;
  wire [19:0] TLB_xor31;
  wire [19:0] TLB_xor65;
  wire [19:0] TLB_xor66;
  wire [19:0] TLB_xor32;
  wire [19:0] TLB_xor15;
  wire [19:0] TLB_xor68;
  wire [19:0] TLB_xor33;
  wire [19:0] TLB_xor69;
  wire [19:0] TLB_xor70;
  wire [19:0] TLB_xor34;
  wire [19:0] TLB_xor16;
  wire [19:0] TLB_xor7;
  wire [19:0] TLB_xor72;
  wire [19:0] TLB_xor35;
  wire [19:0] TLB_xor73;
  wire [19:0] TLB_xor74;
  wire [19:0] TLB_xor36;
  wire [19:0] TLB_xor17;
  wire [19:0] TLB_xor75;
  wire [19:0] TLB_xor76;
  wire [19:0] TLB_xor37;
  wire [19:0] TLB_xor77;
  wire [19:0] TLB_xor78;
  wire [19:0] TLB_xor38;
  wire [19:0] TLB_xor18;
  wire [19:0] TLB_xor8;
  wire [19:0] TLB_xor3;
  wire [19:0] TLB_xor80;
  wire [19:0] TLB_xor39;
  wire [19:0] TLB_xor81;
  wire [19:0] TLB_xor82;
  wire [19:0] TLB_xor40;
  wire [19:0] TLB_xor19;
  wire [19:0] TLB_xor84;
  wire [19:0] TLB_xor41;
  wire [19:0] TLB_xor85;
  wire [19:0] TLB_xor86;
  wire [19:0] TLB_xor42;
  wire [19:0] TLB_xor20;
  wire [19:0] TLB_xor9;
  wire [19:0] TLB_xor88;
  wire [19:0] TLB_xor43;
  wire [19:0] TLB_xor89;
  wire [19:0] TLB_xor90;
  wire [19:0] TLB_xor44;
  wire [19:0] TLB_xor21;
  wire [19:0] TLB_xor91;
  wire [19:0] TLB_xor92;
  wire [19:0] TLB_xor45;
  wire [19:0] TLB_xor93;
  wire [19:0] TLB_xor94;
  wire [19:0] TLB_xor46;
  wire [19:0] TLB_xor22;
  wire [19:0] TLB_xor10;
  wire [19:0] TLB_xor4;
  wire [19:0] TLB_xor1;
  wire [19:0] TLB_xor96;
  wire [19:0] TLB_xor47;
  wire [19:0] TLB_xor97;
  wire [19:0] TLB_xor98;
  wire [19:0] TLB_xor48;
  wire [19:0] TLB_xor23;
  wire [19:0] TLB_xor100;
  wire [19:0] TLB_xor49;
  wire [19:0] TLB_xor101;
  wire [19:0] TLB_xor102;
  wire [19:0] TLB_xor50;
  wire [19:0] TLB_xor24;
  wire [19:0] TLB_xor11;
  wire [19:0] TLB_xor104;
  wire [19:0] TLB_xor51;
  wire [19:0] TLB_xor105;
  wire [19:0] TLB_xor106;
  wire [19:0] TLB_xor52;
  wire [19:0] TLB_xor25;
  wire [19:0] TLB_xor107;
  wire [19:0] TLB_xor108;
  wire [19:0] TLB_xor53;
  wire [19:0] TLB_xor109;
  wire [19:0] TLB_xor110;
  wire [19:0] TLB_xor54;
  wire [19:0] TLB_xor26;
  wire [19:0] TLB_xor12;
  wire [19:0] TLB_xor5;
  wire [19:0] TLB_xor112;
  wire [19:0] TLB_xor55;
  wire [19:0] TLB_xor113;
  wire [19:0] TLB_xor114;
  wire [19:0] TLB_xor56;
  wire [19:0] TLB_xor27;
  wire [19:0] TLB_xor116;
  wire [19:0] TLB_xor57;
  wire [19:0] TLB_xor117;
  wire [19:0] TLB_xor118;
  wire [19:0] TLB_xor58;
  wire [19:0] TLB_xor28;
  wire [19:0] TLB_xor13;
  wire [19:0] TLB_xor120;
  wire [19:0] TLB_xor59;
  wire [19:0] TLB_xor121;
  wire [19:0] TLB_xor122;
  wire [19:0] TLB_xor60;
  wire [19:0] TLB_xor29;
  wire [19:0] TLB_xor123;
  wire [19:0] TLB_xor124;
  wire [19:0] TLB_xor61;
  wire [19:0] TLB_xor125;
  wire [19:0] TLB_xor126;
  wire [19:0] TLB_xor62;
  wire [19:0] TLB_xor30;
  wire [19:0] TLB_xor14;
  wire [19:0] TLB_xor6;
  wire [19:0] TLB_xor2;
  wire [19:0] TLB_xor0;
  wire [29:0] mpu_ppn_barrier_sum;
  wire [29:0] entries_barrier_10_sum;
  wire [29:0] entries_barrier_9_sum;
  wire [29:0] entries_barrier_7_sum;
  wire [29:0] entries_barrier_sum;
  wire [29:0] entries_barrier_6_sum;
  wire [29:0] entries_barrier_12_sum;
  wire [29:0] entries_barrier_1_sum;
  wire [29:0] entries_barrier_11_sum;
  wire [29:0] entries_barrier_8_sum;
  wire [29:0] pmp_sum;
  wire [29:0] entries_barrier_2_sum;
  wire [29:0] entries_barrier_4_sum;
  wire [29:0] entries_barrier_5_sum;
  wire [29:0] entries_barrier_3_sum;
  wire  stopEn0;
  wire  entries_barrier_11_metaAssert_wire;
  wire  entries_barrier_8_metaAssert_wire;
  wire  entries_barrier_3_metaAssert_wire;
  wire  pmp_metaAssert_wire;
  wire  entries_barrier_6_metaAssert_wire;
  wire  entries_barrier_12_metaAssert_wire;
  wire  entries_barrier_9_metaAssert_wire;
  wire  mpu_ppn_barrier_metaAssert_wire;
  wire  entries_barrier_7_metaAssert_wire;
  wire  entries_barrier_metaAssert_wire;
  wire  entries_barrier_5_metaAssert_wire;
  wire  entries_barrier_2_metaAssert_wire;
  wire  entries_barrier_4_metaAssert_wire;
  wire  entries_barrier_1_metaAssert_wire;
  wire  entries_barrier_10_metaAssert_wire;
  wire  TLB_or7;
  wire  TLB_or8;
  wire  TLB_or3;
  wire  TLB_or9;
  wire  TLB_or10;
  wire  TLB_or4;
  wire  TLB_or1;
  wire  TLB_or11;
  wire  TLB_or12;
  wire  TLB_or5;
  wire  TLB_or13;
  wire  TLB_or14;
  wire  TLB_or6;
  wire  TLB_or2;
  wire  TLB_or0;
  reg  TLB_metaAssert;
  reg [31:0] _RAND_103;
  OptimizationBarrier mpu_ppn_barrier ( // @[package.scala 258:25]
    .io_x_ppn(mpu_ppn_barrier_io_x_ppn),
    .io_x_u(mpu_ppn_barrier_io_x_u),
    .io_x_ae(mpu_ppn_barrier_io_x_ae),
    .io_x_sw(mpu_ppn_barrier_io_x_sw),
    .io_x_sx(mpu_ppn_barrier_io_x_sx),
    .io_x_sr(mpu_ppn_barrier_io_x_sr),
    .io_x_pw(mpu_ppn_barrier_io_x_pw),
    .io_x_px(mpu_ppn_barrier_io_x_px),
    .io_x_pr(mpu_ppn_barrier_io_x_pr),
    .io_x_ppp(mpu_ppn_barrier_io_x_ppp),
    .io_x_pal(mpu_ppn_barrier_io_x_pal),
    .io_x_paa(mpu_ppn_barrier_io_x_paa),
    .io_x_eff(mpu_ppn_barrier_io_x_eff),
    .io_x_c(mpu_ppn_barrier_io_x_c),
    .io_y_ppn(mpu_ppn_barrier_io_y_ppn),
    .io_y_u(mpu_ppn_barrier_io_y_u),
    .io_y_ae(mpu_ppn_barrier_io_y_ae),
    .io_y_sw(mpu_ppn_barrier_io_y_sw),
    .io_y_sx(mpu_ppn_barrier_io_y_sx),
    .io_y_sr(mpu_ppn_barrier_io_y_sr),
    .io_y_pw(mpu_ppn_barrier_io_y_pw),
    .io_y_px(mpu_ppn_barrier_io_y_px),
    .io_y_pr(mpu_ppn_barrier_io_y_pr),
    .io_y_ppp(mpu_ppn_barrier_io_y_ppp),
    .io_y_pal(mpu_ppn_barrier_io_y_pal),
    .io_y_paa(mpu_ppn_barrier_io_y_paa),
    .io_y_eff(mpu_ppn_barrier_io_y_eff),
    .io_y_c(mpu_ppn_barrier_io_y_c),
    .io_covSum(mpu_ppn_barrier_io_covSum),
    .metaAssert(mpu_ppn_barrier_metaAssert)
  );
  PMPChecker pmp ( // @[TLB.scala 192:19]
    .io_prv(pmp_io_prv),
    .io_pmp_0_cfg_l(pmp_io_pmp_0_cfg_l),
    .io_pmp_0_cfg_a(pmp_io_pmp_0_cfg_a),
    .io_pmp_0_cfg_x(pmp_io_pmp_0_cfg_x),
    .io_pmp_0_cfg_w(pmp_io_pmp_0_cfg_w),
    .io_pmp_0_cfg_r(pmp_io_pmp_0_cfg_r),
    .io_pmp_0_addr(pmp_io_pmp_0_addr),
    .io_pmp_0_mask(pmp_io_pmp_0_mask),
    .io_pmp_1_cfg_l(pmp_io_pmp_1_cfg_l),
    .io_pmp_1_cfg_a(pmp_io_pmp_1_cfg_a),
    .io_pmp_1_cfg_x(pmp_io_pmp_1_cfg_x),
    .io_pmp_1_cfg_w(pmp_io_pmp_1_cfg_w),
    .io_pmp_1_cfg_r(pmp_io_pmp_1_cfg_r),
    .io_pmp_1_addr(pmp_io_pmp_1_addr),
    .io_pmp_1_mask(pmp_io_pmp_1_mask),
    .io_pmp_2_cfg_l(pmp_io_pmp_2_cfg_l),
    .io_pmp_2_cfg_a(pmp_io_pmp_2_cfg_a),
    .io_pmp_2_cfg_x(pmp_io_pmp_2_cfg_x),
    .io_pmp_2_cfg_w(pmp_io_pmp_2_cfg_w),
    .io_pmp_2_cfg_r(pmp_io_pmp_2_cfg_r),
    .io_pmp_2_addr(pmp_io_pmp_2_addr),
    .io_pmp_2_mask(pmp_io_pmp_2_mask),
    .io_pmp_3_cfg_l(pmp_io_pmp_3_cfg_l),
    .io_pmp_3_cfg_a(pmp_io_pmp_3_cfg_a),
    .io_pmp_3_cfg_x(pmp_io_pmp_3_cfg_x),
    .io_pmp_3_cfg_w(pmp_io_pmp_3_cfg_w),
    .io_pmp_3_cfg_r(pmp_io_pmp_3_cfg_r),
    .io_pmp_3_addr(pmp_io_pmp_3_addr),
    .io_pmp_3_mask(pmp_io_pmp_3_mask),
    .io_pmp_4_cfg_l(pmp_io_pmp_4_cfg_l),
    .io_pmp_4_cfg_a(pmp_io_pmp_4_cfg_a),
    .io_pmp_4_cfg_x(pmp_io_pmp_4_cfg_x),
    .io_pmp_4_cfg_w(pmp_io_pmp_4_cfg_w),
    .io_pmp_4_cfg_r(pmp_io_pmp_4_cfg_r),
    .io_pmp_4_addr(pmp_io_pmp_4_addr),
    .io_pmp_4_mask(pmp_io_pmp_4_mask),
    .io_pmp_5_cfg_l(pmp_io_pmp_5_cfg_l),
    .io_pmp_5_cfg_a(pmp_io_pmp_5_cfg_a),
    .io_pmp_5_cfg_x(pmp_io_pmp_5_cfg_x),
    .io_pmp_5_cfg_w(pmp_io_pmp_5_cfg_w),
    .io_pmp_5_cfg_r(pmp_io_pmp_5_cfg_r),
    .io_pmp_5_addr(pmp_io_pmp_5_addr),
    .io_pmp_5_mask(pmp_io_pmp_5_mask),
    .io_pmp_6_cfg_l(pmp_io_pmp_6_cfg_l),
    .io_pmp_6_cfg_a(pmp_io_pmp_6_cfg_a),
    .io_pmp_6_cfg_x(pmp_io_pmp_6_cfg_x),
    .io_pmp_6_cfg_w(pmp_io_pmp_6_cfg_w),
    .io_pmp_6_cfg_r(pmp_io_pmp_6_cfg_r),
    .io_pmp_6_addr(pmp_io_pmp_6_addr),
    .io_pmp_6_mask(pmp_io_pmp_6_mask),
    .io_pmp_7_cfg_l(pmp_io_pmp_7_cfg_l),
    .io_pmp_7_cfg_a(pmp_io_pmp_7_cfg_a),
    .io_pmp_7_cfg_x(pmp_io_pmp_7_cfg_x),
    .io_pmp_7_cfg_w(pmp_io_pmp_7_cfg_w),
    .io_pmp_7_cfg_r(pmp_io_pmp_7_cfg_r),
    .io_pmp_7_addr(pmp_io_pmp_7_addr),
    .io_pmp_7_mask(pmp_io_pmp_7_mask),
    .io_addr(pmp_io_addr),
    .io_size(pmp_io_size),
    .io_r(pmp_io_r),
    .io_w(pmp_io_w),
    .io_x(pmp_io_x),
    .io_covSum(pmp_io_covSum),
    .metaAssert(pmp_metaAssert)
  );
  OptimizationBarrier entries_barrier ( // @[package.scala 258:25]
    .io_x_ppn(entries_barrier_io_x_ppn),
    .io_x_u(entries_barrier_io_x_u),
    .io_x_ae(entries_barrier_io_x_ae),
    .io_x_sw(entries_barrier_io_x_sw),
    .io_x_sx(entries_barrier_io_x_sx),
    .io_x_sr(entries_barrier_io_x_sr),
    .io_x_pw(entries_barrier_io_x_pw),
    .io_x_px(entries_barrier_io_x_px),
    .io_x_pr(entries_barrier_io_x_pr),
    .io_x_ppp(entries_barrier_io_x_ppp),
    .io_x_pal(entries_barrier_io_x_pal),
    .io_x_paa(entries_barrier_io_x_paa),
    .io_x_eff(entries_barrier_io_x_eff),
    .io_x_c(entries_barrier_io_x_c),
    .io_y_ppn(entries_barrier_io_y_ppn),
    .io_y_u(entries_barrier_io_y_u),
    .io_y_ae(entries_barrier_io_y_ae),
    .io_y_sw(entries_barrier_io_y_sw),
    .io_y_sx(entries_barrier_io_y_sx),
    .io_y_sr(entries_barrier_io_y_sr),
    .io_y_pw(entries_barrier_io_y_pw),
    .io_y_px(entries_barrier_io_y_px),
    .io_y_pr(entries_barrier_io_y_pr),
    .io_y_ppp(entries_barrier_io_y_ppp),
    .io_y_pal(entries_barrier_io_y_pal),
    .io_y_paa(entries_barrier_io_y_paa),
    .io_y_eff(entries_barrier_io_y_eff),
    .io_y_c(entries_barrier_io_y_c),
    .io_covSum(entries_barrier_io_covSum),
    .metaAssert(entries_barrier_metaAssert)
  );
  OptimizationBarrier entries_barrier_1 ( // @[package.scala 258:25]
    .io_x_ppn(entries_barrier_1_io_x_ppn),
    .io_x_u(entries_barrier_1_io_x_u),
    .io_x_ae(entries_barrier_1_io_x_ae),
    .io_x_sw(entries_barrier_1_io_x_sw),
    .io_x_sx(entries_barrier_1_io_x_sx),
    .io_x_sr(entries_barrier_1_io_x_sr),
    .io_x_pw(entries_barrier_1_io_x_pw),
    .io_x_px(entries_barrier_1_io_x_px),
    .io_x_pr(entries_barrier_1_io_x_pr),
    .io_x_ppp(entries_barrier_1_io_x_ppp),
    .io_x_pal(entries_barrier_1_io_x_pal),
    .io_x_paa(entries_barrier_1_io_x_paa),
    .io_x_eff(entries_barrier_1_io_x_eff),
    .io_x_c(entries_barrier_1_io_x_c),
    .io_y_ppn(entries_barrier_1_io_y_ppn),
    .io_y_u(entries_barrier_1_io_y_u),
    .io_y_ae(entries_barrier_1_io_y_ae),
    .io_y_sw(entries_barrier_1_io_y_sw),
    .io_y_sx(entries_barrier_1_io_y_sx),
    .io_y_sr(entries_barrier_1_io_y_sr),
    .io_y_pw(entries_barrier_1_io_y_pw),
    .io_y_px(entries_barrier_1_io_y_px),
    .io_y_pr(entries_barrier_1_io_y_pr),
    .io_y_ppp(entries_barrier_1_io_y_ppp),
    .io_y_pal(entries_barrier_1_io_y_pal),
    .io_y_paa(entries_barrier_1_io_y_paa),
    .io_y_eff(entries_barrier_1_io_y_eff),
    .io_y_c(entries_barrier_1_io_y_c),
    .io_covSum(entries_barrier_1_io_covSum),
    .metaAssert(entries_barrier_1_metaAssert)
  );
  OptimizationBarrier entries_barrier_2 ( // @[package.scala 258:25]
    .io_x_ppn(entries_barrier_2_io_x_ppn),
    .io_x_u(entries_barrier_2_io_x_u),
    .io_x_ae(entries_barrier_2_io_x_ae),
    .io_x_sw(entries_barrier_2_io_x_sw),
    .io_x_sx(entries_barrier_2_io_x_sx),
    .io_x_sr(entries_barrier_2_io_x_sr),
    .io_x_pw(entries_barrier_2_io_x_pw),
    .io_x_px(entries_barrier_2_io_x_px),
    .io_x_pr(entries_barrier_2_io_x_pr),
    .io_x_ppp(entries_barrier_2_io_x_ppp),
    .io_x_pal(entries_barrier_2_io_x_pal),
    .io_x_paa(entries_barrier_2_io_x_paa),
    .io_x_eff(entries_barrier_2_io_x_eff),
    .io_x_c(entries_barrier_2_io_x_c),
    .io_y_ppn(entries_barrier_2_io_y_ppn),
    .io_y_u(entries_barrier_2_io_y_u),
    .io_y_ae(entries_barrier_2_io_y_ae),
    .io_y_sw(entries_barrier_2_io_y_sw),
    .io_y_sx(entries_barrier_2_io_y_sx),
    .io_y_sr(entries_barrier_2_io_y_sr),
    .io_y_pw(entries_barrier_2_io_y_pw),
    .io_y_px(entries_barrier_2_io_y_px),
    .io_y_pr(entries_barrier_2_io_y_pr),
    .io_y_ppp(entries_barrier_2_io_y_ppp),
    .io_y_pal(entries_barrier_2_io_y_pal),
    .io_y_paa(entries_barrier_2_io_y_paa),
    .io_y_eff(entries_barrier_2_io_y_eff),
    .io_y_c(entries_barrier_2_io_y_c),
    .io_covSum(entries_barrier_2_io_covSum),
    .metaAssert(entries_barrier_2_metaAssert)
  );
  OptimizationBarrier entries_barrier_3 ( // @[package.scala 258:25]
    .io_x_ppn(entries_barrier_3_io_x_ppn),
    .io_x_u(entries_barrier_3_io_x_u),
    .io_x_ae(entries_barrier_3_io_x_ae),
    .io_x_sw(entries_barrier_3_io_x_sw),
    .io_x_sx(entries_barrier_3_io_x_sx),
    .io_x_sr(entries_barrier_3_io_x_sr),
    .io_x_pw(entries_barrier_3_io_x_pw),
    .io_x_px(entries_barrier_3_io_x_px),
    .io_x_pr(entries_barrier_3_io_x_pr),
    .io_x_ppp(entries_barrier_3_io_x_ppp),
    .io_x_pal(entries_barrier_3_io_x_pal),
    .io_x_paa(entries_barrier_3_io_x_paa),
    .io_x_eff(entries_barrier_3_io_x_eff),
    .io_x_c(entries_barrier_3_io_x_c),
    .io_y_ppn(entries_barrier_3_io_y_ppn),
    .io_y_u(entries_barrier_3_io_y_u),
    .io_y_ae(entries_barrier_3_io_y_ae),
    .io_y_sw(entries_barrier_3_io_y_sw),
    .io_y_sx(entries_barrier_3_io_y_sx),
    .io_y_sr(entries_barrier_3_io_y_sr),
    .io_y_pw(entries_barrier_3_io_y_pw),
    .io_y_px(entries_barrier_3_io_y_px),
    .io_y_pr(entries_barrier_3_io_y_pr),
    .io_y_ppp(entries_barrier_3_io_y_ppp),
    .io_y_pal(entries_barrier_3_io_y_pal),
    .io_y_paa(entries_barrier_3_io_y_paa),
    .io_y_eff(entries_barrier_3_io_y_eff),
    .io_y_c(entries_barrier_3_io_y_c),
    .io_covSum(entries_barrier_3_io_covSum),
    .metaAssert(entries_barrier_3_metaAssert)
  );
  OptimizationBarrier entries_barrier_4 ( // @[package.scala 258:25]
    .io_x_ppn(entries_barrier_4_io_x_ppn),
    .io_x_u(entries_barrier_4_io_x_u),
    .io_x_ae(entries_barrier_4_io_x_ae),
    .io_x_sw(entries_barrier_4_io_x_sw),
    .io_x_sx(entries_barrier_4_io_x_sx),
    .io_x_sr(entries_barrier_4_io_x_sr),
    .io_x_pw(entries_barrier_4_io_x_pw),
    .io_x_px(entries_barrier_4_io_x_px),
    .io_x_pr(entries_barrier_4_io_x_pr),
    .io_x_ppp(entries_barrier_4_io_x_ppp),
    .io_x_pal(entries_barrier_4_io_x_pal),
    .io_x_paa(entries_barrier_4_io_x_paa),
    .io_x_eff(entries_barrier_4_io_x_eff),
    .io_x_c(entries_barrier_4_io_x_c),
    .io_y_ppn(entries_barrier_4_io_y_ppn),
    .io_y_u(entries_barrier_4_io_y_u),
    .io_y_ae(entries_barrier_4_io_y_ae),
    .io_y_sw(entries_barrier_4_io_y_sw),
    .io_y_sx(entries_barrier_4_io_y_sx),
    .io_y_sr(entries_barrier_4_io_y_sr),
    .io_y_pw(entries_barrier_4_io_y_pw),
    .io_y_px(entries_barrier_4_io_y_px),
    .io_y_pr(entries_barrier_4_io_y_pr),
    .io_y_ppp(entries_barrier_4_io_y_ppp),
    .io_y_pal(entries_barrier_4_io_y_pal),
    .io_y_paa(entries_barrier_4_io_y_paa),
    .io_y_eff(entries_barrier_4_io_y_eff),
    .io_y_c(entries_barrier_4_io_y_c),
    .io_covSum(entries_barrier_4_io_covSum),
    .metaAssert(entries_barrier_4_metaAssert)
  );
  OptimizationBarrier entries_barrier_5 ( // @[package.scala 258:25]
    .io_x_ppn(entries_barrier_5_io_x_ppn),
    .io_x_u(entries_barrier_5_io_x_u),
    .io_x_ae(entries_barrier_5_io_x_ae),
    .io_x_sw(entries_barrier_5_io_x_sw),
    .io_x_sx(entries_barrier_5_io_x_sx),
    .io_x_sr(entries_barrier_5_io_x_sr),
    .io_x_pw(entries_barrier_5_io_x_pw),
    .io_x_px(entries_barrier_5_io_x_px),
    .io_x_pr(entries_barrier_5_io_x_pr),
    .io_x_ppp(entries_barrier_5_io_x_ppp),
    .io_x_pal(entries_barrier_5_io_x_pal),
    .io_x_paa(entries_barrier_5_io_x_paa),
    .io_x_eff(entries_barrier_5_io_x_eff),
    .io_x_c(entries_barrier_5_io_x_c),
    .io_y_ppn(entries_barrier_5_io_y_ppn),
    .io_y_u(entries_barrier_5_io_y_u),
    .io_y_ae(entries_barrier_5_io_y_ae),
    .io_y_sw(entries_barrier_5_io_y_sw),
    .io_y_sx(entries_barrier_5_io_y_sx),
    .io_y_sr(entries_barrier_5_io_y_sr),
    .io_y_pw(entries_barrier_5_io_y_pw),
    .io_y_px(entries_barrier_5_io_y_px),
    .io_y_pr(entries_barrier_5_io_y_pr),
    .io_y_ppp(entries_barrier_5_io_y_ppp),
    .io_y_pal(entries_barrier_5_io_y_pal),
    .io_y_paa(entries_barrier_5_io_y_paa),
    .io_y_eff(entries_barrier_5_io_y_eff),
    .io_y_c(entries_barrier_5_io_y_c),
    .io_covSum(entries_barrier_5_io_covSum),
    .metaAssert(entries_barrier_5_metaAssert)
  );
  OptimizationBarrier entries_barrier_6 ( // @[package.scala 258:25]
    .io_x_ppn(entries_barrier_6_io_x_ppn),
    .io_x_u(entries_barrier_6_io_x_u),
    .io_x_ae(entries_barrier_6_io_x_ae),
    .io_x_sw(entries_barrier_6_io_x_sw),
    .io_x_sx(entries_barrier_6_io_x_sx),
    .io_x_sr(entries_barrier_6_io_x_sr),
    .io_x_pw(entries_barrier_6_io_x_pw),
    .io_x_px(entries_barrier_6_io_x_px),
    .io_x_pr(entries_barrier_6_io_x_pr),
    .io_x_ppp(entries_barrier_6_io_x_ppp),
    .io_x_pal(entries_barrier_6_io_x_pal),
    .io_x_paa(entries_barrier_6_io_x_paa),
    .io_x_eff(entries_barrier_6_io_x_eff),
    .io_x_c(entries_barrier_6_io_x_c),
    .io_y_ppn(entries_barrier_6_io_y_ppn),
    .io_y_u(entries_barrier_6_io_y_u),
    .io_y_ae(entries_barrier_6_io_y_ae),
    .io_y_sw(entries_barrier_6_io_y_sw),
    .io_y_sx(entries_barrier_6_io_y_sx),
    .io_y_sr(entries_barrier_6_io_y_sr),
    .io_y_pw(entries_barrier_6_io_y_pw),
    .io_y_px(entries_barrier_6_io_y_px),
    .io_y_pr(entries_barrier_6_io_y_pr),
    .io_y_ppp(entries_barrier_6_io_y_ppp),
    .io_y_pal(entries_barrier_6_io_y_pal),
    .io_y_paa(entries_barrier_6_io_y_paa),
    .io_y_eff(entries_barrier_6_io_y_eff),
    .io_y_c(entries_barrier_6_io_y_c),
    .io_covSum(entries_barrier_6_io_covSum),
    .metaAssert(entries_barrier_6_metaAssert)
  );
  OptimizationBarrier entries_barrier_7 ( // @[package.scala 258:25]
    .io_x_ppn(entries_barrier_7_io_x_ppn),
    .io_x_u(entries_barrier_7_io_x_u),
    .io_x_ae(entries_barrier_7_io_x_ae),
    .io_x_sw(entries_barrier_7_io_x_sw),
    .io_x_sx(entries_barrier_7_io_x_sx),
    .io_x_sr(entries_barrier_7_io_x_sr),
    .io_x_pw(entries_barrier_7_io_x_pw),
    .io_x_px(entries_barrier_7_io_x_px),
    .io_x_pr(entries_barrier_7_io_x_pr),
    .io_x_ppp(entries_barrier_7_io_x_ppp),
    .io_x_pal(entries_barrier_7_io_x_pal),
    .io_x_paa(entries_barrier_7_io_x_paa),
    .io_x_eff(entries_barrier_7_io_x_eff),
    .io_x_c(entries_barrier_7_io_x_c),
    .io_y_ppn(entries_barrier_7_io_y_ppn),
    .io_y_u(entries_barrier_7_io_y_u),
    .io_y_ae(entries_barrier_7_io_y_ae),
    .io_y_sw(entries_barrier_7_io_y_sw),
    .io_y_sx(entries_barrier_7_io_y_sx),
    .io_y_sr(entries_barrier_7_io_y_sr),
    .io_y_pw(entries_barrier_7_io_y_pw),
    .io_y_px(entries_barrier_7_io_y_px),
    .io_y_pr(entries_barrier_7_io_y_pr),
    .io_y_ppp(entries_barrier_7_io_y_ppp),
    .io_y_pal(entries_barrier_7_io_y_pal),
    .io_y_paa(entries_barrier_7_io_y_paa),
    .io_y_eff(entries_barrier_7_io_y_eff),
    .io_y_c(entries_barrier_7_io_y_c),
    .io_covSum(entries_barrier_7_io_covSum),
    .metaAssert(entries_barrier_7_metaAssert)
  );
  OptimizationBarrier entries_barrier_8 ( // @[package.scala 258:25]
    .io_x_ppn(entries_barrier_8_io_x_ppn),
    .io_x_u(entries_barrier_8_io_x_u),
    .io_x_ae(entries_barrier_8_io_x_ae),
    .io_x_sw(entries_barrier_8_io_x_sw),
    .io_x_sx(entries_barrier_8_io_x_sx),
    .io_x_sr(entries_barrier_8_io_x_sr),
    .io_x_pw(entries_barrier_8_io_x_pw),
    .io_x_px(entries_barrier_8_io_x_px),
    .io_x_pr(entries_barrier_8_io_x_pr),
    .io_x_ppp(entries_barrier_8_io_x_ppp),
    .io_x_pal(entries_barrier_8_io_x_pal),
    .io_x_paa(entries_barrier_8_io_x_paa),
    .io_x_eff(entries_barrier_8_io_x_eff),
    .io_x_c(entries_barrier_8_io_x_c),
    .io_y_ppn(entries_barrier_8_io_y_ppn),
    .io_y_u(entries_barrier_8_io_y_u),
    .io_y_ae(entries_barrier_8_io_y_ae),
    .io_y_sw(entries_barrier_8_io_y_sw),
    .io_y_sx(entries_barrier_8_io_y_sx),
    .io_y_sr(entries_barrier_8_io_y_sr),
    .io_y_pw(entries_barrier_8_io_y_pw),
    .io_y_px(entries_barrier_8_io_y_px),
    .io_y_pr(entries_barrier_8_io_y_pr),
    .io_y_ppp(entries_barrier_8_io_y_ppp),
    .io_y_pal(entries_barrier_8_io_y_pal),
    .io_y_paa(entries_barrier_8_io_y_paa),
    .io_y_eff(entries_barrier_8_io_y_eff),
    .io_y_c(entries_barrier_8_io_y_c),
    .io_covSum(entries_barrier_8_io_covSum),
    .metaAssert(entries_barrier_8_metaAssert)
  );
  OptimizationBarrier entries_barrier_9 ( // @[package.scala 258:25]
    .io_x_ppn(entries_barrier_9_io_x_ppn),
    .io_x_u(entries_barrier_9_io_x_u),
    .io_x_ae(entries_barrier_9_io_x_ae),
    .io_x_sw(entries_barrier_9_io_x_sw),
    .io_x_sx(entries_barrier_9_io_x_sx),
    .io_x_sr(entries_barrier_9_io_x_sr),
    .io_x_pw(entries_barrier_9_io_x_pw),
    .io_x_px(entries_barrier_9_io_x_px),
    .io_x_pr(entries_barrier_9_io_x_pr),
    .io_x_ppp(entries_barrier_9_io_x_ppp),
    .io_x_pal(entries_barrier_9_io_x_pal),
    .io_x_paa(entries_barrier_9_io_x_paa),
    .io_x_eff(entries_barrier_9_io_x_eff),
    .io_x_c(entries_barrier_9_io_x_c),
    .io_y_ppn(entries_barrier_9_io_y_ppn),
    .io_y_u(entries_barrier_9_io_y_u),
    .io_y_ae(entries_barrier_9_io_y_ae),
    .io_y_sw(entries_barrier_9_io_y_sw),
    .io_y_sx(entries_barrier_9_io_y_sx),
    .io_y_sr(entries_barrier_9_io_y_sr),
    .io_y_pw(entries_barrier_9_io_y_pw),
    .io_y_px(entries_barrier_9_io_y_px),
    .io_y_pr(entries_barrier_9_io_y_pr),
    .io_y_ppp(entries_barrier_9_io_y_ppp),
    .io_y_pal(entries_barrier_9_io_y_pal),
    .io_y_paa(entries_barrier_9_io_y_paa),
    .io_y_eff(entries_barrier_9_io_y_eff),
    .io_y_c(entries_barrier_9_io_y_c),
    .io_covSum(entries_barrier_9_io_covSum),
    .metaAssert(entries_barrier_9_metaAssert)
  );
  OptimizationBarrier entries_barrier_10 ( // @[package.scala 258:25]
    .io_x_ppn(entries_barrier_10_io_x_ppn),
    .io_x_u(entries_barrier_10_io_x_u),
    .io_x_ae(entries_barrier_10_io_x_ae),
    .io_x_sw(entries_barrier_10_io_x_sw),
    .io_x_sx(entries_barrier_10_io_x_sx),
    .io_x_sr(entries_barrier_10_io_x_sr),
    .io_x_pw(entries_barrier_10_io_x_pw),
    .io_x_px(entries_barrier_10_io_x_px),
    .io_x_pr(entries_barrier_10_io_x_pr),
    .io_x_ppp(entries_barrier_10_io_x_ppp),
    .io_x_pal(entries_barrier_10_io_x_pal),
    .io_x_paa(entries_barrier_10_io_x_paa),
    .io_x_eff(entries_barrier_10_io_x_eff),
    .io_x_c(entries_barrier_10_io_x_c),
    .io_y_ppn(entries_barrier_10_io_y_ppn),
    .io_y_u(entries_barrier_10_io_y_u),
    .io_y_ae(entries_barrier_10_io_y_ae),
    .io_y_sw(entries_barrier_10_io_y_sw),
    .io_y_sx(entries_barrier_10_io_y_sx),
    .io_y_sr(entries_barrier_10_io_y_sr),
    .io_y_pw(entries_barrier_10_io_y_pw),
    .io_y_px(entries_barrier_10_io_y_px),
    .io_y_pr(entries_barrier_10_io_y_pr),
    .io_y_ppp(entries_barrier_10_io_y_ppp),
    .io_y_pal(entries_barrier_10_io_y_pal),
    .io_y_paa(entries_barrier_10_io_y_paa),
    .io_y_eff(entries_barrier_10_io_y_eff),
    .io_y_c(entries_barrier_10_io_y_c),
    .io_covSum(entries_barrier_10_io_covSum),
    .metaAssert(entries_barrier_10_metaAssert)
  );
  OptimizationBarrier entries_barrier_11 ( // @[package.scala 258:25]
    .io_x_ppn(entries_barrier_11_io_x_ppn),
    .io_x_u(entries_barrier_11_io_x_u),
    .io_x_ae(entries_barrier_11_io_x_ae),
    .io_x_sw(entries_barrier_11_io_x_sw),
    .io_x_sx(entries_barrier_11_io_x_sx),
    .io_x_sr(entries_barrier_11_io_x_sr),
    .io_x_pw(entries_barrier_11_io_x_pw),
    .io_x_px(entries_barrier_11_io_x_px),
    .io_x_pr(entries_barrier_11_io_x_pr),
    .io_x_ppp(entries_barrier_11_io_x_ppp),
    .io_x_pal(entries_barrier_11_io_x_pal),
    .io_x_paa(entries_barrier_11_io_x_paa),
    .io_x_eff(entries_barrier_11_io_x_eff),
    .io_x_c(entries_barrier_11_io_x_c),
    .io_y_ppn(entries_barrier_11_io_y_ppn),
    .io_y_u(entries_barrier_11_io_y_u),
    .io_y_ae(entries_barrier_11_io_y_ae),
    .io_y_sw(entries_barrier_11_io_y_sw),
    .io_y_sx(entries_barrier_11_io_y_sx),
    .io_y_sr(entries_barrier_11_io_y_sr),
    .io_y_pw(entries_barrier_11_io_y_pw),
    .io_y_px(entries_barrier_11_io_y_px),
    .io_y_pr(entries_barrier_11_io_y_pr),
    .io_y_ppp(entries_barrier_11_io_y_ppp),
    .io_y_pal(entries_barrier_11_io_y_pal),
    .io_y_paa(entries_barrier_11_io_y_paa),
    .io_y_eff(entries_barrier_11_io_y_eff),
    .io_y_c(entries_barrier_11_io_y_c),
    .io_covSum(entries_barrier_11_io_covSum),
    .metaAssert(entries_barrier_11_metaAssert)
  );
  OptimizationBarrier entries_barrier_12 ( // @[package.scala 258:25]
    .io_x_ppn(entries_barrier_12_io_x_ppn),
    .io_x_u(entries_barrier_12_io_x_u),
    .io_x_ae(entries_barrier_12_io_x_ae),
    .io_x_sw(entries_barrier_12_io_x_sw),
    .io_x_sx(entries_barrier_12_io_x_sx),
    .io_x_sr(entries_barrier_12_io_x_sr),
    .io_x_pw(entries_barrier_12_io_x_pw),
    .io_x_px(entries_barrier_12_io_x_px),
    .io_x_pr(entries_barrier_12_io_x_pr),
    .io_x_ppp(entries_barrier_12_io_x_ppp),
    .io_x_pal(entries_barrier_12_io_x_pal),
    .io_x_paa(entries_barrier_12_io_x_paa),
    .io_x_eff(entries_barrier_12_io_x_eff),
    .io_x_c(entries_barrier_12_io_x_c),
    .io_y_ppn(entries_barrier_12_io_y_ppn),
    .io_y_u(entries_barrier_12_io_y_u),
    .io_y_ae(entries_barrier_12_io_y_ae),
    .io_y_sw(entries_barrier_12_io_y_sw),
    .io_y_sx(entries_barrier_12_io_y_sx),
    .io_y_sr(entries_barrier_12_io_y_sr),
    .io_y_pw(entries_barrier_12_io_y_pw),
    .io_y_px(entries_barrier_12_io_y_px),
    .io_y_pr(entries_barrier_12_io_y_pr),
    .io_y_ppp(entries_barrier_12_io_y_ppp),
    .io_y_pal(entries_barrier_12_io_y_pal),
    .io_y_paa(entries_barrier_12_io_y_paa),
    .io_y_eff(entries_barrier_12_io_y_eff),
    .io_y_c(entries_barrier_12_io_y_c),
    .io_covSum(entries_barrier_12_io_covSum),
    .metaAssert(entries_barrier_12_metaAssert)
  );
  assign vpn = io_req_bits_vaddr[38:12]; // @[TLB.scala 162:30]
  assign priv_s = io_ptw_status_dprv[0]; // @[TLB.scala 180:20]
  assign priv_uses_vm = io_ptw_status_dprv <= 2'h1; // @[TLB.scala 181:27]
  assign _vm_enabled_T_2 = io_ptw_ptbr_mode[3] & priv_uses_vm; // @[TLB.scala 182:83]
  assign vm_enabled = _vm_enabled_T_2 & ~io_req_bits_passthrough; // @[TLB.scala 182:99]
  assign refill_ppn = io_ptw_resp_bits_pte_ppn[19:0]; // @[TLB.scala 185:44]
  assign _invalidate_refill_T = state == 2'h1; // @[package.scala 15:47]
  assign _invalidate_refill_T_1 = state == 2'h3; // @[package.scala 15:47]
  assign _invalidate_refill_T_2 = _invalidate_refill_T | _invalidate_refill_T_1; // @[package.scala 72:59]
  assign invalidate_refill = _invalidate_refill_T_2 | io_sfence_valid; // @[TLB.scala 187:88]
  assign mpu_ppn_hi = mpu_ppn_barrier_io_y_ppn[19:18]; // @[TLB.scala 105:26]
  assign mpu_ppn_ignore = special_entry_level < 2'h1; // @[TLB.scala 107:28]
  assign _mpu_ppn_T_17 = mpu_ppn_ignore ? vpn : 27'h0; // @[TLB.scala 108:28]
  assign _GEN_919 = {{7'd0}, mpu_ppn_barrier_io_y_ppn}; // @[TLB.scala 108:47]
  assign _mpu_ppn_T_18 = _mpu_ppn_T_17 | _GEN_919; // @[TLB.scala 108:47]
  assign mpu_ppn_lo = _mpu_ppn_T_18[17:9]; // @[TLB.scala 108:58]
  assign mpu_ppn_ignore_1 = special_entry_level < 2'h2; // @[TLB.scala 107:28]
  assign _mpu_ppn_T_19 = mpu_ppn_ignore_1 ? vpn : 27'h0; // @[TLB.scala 108:28]
  assign _mpu_ppn_T_20 = _mpu_ppn_T_19 | _GEN_919; // @[TLB.scala 108:47]
  assign mpu_ppn_lo_1 = _mpu_ppn_T_20[8:0]; // @[TLB.scala 108:58]
  assign _mpu_ppn_T_21 = {mpu_ppn_hi,mpu_ppn_lo,mpu_ppn_lo_1}; // @[Cat.scala 30:58]
  assign _mpu_ppn_T_23 = vm_enabled ? {{8'd0}, _mpu_ppn_T_21} : io_req_bits_vaddr[39:12]; // @[TLB.scala 189:20]
  assign mpu_ppn = io_ptw_resp_valid ? {{8'd0}, refill_ppn} : _mpu_ppn_T_23; // @[TLB.scala 188:20]
  assign mpu_physaddr_lo = io_req_bits_vaddr[11:0]; // @[TLB.scala 190:52]
  assign mpu_physaddr = {mpu_ppn,mpu_physaddr_lo}; // @[Cat.scala 30:58]
  assign _mpu_priv_T = io_ptw_resp_valid | io_req_bits_passthrough; // @[TLB.scala 191:56]
  assign _mpu_priv_T_2 = {io_ptw_status_debug,io_ptw_status_dprv}; // @[Cat.scala 30:58]
  assign mpu_priv = _mpu_priv_T ? 3'h1 : _mpu_priv_T_2; // @[TLB.scala 191:27]
  assign _legal_address_T = mpu_physaddr ^ 40'h3000; // @[Parameters.scala 137:31]
  assign _legal_address_T_1 = {1'b0,$signed(_legal_address_T)}; // @[Parameters.scala 137:49]
  assign _legal_address_T_3 = $signed(_legal_address_T_1) & -41'sh1000; // @[Parameters.scala 137:52]
  assign _legal_address_T_4 = $signed(_legal_address_T_3) == 41'sh0; // @[Parameters.scala 137:67]
  assign _legal_address_T_5 = mpu_physaddr ^ 40'hc000000; // @[Parameters.scala 137:31]
  assign _legal_address_T_6 = {1'b0,$signed(_legal_address_T_5)}; // @[Parameters.scala 137:49]
  assign _legal_address_T_8 = $signed(_legal_address_T_6) & -41'sh4000000; // @[Parameters.scala 137:52]
  assign _legal_address_T_9 = $signed(_legal_address_T_8) == 41'sh0; // @[Parameters.scala 137:67]
  assign _legal_address_T_10 = mpu_physaddr ^ 40'h2000000; // @[Parameters.scala 137:31]
  assign _legal_address_T_11 = {1'b0,$signed(_legal_address_T_10)}; // @[Parameters.scala 137:49]
  assign _legal_address_T_13 = $signed(_legal_address_T_11) & -41'sh10000; // @[Parameters.scala 137:52]
  assign _legal_address_T_14 = $signed(_legal_address_T_13) == 41'sh0; // @[Parameters.scala 137:67]
  assign _legal_address_T_16 = {1'b0,$signed(mpu_physaddr)}; // @[Parameters.scala 137:49]
  assign _legal_address_T_18 = $signed(_legal_address_T_16) & -41'sh1000; // @[Parameters.scala 137:52]
  assign _legal_address_T_19 = $signed(_legal_address_T_18) == 41'sh0; // @[Parameters.scala 137:67]
  assign _legal_address_T_20 = mpu_physaddr ^ 40'h10000; // @[Parameters.scala 137:31]
  assign _legal_address_T_21 = {1'b0,$signed(_legal_address_T_20)}; // @[Parameters.scala 137:49]
  assign _legal_address_T_23 = $signed(_legal_address_T_21) & -41'sh10000; // @[Parameters.scala 137:52]
  assign _legal_address_T_24 = $signed(_legal_address_T_23) == 41'sh0; // @[Parameters.scala 137:67]
  assign _legal_address_T_25 = mpu_physaddr ^ 40'h80000000; // @[Parameters.scala 137:31]
  assign _legal_address_T_26 = {1'b0,$signed(_legal_address_T_25)}; // @[Parameters.scala 137:49]
  assign _legal_address_T_28 = $signed(_legal_address_T_26) & -41'sh10000000; // @[Parameters.scala 137:52]
  assign _legal_address_T_29 = $signed(_legal_address_T_28) == 41'sh0; // @[Parameters.scala 137:67]
  assign _legal_address_T_30 = mpu_physaddr ^ 40'h60000000; // @[Parameters.scala 137:31]
  assign _legal_address_T_31 = {1'b0,$signed(_legal_address_T_30)}; // @[Parameters.scala 137:49]
  assign _legal_address_T_33 = $signed(_legal_address_T_31) & -41'sh20000000; // @[Parameters.scala 137:52]
  assign _legal_address_T_34 = $signed(_legal_address_T_33) == 41'sh0; // @[Parameters.scala 137:67]
  assign _legal_address_T_35 = _legal_address_T_4 | _legal_address_T_9; // @[TLB.scala 197:67]
  assign _legal_address_T_36 = _legal_address_T_35 | _legal_address_T_14; // @[TLB.scala 197:67]
  assign _legal_address_T_37 = _legal_address_T_36 | _legal_address_T_19; // @[TLB.scala 197:67]
  assign _legal_address_T_38 = _legal_address_T_37 | _legal_address_T_24; // @[TLB.scala 197:67]
  assign _legal_address_T_39 = _legal_address_T_38 | _legal_address_T_29; // @[TLB.scala 197:67]
  assign legal_address = _legal_address_T_39 | _legal_address_T_34; // @[TLB.scala 197:67]
  assign _cacheable_T_8 = $signed(_legal_address_T_26) & 41'sh80000000; // @[Parameters.scala 137:52]
  assign _cacheable_T_9 = $signed(_cacheable_T_8) == 41'sh0; // @[Parameters.scala 137:67]
  assign cacheable = legal_address & _cacheable_T_9; // @[TLB.scala 199:19]
  assign _homogeneous_T_54 = mpu_physaddr ^ 40'h8000000; // @[Parameters.scala 137:31]
  assign _homogeneous_T_55 = {1'b0,$signed(_homogeneous_T_54)}; // @[Parameters.scala 137:49]
  assign _homogeneous_T_57 = $signed(_homogeneous_T_55) & 41'shc8000000; // @[Parameters.scala 137:52]
  assign _homogeneous_T_58 = $signed(_homogeneous_T_57) == 41'sh0; // @[Parameters.scala 137:67]
  assign _homogeneous_T_71 = $signed(_legal_address_T_16) & 41'shc8010000; // @[Parameters.scala 137:52]
  assign _homogeneous_T_72 = $signed(_homogeneous_T_71) == 41'sh0; // @[Parameters.scala 137:67]
  assign _homogeneous_T_79 = _homogeneous_T_72 | _homogeneous_T_58; // @[TLBPermissions.scala 83:66]
  assign _deny_access_to_debug_T = mpu_priv <= 3'h3; // @[TLB.scala 202:39]
  assign deny_access_to_debug = _deny_access_to_debug_T & _legal_address_T_19; // @[TLB.scala 202:48]
  assign _prot_r_T_7 = legal_address & ~deny_access_to_debug; // @[TLB.scala 203:41]
  assign prot_r = _prot_r_T_7 & pmp_io_r; // @[TLB.scala 203:66]
  assign _prot_w_T_10 = mpu_physaddr ^ 40'h40000000; // @[Parameters.scala 137:31]
  assign _prot_w_T_11 = {1'b0,$signed(_prot_w_T_10)}; // @[Parameters.scala 137:49]
  assign _prot_w_T_13 = $signed(_prot_w_T_11) & 41'shc0000000; // @[Parameters.scala 137:52]
  assign _prot_w_T_14 = $signed(_prot_w_T_13) == 41'sh0; // @[Parameters.scala 137:67]
  assign _prot_w_T_18 = $signed(_legal_address_T_26) & 41'shc0000000; // @[Parameters.scala 137:52]
  assign _prot_w_T_19 = $signed(_prot_w_T_18) == 41'sh0; // @[Parameters.scala 137:67]
  assign _prot_w_T_21 = _homogeneous_T_79 | _prot_w_T_14; // @[Parameters.scala 615:89]
  assign _prot_w_T_22 = _prot_w_T_21 | _prot_w_T_19; // @[Parameters.scala 615:89]
  assign _prot_w_T_31 = legal_address & _prot_w_T_22; // @[TLB.scala 199:19]
  assign _prot_w_T_33 = _prot_w_T_31 & ~deny_access_to_debug; // @[TLB.scala 204:45]
  assign prot_w = _prot_w_T_33 & pmp_io_w; // @[TLB.scala 204:70]
  assign prot_al = legal_address & _homogeneous_T_79; // @[TLB.scala 199:19]
  assign _prot_x_T_3 = $signed(_legal_address_T_16) & 41'shca000000; // @[Parameters.scala 137:52]
  assign _prot_x_T_4 = $signed(_prot_x_T_3) == 41'sh0; // @[Parameters.scala 137:67]
  assign _prot_x_T_15 = _prot_x_T_4 | _prot_w_T_14; // @[Parameters.scala 615:89]
  assign _prot_x_T_16 = _prot_x_T_15 | _prot_w_T_19; // @[Parameters.scala 615:89]
  assign _prot_x_T_31 = legal_address & _prot_x_T_16; // @[TLB.scala 199:19]
  assign _prot_x_T_33 = _prot_x_T_31 & ~deny_access_to_debug; // @[TLB.scala 208:40]
  assign prot_x = _prot_x_T_33 & pmp_io_x; // @[TLB.scala 208:65]
  assign _prot_eff_T_20 = $signed(_legal_address_T_16) & 41'shca012000; // @[Parameters.scala 137:52]
  assign _prot_eff_T_21 = $signed(_prot_eff_T_20) == 41'sh0; // @[Parameters.scala 137:67]
  assign _prot_eff_T_25 = $signed(_legal_address_T_11) & 41'shca010000; // @[Parameters.scala 137:52]
  assign _prot_eff_T_26 = $signed(_prot_eff_T_25) == 41'sh0; // @[Parameters.scala 137:67]
  assign _prot_eff_T_37 = _prot_eff_T_21 | _prot_eff_T_26; // @[Parameters.scala 615:89]
  assign _prot_eff_T_38 = _prot_eff_T_37 | _homogeneous_T_58; // @[Parameters.scala 615:89]
  assign _prot_eff_T_39 = _prot_eff_T_38 | _prot_w_T_14; // @[Parameters.scala 615:89]
  assign prot_eff = legal_address & _prot_eff_T_39; // @[TLB.scala 199:19]
  assign _sector_hits_T = sectored_entries_0_0_valid_0 | sectored_entries_0_0_valid_1; // @[package.scala 72:59]
  assign _sector_hits_T_1 = _sector_hits_T | sectored_entries_0_0_valid_2; // @[package.scala 72:59]
  assign _sector_hits_T_2 = _sector_hits_T_1 | sectored_entries_0_0_valid_3; // @[package.scala 72:59]
  assign _sector_hits_T_3 = sectored_entries_0_0_tag ^ vpn; // @[TLB.scala 88:41]
  assign _sector_hits_T_5 = _sector_hits_T_3[26:2] == 25'h0; // @[TLB.scala 88:66]
  assign sector_hits_0 = _sector_hits_T_2 & _sector_hits_T_5; // @[TLB.scala 87:40]
  assign _sector_hits_T_6 = sectored_entries_0_1_valid_0 | sectored_entries_0_1_valid_1; // @[package.scala 72:59]
  assign _sector_hits_T_7 = _sector_hits_T_6 | sectored_entries_0_1_valid_2; // @[package.scala 72:59]
  assign _sector_hits_T_8 = _sector_hits_T_7 | sectored_entries_0_1_valid_3; // @[package.scala 72:59]
  assign _sector_hits_T_9 = sectored_entries_0_1_tag ^ vpn; // @[TLB.scala 88:41]
  assign _sector_hits_T_11 = _sector_hits_T_9[26:2] == 25'h0; // @[TLB.scala 88:66]
  assign sector_hits_1 = _sector_hits_T_8 & _sector_hits_T_11; // @[TLB.scala 87:40]
  assign _sector_hits_T_12 = sectored_entries_0_2_valid_0 | sectored_entries_0_2_valid_1; // @[package.scala 72:59]
  assign _sector_hits_T_13 = _sector_hits_T_12 | sectored_entries_0_2_valid_2; // @[package.scala 72:59]
  assign _sector_hits_T_14 = _sector_hits_T_13 | sectored_entries_0_2_valid_3; // @[package.scala 72:59]
  assign _sector_hits_T_15 = sectored_entries_0_2_tag ^ vpn; // @[TLB.scala 88:41]
  assign _sector_hits_T_17 = _sector_hits_T_15[26:2] == 25'h0; // @[TLB.scala 88:66]
  assign sector_hits_2 = _sector_hits_T_14 & _sector_hits_T_17; // @[TLB.scala 87:40]
  assign _sector_hits_T_18 = sectored_entries_0_3_valid_0 | sectored_entries_0_3_valid_1; // @[package.scala 72:59]
  assign _sector_hits_T_19 = _sector_hits_T_18 | sectored_entries_0_3_valid_2; // @[package.scala 72:59]
  assign _sector_hits_T_20 = _sector_hits_T_19 | sectored_entries_0_3_valid_3; // @[package.scala 72:59]
  assign _sector_hits_T_21 = sectored_entries_0_3_tag ^ vpn; // @[TLB.scala 88:41]
  assign _sector_hits_T_23 = _sector_hits_T_21[26:2] == 25'h0; // @[TLB.scala 88:66]
  assign sector_hits_3 = _sector_hits_T_20 & _sector_hits_T_23; // @[TLB.scala 87:40]
  assign _sector_hits_T_24 = sectored_entries_0_4_valid_0 | sectored_entries_0_4_valid_1; // @[package.scala 72:59]
  assign _sector_hits_T_25 = _sector_hits_T_24 | sectored_entries_0_4_valid_2; // @[package.scala 72:59]
  assign _sector_hits_T_26 = _sector_hits_T_25 | sectored_entries_0_4_valid_3; // @[package.scala 72:59]
  assign _sector_hits_T_27 = sectored_entries_0_4_tag ^ vpn; // @[TLB.scala 88:41]
  assign _sector_hits_T_29 = _sector_hits_T_27[26:2] == 25'h0; // @[TLB.scala 88:66]
  assign sector_hits_4 = _sector_hits_T_26 & _sector_hits_T_29; // @[TLB.scala 87:40]
  assign _sector_hits_T_30 = sectored_entries_0_5_valid_0 | sectored_entries_0_5_valid_1; // @[package.scala 72:59]
  assign _sector_hits_T_31 = _sector_hits_T_30 | sectored_entries_0_5_valid_2; // @[package.scala 72:59]
  assign _sector_hits_T_32 = _sector_hits_T_31 | sectored_entries_0_5_valid_3; // @[package.scala 72:59]
  assign _sector_hits_T_33 = sectored_entries_0_5_tag ^ vpn; // @[TLB.scala 88:41]
  assign _sector_hits_T_35 = _sector_hits_T_33[26:2] == 25'h0; // @[TLB.scala 88:66]
  assign sector_hits_5 = _sector_hits_T_32 & _sector_hits_T_35; // @[TLB.scala 87:40]
  assign _sector_hits_T_36 = sectored_entries_0_6_valid_0 | sectored_entries_0_6_valid_1; // @[package.scala 72:59]
  assign _sector_hits_T_37 = _sector_hits_T_36 | sectored_entries_0_6_valid_2; // @[package.scala 72:59]
  assign _sector_hits_T_38 = _sector_hits_T_37 | sectored_entries_0_6_valid_3; // @[package.scala 72:59]
  assign _sector_hits_T_39 = sectored_entries_0_6_tag ^ vpn; // @[TLB.scala 88:41]
  assign _sector_hits_T_41 = _sector_hits_T_39[26:2] == 25'h0; // @[TLB.scala 88:66]
  assign sector_hits_6 = _sector_hits_T_38 & _sector_hits_T_41; // @[TLB.scala 87:40]
  assign _sector_hits_T_42 = sectored_entries_0_7_valid_0 | sectored_entries_0_7_valid_1; // @[package.scala 72:59]
  assign _sector_hits_T_43 = _sector_hits_T_42 | sectored_entries_0_7_valid_2; // @[package.scala 72:59]
  assign _sector_hits_T_44 = _sector_hits_T_43 | sectored_entries_0_7_valid_3; // @[package.scala 72:59]
  assign _sector_hits_T_45 = sectored_entries_0_7_tag ^ vpn; // @[TLB.scala 88:41]
  assign _sector_hits_T_47 = _sector_hits_T_45[26:2] == 25'h0; // @[TLB.scala 88:66]
  assign sector_hits_7 = _sector_hits_T_44 & _sector_hits_T_47; // @[TLB.scala 87:40]
  assign _superpage_hits_T_2 = superpage_entries_0_tag[26:18] == vpn[26:18]; // @[TLB.scala 95:77]
  assign _superpage_hits_T_4 = superpage_entries_0_valid_0 & _superpage_hits_T_2; // @[TLB.scala 95:29]
  assign superpage_hits_ignore_1 = superpage_entries_0_level < 2'h1; // @[TLB.scala 94:28]
  assign _superpage_hits_T_7 = superpage_entries_0_tag[17:9] == vpn[17:9]; // @[TLB.scala 95:77]
  assign _superpage_hits_T_8 = superpage_hits_ignore_1 | _superpage_hits_T_7; // @[TLB.scala 95:40]
  assign superpage_hits_0 = _superpage_hits_T_4 & _superpage_hits_T_8; // @[TLB.scala 95:29]
  assign _superpage_hits_T_16 = superpage_entries_1_tag[26:18] == vpn[26:18]; // @[TLB.scala 95:77]
  assign _superpage_hits_T_18 = superpage_entries_1_valid_0 & _superpage_hits_T_16; // @[TLB.scala 95:29]
  assign superpage_hits_ignore_4 = superpage_entries_1_level < 2'h1; // @[TLB.scala 94:28]
  assign _superpage_hits_T_21 = superpage_entries_1_tag[17:9] == vpn[17:9]; // @[TLB.scala 95:77]
  assign _superpage_hits_T_22 = superpage_hits_ignore_4 | _superpage_hits_T_21; // @[TLB.scala 95:40]
  assign superpage_hits_1 = _superpage_hits_T_18 & _superpage_hits_T_22; // @[TLB.scala 95:29]
  assign _superpage_hits_T_30 = superpage_entries_2_tag[26:18] == vpn[26:18]; // @[TLB.scala 95:77]
  assign _superpage_hits_T_32 = superpage_entries_2_valid_0 & _superpage_hits_T_30; // @[TLB.scala 95:29]
  assign superpage_hits_ignore_7 = superpage_entries_2_level < 2'h1; // @[TLB.scala 94:28]
  assign _superpage_hits_T_35 = superpage_entries_2_tag[17:9] == vpn[17:9]; // @[TLB.scala 95:77]
  assign _superpage_hits_T_36 = superpage_hits_ignore_7 | _superpage_hits_T_35; // @[TLB.scala 95:40]
  assign superpage_hits_2 = _superpage_hits_T_32 & _superpage_hits_T_36; // @[TLB.scala 95:29]
  assign _superpage_hits_T_44 = superpage_entries_3_tag[26:18] == vpn[26:18]; // @[TLB.scala 95:77]
  assign _superpage_hits_T_46 = superpage_entries_3_valid_0 & _superpage_hits_T_44; // @[TLB.scala 95:29]
  assign superpage_hits_ignore_10 = superpage_entries_3_level < 2'h1; // @[TLB.scala 94:28]
  assign _superpage_hits_T_49 = superpage_entries_3_tag[17:9] == vpn[17:9]; // @[TLB.scala 95:77]
  assign _superpage_hits_T_50 = superpage_hits_ignore_10 | _superpage_hits_T_49; // @[TLB.scala 95:40]
  assign superpage_hits_3 = _superpage_hits_T_46 & _superpage_hits_T_50; // @[TLB.scala 95:29]
  assign hitsVec_idx = vpn[1:0]; // @[package.scala 154:13]
  assign _GEN_1 = 2'h1 == hitsVec_idx ? sectored_entries_0_0_valid_1 : sectored_entries_0_0_valid_0; // @[TLB.scala 100:18]
  assign _GEN_2 = 2'h2 == hitsVec_idx ? sectored_entries_0_0_valid_2 : _GEN_1; // @[TLB.scala 100:18]
  assign _GEN_3 = 2'h3 == hitsVec_idx ? sectored_entries_0_0_valid_3 : _GEN_2; // @[TLB.scala 100:18]
  assign _hitsVec_T_3 = _GEN_3 & _sector_hits_T_5; // @[TLB.scala 100:18]
  assign hitsVec_0 = vm_enabled & _hitsVec_T_3; // @[TLB.scala 213:44]
  assign _GEN_5 = 2'h1 == hitsVec_idx ? sectored_entries_0_1_valid_1 : sectored_entries_0_1_valid_0; // @[TLB.scala 100:18]
  assign _GEN_6 = 2'h2 == hitsVec_idx ? sectored_entries_0_1_valid_2 : _GEN_5; // @[TLB.scala 100:18]
  assign _GEN_7 = 2'h3 == hitsVec_idx ? sectored_entries_0_1_valid_3 : _GEN_6; // @[TLB.scala 100:18]
  assign _hitsVec_T_7 = _GEN_7 & _sector_hits_T_11; // @[TLB.scala 100:18]
  assign hitsVec_1 = vm_enabled & _hitsVec_T_7; // @[TLB.scala 213:44]
  assign _GEN_9 = 2'h1 == hitsVec_idx ? sectored_entries_0_2_valid_1 : sectored_entries_0_2_valid_0; // @[TLB.scala 100:18]
  assign _GEN_10 = 2'h2 == hitsVec_idx ? sectored_entries_0_2_valid_2 : _GEN_9; // @[TLB.scala 100:18]
  assign _GEN_11 = 2'h3 == hitsVec_idx ? sectored_entries_0_2_valid_3 : _GEN_10; // @[TLB.scala 100:18]
  assign _hitsVec_T_11 = _GEN_11 & _sector_hits_T_17; // @[TLB.scala 100:18]
  assign hitsVec_2 = vm_enabled & _hitsVec_T_11; // @[TLB.scala 213:44]
  assign _GEN_13 = 2'h1 == hitsVec_idx ? sectored_entries_0_3_valid_1 : sectored_entries_0_3_valid_0; // @[TLB.scala 100:18]
  assign _GEN_14 = 2'h2 == hitsVec_idx ? sectored_entries_0_3_valid_2 : _GEN_13; // @[TLB.scala 100:18]
  assign _GEN_15 = 2'h3 == hitsVec_idx ? sectored_entries_0_3_valid_3 : _GEN_14; // @[TLB.scala 100:18]
  assign _hitsVec_T_15 = _GEN_15 & _sector_hits_T_23; // @[TLB.scala 100:18]
  assign hitsVec_3 = vm_enabled & _hitsVec_T_15; // @[TLB.scala 213:44]
  assign _GEN_17 = 2'h1 == hitsVec_idx ? sectored_entries_0_4_valid_1 : sectored_entries_0_4_valid_0; // @[TLB.scala 100:18]
  assign _GEN_18 = 2'h2 == hitsVec_idx ? sectored_entries_0_4_valid_2 : _GEN_17; // @[TLB.scala 100:18]
  assign _GEN_19 = 2'h3 == hitsVec_idx ? sectored_entries_0_4_valid_3 : _GEN_18; // @[TLB.scala 100:18]
  assign _hitsVec_T_19 = _GEN_19 & _sector_hits_T_29; // @[TLB.scala 100:18]
  assign hitsVec_4 = vm_enabled & _hitsVec_T_19; // @[TLB.scala 213:44]
  assign _GEN_21 = 2'h1 == hitsVec_idx ? sectored_entries_0_5_valid_1 : sectored_entries_0_5_valid_0; // @[TLB.scala 100:18]
  assign _GEN_22 = 2'h2 == hitsVec_idx ? sectored_entries_0_5_valid_2 : _GEN_21; // @[TLB.scala 100:18]
  assign _GEN_23 = 2'h3 == hitsVec_idx ? sectored_entries_0_5_valid_3 : _GEN_22; // @[TLB.scala 100:18]
  assign _hitsVec_T_23 = _GEN_23 & _sector_hits_T_35; // @[TLB.scala 100:18]
  assign hitsVec_5 = vm_enabled & _hitsVec_T_23; // @[TLB.scala 213:44]
  assign _GEN_25 = 2'h1 == hitsVec_idx ? sectored_entries_0_6_valid_1 : sectored_entries_0_6_valid_0; // @[TLB.scala 100:18]
  assign _GEN_26 = 2'h2 == hitsVec_idx ? sectored_entries_0_6_valid_2 : _GEN_25; // @[TLB.scala 100:18]
  assign _GEN_27 = 2'h3 == hitsVec_idx ? sectored_entries_0_6_valid_3 : _GEN_26; // @[TLB.scala 100:18]
  assign _hitsVec_T_27 = _GEN_27 & _sector_hits_T_41; // @[TLB.scala 100:18]
  assign hitsVec_6 = vm_enabled & _hitsVec_T_27; // @[TLB.scala 213:44]
  assign _GEN_29 = 2'h1 == hitsVec_idx ? sectored_entries_0_7_valid_1 : sectored_entries_0_7_valid_0; // @[TLB.scala 100:18]
  assign _GEN_30 = 2'h2 == hitsVec_idx ? sectored_entries_0_7_valid_2 : _GEN_29; // @[TLB.scala 100:18]
  assign _GEN_31 = 2'h3 == hitsVec_idx ? sectored_entries_0_7_valid_3 : _GEN_30; // @[TLB.scala 100:18]
  assign _hitsVec_T_31 = _GEN_31 & _sector_hits_T_47; // @[TLB.scala 100:18]
  assign hitsVec_7 = vm_enabled & _hitsVec_T_31; // @[TLB.scala 213:44]
  assign hitsVec_8 = vm_enabled & superpage_hits_0; // @[TLB.scala 213:44]
  assign hitsVec_9 = vm_enabled & superpage_hits_1; // @[TLB.scala 213:44]
  assign hitsVec_10 = vm_enabled & superpage_hits_2; // @[TLB.scala 213:44]
  assign hitsVec_11 = vm_enabled & superpage_hits_3; // @[TLB.scala 213:44]
  assign _hitsVec_T_94 = special_entry_tag[26:18] == vpn[26:18]; // @[TLB.scala 95:77]
  assign _hitsVec_T_96 = special_entry_valid_0 & _hitsVec_T_94; // @[TLB.scala 95:29]
  assign _hitsVec_T_99 = special_entry_tag[17:9] == vpn[17:9]; // @[TLB.scala 95:77]
  assign _hitsVec_T_100 = mpu_ppn_ignore | _hitsVec_T_99; // @[TLB.scala 95:40]
  assign _hitsVec_T_101 = _hitsVec_T_96 & _hitsVec_T_100; // @[TLB.scala 95:29]
  assign _hitsVec_T_104 = special_entry_tag[8:0] == vpn[8:0]; // @[TLB.scala 95:77]
  assign _hitsVec_T_105 = mpu_ppn_ignore_1 | _hitsVec_T_104; // @[TLB.scala 95:40]
  assign _hitsVec_T_106 = _hitsVec_T_101 & _hitsVec_T_105; // @[TLB.scala 95:29]
  assign hitsVec_12 = vm_enabled & _hitsVec_T_106; // @[TLB.scala 213:44]
  assign real_hits_lo = {hitsVec_5,hitsVec_4,hitsVec_3,hitsVec_2,hitsVec_1,hitsVec_0}; // @[Cat.scala 30:58]
  assign real_hits = {hitsVec_12,hitsVec_11,hitsVec_10,hitsVec_9,hitsVec_8,hitsVec_7,hitsVec_6,real_hits_lo}; // @[Cat.scala 30:58]
  assign hits_hi = ~vm_enabled; // @[TLB.scala 215:18]
  assign hits = {hits_hi,hitsVec_12,hitsVec_11,hitsVec_10,hitsVec_9,hitsVec_8,hitsVec_7,hitsVec_6,real_hits_lo}; // @[Cat.scala 30:58]
  assign newEntry_g = io_ptw_resp_bits_pte_g & io_ptw_resp_bits_pte_v; // @[TLB.scala 224:25]
  assign _newEntry_sr_T_1 = io_ptw_resp_bits_pte_x & ~io_ptw_resp_bits_pte_w; // @[PTW.scala 73:44]
  assign _newEntry_sr_T_2 = io_ptw_resp_bits_pte_r | _newEntry_sr_T_1; // @[PTW.scala 73:38]
  assign _newEntry_sr_T_3 = io_ptw_resp_bits_pte_v & _newEntry_sr_T_2; // @[PTW.scala 73:32]
  assign _newEntry_sr_T_4 = _newEntry_sr_T_3 & io_ptw_resp_bits_pte_a; // @[PTW.scala 73:52]
  assign newEntry_sr = _newEntry_sr_T_4 & io_ptw_resp_bits_pte_r; // @[PTW.scala 77:35]
  assign _newEntry_sw_T_5 = _newEntry_sr_T_4 & io_ptw_resp_bits_pte_w; // @[PTW.scala 78:35]
  assign newEntry_sw = _newEntry_sw_T_5 & io_ptw_resp_bits_pte_d; // @[PTW.scala 78:40]
  assign newEntry_sx = _newEntry_sr_T_4 & io_ptw_resp_bits_pte_x; // @[PTW.scala 79:35]
  assign special_entry_data_0_lo = {prot_x,prot_r,_prot_w_T_31,prot_al,prot_al,prot_eff,cacheable,1'h0}; // @[TLB.scala 122:24]
  assign _special_entry_data_0_T = {refill_ppn,io_ptw_resp_bits_pte_u,newEntry_g,io_ptw_resp_bits_ae,newEntry_sw,newEntry_sx,newEntry_sr,prot_w,special_entry_data_0_lo}; // @[TLB.scala 122:24]
  assign _GEN_32 = invalidate_refill ? 1'h0 : 1'h1; // @[TLB.scala 241:34]
  assign _T_2 = io_ptw_resp_bits_level < 2'h2; // @[TLB.scala 243:40]
  assign _T_3 = r_superpage_repl_addr == 2'h0; // @[TLB.scala 244:82]
  assign _GEN_35 = _T_3 ? _GEN_32 : superpage_entries_0_valid_0; // @[TLB.scala 244:89]
  assign _T_4 = r_superpage_repl_addr == 2'h1; // @[TLB.scala 244:82]
  assign _GEN_39 = _T_4 ? _GEN_32 : superpage_entries_1_valid_0; // @[TLB.scala 244:89]
  assign _T_5 = r_superpage_repl_addr == 2'h2; // @[TLB.scala 244:82]
  assign _GEN_43 = _T_5 ? _GEN_32 : superpage_entries_2_valid_0; // @[TLB.scala 244:89]
  assign _T_6 = r_superpage_repl_addr == 2'h3; // @[TLB.scala 244:82]
  assign _GEN_47 = _T_6 ? _GEN_32 : superpage_entries_3_valid_0; // @[TLB.scala 244:89]
  assign waddr = r_sectored_hit ? r_sectored_hit_addr : r_sectored_repl_addr; // @[TLB.scala 250:22]
  assign _T_7 = waddr == 3'h0; // @[TLB.scala 251:75]
  assign _GEN_49 = r_sectored_hit ? sectored_entries_0_0_valid_0 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_50 = r_sectored_hit ? sectored_entries_0_0_valid_1 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_51 = r_sectored_hit ? sectored_entries_0_0_valid_2 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_52 = r_sectored_hit ? sectored_entries_0_0_valid_3 : 1'h0; // @[TLB.scala 252:32]
  assign idx = r_refill_tag[1:0]; // @[package.scala 154:13]
  assign _GEN_921 = 2'h0 == idx; // @[TLB.scala 121:16]
  assign _GEN_53 = _GEN_921 | _GEN_49; // @[TLB.scala 121:16]
  assign _GEN_922 = 2'h1 == idx; // @[TLB.scala 121:16]
  assign _GEN_54 = _GEN_922 | _GEN_50; // @[TLB.scala 121:16]
  assign _GEN_923 = 2'h2 == idx; // @[TLB.scala 121:16]
  assign _GEN_55 = _GEN_923 | _GEN_51; // @[TLB.scala 121:16]
  assign _GEN_924 = 2'h3 == idx; // @[TLB.scala 121:16]
  assign _GEN_56 = _GEN_924 | _GEN_52; // @[TLB.scala 121:16]
  assign _GEN_61 = invalidate_refill ? 1'h0 : _GEN_53; // @[TLB.scala 254:34]
  assign _GEN_62 = invalidate_refill ? 1'h0 : _GEN_54; // @[TLB.scala 254:34]
  assign _GEN_63 = invalidate_refill ? 1'h0 : _GEN_55; // @[TLB.scala 254:34]
  assign _GEN_64 = invalidate_refill ? 1'h0 : _GEN_56; // @[TLB.scala 254:34]
  assign _GEN_65 = _T_7 ? _GEN_61 : sectored_entries_0_0_valid_0; // @[TLB.scala 251:82]
  assign _GEN_66 = _T_7 ? _GEN_62 : sectored_entries_0_0_valid_1; // @[TLB.scala 251:82]
  assign _GEN_67 = _T_7 ? _GEN_63 : sectored_entries_0_0_valid_2; // @[TLB.scala 251:82]
  assign _GEN_68 = _T_7 ? _GEN_64 : sectored_entries_0_0_valid_3; // @[TLB.scala 251:82]
  assign _T_9 = waddr == 3'h1; // @[TLB.scala 251:75]
  assign _GEN_75 = r_sectored_hit ? sectored_entries_0_1_valid_0 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_76 = r_sectored_hit ? sectored_entries_0_1_valid_1 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_77 = r_sectored_hit ? sectored_entries_0_1_valid_2 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_78 = r_sectored_hit ? sectored_entries_0_1_valid_3 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_79 = _GEN_921 | _GEN_75; // @[TLB.scala 121:16]
  assign _GEN_80 = _GEN_922 | _GEN_76; // @[TLB.scala 121:16]
  assign _GEN_81 = _GEN_923 | _GEN_77; // @[TLB.scala 121:16]
  assign _GEN_82 = _GEN_924 | _GEN_78; // @[TLB.scala 121:16]
  assign _GEN_87 = invalidate_refill ? 1'h0 : _GEN_79; // @[TLB.scala 254:34]
  assign _GEN_88 = invalidate_refill ? 1'h0 : _GEN_80; // @[TLB.scala 254:34]
  assign _GEN_89 = invalidate_refill ? 1'h0 : _GEN_81; // @[TLB.scala 254:34]
  assign _GEN_90 = invalidate_refill ? 1'h0 : _GEN_82; // @[TLB.scala 254:34]
  assign _GEN_91 = _T_9 ? _GEN_87 : sectored_entries_0_1_valid_0; // @[TLB.scala 251:82]
  assign _GEN_92 = _T_9 ? _GEN_88 : sectored_entries_0_1_valid_1; // @[TLB.scala 251:82]
  assign _GEN_93 = _T_9 ? _GEN_89 : sectored_entries_0_1_valid_2; // @[TLB.scala 251:82]
  assign _GEN_94 = _T_9 ? _GEN_90 : sectored_entries_0_1_valid_3; // @[TLB.scala 251:82]
  assign _T_11 = waddr == 3'h2; // @[TLB.scala 251:75]
  assign _GEN_101 = r_sectored_hit ? sectored_entries_0_2_valid_0 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_102 = r_sectored_hit ? sectored_entries_0_2_valid_1 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_103 = r_sectored_hit ? sectored_entries_0_2_valid_2 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_104 = r_sectored_hit ? sectored_entries_0_2_valid_3 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_105 = _GEN_921 | _GEN_101; // @[TLB.scala 121:16]
  assign _GEN_106 = _GEN_922 | _GEN_102; // @[TLB.scala 121:16]
  assign _GEN_107 = _GEN_923 | _GEN_103; // @[TLB.scala 121:16]
  assign _GEN_108 = _GEN_924 | _GEN_104; // @[TLB.scala 121:16]
  assign _GEN_113 = invalidate_refill ? 1'h0 : _GEN_105; // @[TLB.scala 254:34]
  assign _GEN_114 = invalidate_refill ? 1'h0 : _GEN_106; // @[TLB.scala 254:34]
  assign _GEN_115 = invalidate_refill ? 1'h0 : _GEN_107; // @[TLB.scala 254:34]
  assign _GEN_116 = invalidate_refill ? 1'h0 : _GEN_108; // @[TLB.scala 254:34]
  assign _GEN_117 = _T_11 ? _GEN_113 : sectored_entries_0_2_valid_0; // @[TLB.scala 251:82]
  assign _GEN_118 = _T_11 ? _GEN_114 : sectored_entries_0_2_valid_1; // @[TLB.scala 251:82]
  assign _GEN_119 = _T_11 ? _GEN_115 : sectored_entries_0_2_valid_2; // @[TLB.scala 251:82]
  assign _GEN_120 = _T_11 ? _GEN_116 : sectored_entries_0_2_valid_3; // @[TLB.scala 251:82]
  assign _T_13 = waddr == 3'h3; // @[TLB.scala 251:75]
  assign _GEN_127 = r_sectored_hit ? sectored_entries_0_3_valid_0 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_128 = r_sectored_hit ? sectored_entries_0_3_valid_1 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_129 = r_sectored_hit ? sectored_entries_0_3_valid_2 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_130 = r_sectored_hit ? sectored_entries_0_3_valid_3 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_131 = _GEN_921 | _GEN_127; // @[TLB.scala 121:16]
  assign _GEN_132 = _GEN_922 | _GEN_128; // @[TLB.scala 121:16]
  assign _GEN_133 = _GEN_923 | _GEN_129; // @[TLB.scala 121:16]
  assign _GEN_134 = _GEN_924 | _GEN_130; // @[TLB.scala 121:16]
  assign _GEN_139 = invalidate_refill ? 1'h0 : _GEN_131; // @[TLB.scala 254:34]
  assign _GEN_140 = invalidate_refill ? 1'h0 : _GEN_132; // @[TLB.scala 254:34]
  assign _GEN_141 = invalidate_refill ? 1'h0 : _GEN_133; // @[TLB.scala 254:34]
  assign _GEN_142 = invalidate_refill ? 1'h0 : _GEN_134; // @[TLB.scala 254:34]
  assign _GEN_143 = _T_13 ? _GEN_139 : sectored_entries_0_3_valid_0; // @[TLB.scala 251:82]
  assign _GEN_144 = _T_13 ? _GEN_140 : sectored_entries_0_3_valid_1; // @[TLB.scala 251:82]
  assign _GEN_145 = _T_13 ? _GEN_141 : sectored_entries_0_3_valid_2; // @[TLB.scala 251:82]
  assign _GEN_146 = _T_13 ? _GEN_142 : sectored_entries_0_3_valid_3; // @[TLB.scala 251:82]
  assign _T_15 = waddr == 3'h4; // @[TLB.scala 251:75]
  assign _GEN_153 = r_sectored_hit ? sectored_entries_0_4_valid_0 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_154 = r_sectored_hit ? sectored_entries_0_4_valid_1 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_155 = r_sectored_hit ? sectored_entries_0_4_valid_2 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_156 = r_sectored_hit ? sectored_entries_0_4_valid_3 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_157 = _GEN_921 | _GEN_153; // @[TLB.scala 121:16]
  assign _GEN_158 = _GEN_922 | _GEN_154; // @[TLB.scala 121:16]
  assign _GEN_159 = _GEN_923 | _GEN_155; // @[TLB.scala 121:16]
  assign _GEN_160 = _GEN_924 | _GEN_156; // @[TLB.scala 121:16]
  assign _GEN_165 = invalidate_refill ? 1'h0 : _GEN_157; // @[TLB.scala 254:34]
  assign _GEN_166 = invalidate_refill ? 1'h0 : _GEN_158; // @[TLB.scala 254:34]
  assign _GEN_167 = invalidate_refill ? 1'h0 : _GEN_159; // @[TLB.scala 254:34]
  assign _GEN_168 = invalidate_refill ? 1'h0 : _GEN_160; // @[TLB.scala 254:34]
  assign _GEN_169 = _T_15 ? _GEN_165 : sectored_entries_0_4_valid_0; // @[TLB.scala 251:82]
  assign _GEN_170 = _T_15 ? _GEN_166 : sectored_entries_0_4_valid_1; // @[TLB.scala 251:82]
  assign _GEN_171 = _T_15 ? _GEN_167 : sectored_entries_0_4_valid_2; // @[TLB.scala 251:82]
  assign _GEN_172 = _T_15 ? _GEN_168 : sectored_entries_0_4_valid_3; // @[TLB.scala 251:82]
  assign _T_17 = waddr == 3'h5; // @[TLB.scala 251:75]
  assign _GEN_179 = r_sectored_hit ? sectored_entries_0_5_valid_0 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_180 = r_sectored_hit ? sectored_entries_0_5_valid_1 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_181 = r_sectored_hit ? sectored_entries_0_5_valid_2 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_182 = r_sectored_hit ? sectored_entries_0_5_valid_3 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_183 = _GEN_921 | _GEN_179; // @[TLB.scala 121:16]
  assign _GEN_184 = _GEN_922 | _GEN_180; // @[TLB.scala 121:16]
  assign _GEN_185 = _GEN_923 | _GEN_181; // @[TLB.scala 121:16]
  assign _GEN_186 = _GEN_924 | _GEN_182; // @[TLB.scala 121:16]
  assign _GEN_191 = invalidate_refill ? 1'h0 : _GEN_183; // @[TLB.scala 254:34]
  assign _GEN_192 = invalidate_refill ? 1'h0 : _GEN_184; // @[TLB.scala 254:34]
  assign _GEN_193 = invalidate_refill ? 1'h0 : _GEN_185; // @[TLB.scala 254:34]
  assign _GEN_194 = invalidate_refill ? 1'h0 : _GEN_186; // @[TLB.scala 254:34]
  assign _GEN_195 = _T_17 ? _GEN_191 : sectored_entries_0_5_valid_0; // @[TLB.scala 251:82]
  assign _GEN_196 = _T_17 ? _GEN_192 : sectored_entries_0_5_valid_1; // @[TLB.scala 251:82]
  assign _GEN_197 = _T_17 ? _GEN_193 : sectored_entries_0_5_valid_2; // @[TLB.scala 251:82]
  assign _GEN_198 = _T_17 ? _GEN_194 : sectored_entries_0_5_valid_3; // @[TLB.scala 251:82]
  assign _T_19 = waddr == 3'h6; // @[TLB.scala 251:75]
  assign _GEN_205 = r_sectored_hit ? sectored_entries_0_6_valid_0 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_206 = r_sectored_hit ? sectored_entries_0_6_valid_1 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_207 = r_sectored_hit ? sectored_entries_0_6_valid_2 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_208 = r_sectored_hit ? sectored_entries_0_6_valid_3 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_209 = _GEN_921 | _GEN_205; // @[TLB.scala 121:16]
  assign _GEN_210 = _GEN_922 | _GEN_206; // @[TLB.scala 121:16]
  assign _GEN_211 = _GEN_923 | _GEN_207; // @[TLB.scala 121:16]
  assign _GEN_212 = _GEN_924 | _GEN_208; // @[TLB.scala 121:16]
  assign _GEN_217 = invalidate_refill ? 1'h0 : _GEN_209; // @[TLB.scala 254:34]
  assign _GEN_218 = invalidate_refill ? 1'h0 : _GEN_210; // @[TLB.scala 254:34]
  assign _GEN_219 = invalidate_refill ? 1'h0 : _GEN_211; // @[TLB.scala 254:34]
  assign _GEN_220 = invalidate_refill ? 1'h0 : _GEN_212; // @[TLB.scala 254:34]
  assign _GEN_221 = _T_19 ? _GEN_217 : sectored_entries_0_6_valid_0; // @[TLB.scala 251:82]
  assign _GEN_222 = _T_19 ? _GEN_218 : sectored_entries_0_6_valid_1; // @[TLB.scala 251:82]
  assign _GEN_223 = _T_19 ? _GEN_219 : sectored_entries_0_6_valid_2; // @[TLB.scala 251:82]
  assign _GEN_224 = _T_19 ? _GEN_220 : sectored_entries_0_6_valid_3; // @[TLB.scala 251:82]
  assign _T_21 = waddr == 3'h7; // @[TLB.scala 251:75]
  assign _GEN_231 = r_sectored_hit ? sectored_entries_0_7_valid_0 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_232 = r_sectored_hit ? sectored_entries_0_7_valid_1 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_233 = r_sectored_hit ? sectored_entries_0_7_valid_2 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_234 = r_sectored_hit ? sectored_entries_0_7_valid_3 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_235 = _GEN_921 | _GEN_231; // @[TLB.scala 121:16]
  assign _GEN_236 = _GEN_922 | _GEN_232; // @[TLB.scala 121:16]
  assign _GEN_237 = _GEN_923 | _GEN_233; // @[TLB.scala 121:16]
  assign _GEN_238 = _GEN_924 | _GEN_234; // @[TLB.scala 121:16]
  assign _GEN_243 = invalidate_refill ? 1'h0 : _GEN_235; // @[TLB.scala 254:34]
  assign _GEN_244 = invalidate_refill ? 1'h0 : _GEN_236; // @[TLB.scala 254:34]
  assign _GEN_245 = invalidate_refill ? 1'h0 : _GEN_237; // @[TLB.scala 254:34]
  assign _GEN_246 = invalidate_refill ? 1'h0 : _GEN_238; // @[TLB.scala 254:34]
  assign _GEN_247 = _T_21 ? _GEN_243 : sectored_entries_0_7_valid_0; // @[TLB.scala 251:82]
  assign _GEN_248 = _T_21 ? _GEN_244 : sectored_entries_0_7_valid_1; // @[TLB.scala 251:82]
  assign _GEN_249 = _T_21 ? _GEN_245 : sectored_entries_0_7_valid_2; // @[TLB.scala 251:82]
  assign _GEN_250 = _T_21 ? _GEN_246 : sectored_entries_0_7_valid_3; // @[TLB.scala 251:82]
  assign _GEN_259 = _T_2 ? _GEN_35 : superpage_entries_0_valid_0; // @[TLB.scala 243:54]
  assign _GEN_263 = _T_2 ? _GEN_39 : superpage_entries_1_valid_0; // @[TLB.scala 243:54]
  assign _GEN_267 = _T_2 ? _GEN_43 : superpage_entries_2_valid_0; // @[TLB.scala 243:54]
  assign _GEN_271 = _T_2 ? _GEN_47 : superpage_entries_3_valid_0; // @[TLB.scala 243:54]
  assign _GEN_273 = _T_2 ? sectored_entries_0_0_valid_0 : _GEN_65; // @[TLB.scala 243:54]
  assign _GEN_274 = _T_2 ? sectored_entries_0_0_valid_1 : _GEN_66; // @[TLB.scala 243:54]
  assign _GEN_275 = _T_2 ? sectored_entries_0_0_valid_2 : _GEN_67; // @[TLB.scala 243:54]
  assign _GEN_276 = _T_2 ? sectored_entries_0_0_valid_3 : _GEN_68; // @[TLB.scala 243:54]
  assign _GEN_283 = _T_2 ? sectored_entries_0_1_valid_0 : _GEN_91; // @[TLB.scala 243:54]
  assign _GEN_284 = _T_2 ? sectored_entries_0_1_valid_1 : _GEN_92; // @[TLB.scala 243:54]
  assign _GEN_285 = _T_2 ? sectored_entries_0_1_valid_2 : _GEN_93; // @[TLB.scala 243:54]
  assign _GEN_286 = _T_2 ? sectored_entries_0_1_valid_3 : _GEN_94; // @[TLB.scala 243:54]
  assign _GEN_293 = _T_2 ? sectored_entries_0_2_valid_0 : _GEN_117; // @[TLB.scala 243:54]
  assign _GEN_294 = _T_2 ? sectored_entries_0_2_valid_1 : _GEN_118; // @[TLB.scala 243:54]
  assign _GEN_295 = _T_2 ? sectored_entries_0_2_valid_2 : _GEN_119; // @[TLB.scala 243:54]
  assign _GEN_296 = _T_2 ? sectored_entries_0_2_valid_3 : _GEN_120; // @[TLB.scala 243:54]
  assign _GEN_303 = _T_2 ? sectored_entries_0_3_valid_0 : _GEN_143; // @[TLB.scala 243:54]
  assign _GEN_304 = _T_2 ? sectored_entries_0_3_valid_1 : _GEN_144; // @[TLB.scala 243:54]
  assign _GEN_305 = _T_2 ? sectored_entries_0_3_valid_2 : _GEN_145; // @[TLB.scala 243:54]
  assign _GEN_306 = _T_2 ? sectored_entries_0_3_valid_3 : _GEN_146; // @[TLB.scala 243:54]
  assign _GEN_313 = _T_2 ? sectored_entries_0_4_valid_0 : _GEN_169; // @[TLB.scala 243:54]
  assign _GEN_314 = _T_2 ? sectored_entries_0_4_valid_1 : _GEN_170; // @[TLB.scala 243:54]
  assign _GEN_315 = _T_2 ? sectored_entries_0_4_valid_2 : _GEN_171; // @[TLB.scala 243:54]
  assign _GEN_316 = _T_2 ? sectored_entries_0_4_valid_3 : _GEN_172; // @[TLB.scala 243:54]
  assign _GEN_323 = _T_2 ? sectored_entries_0_5_valid_0 : _GEN_195; // @[TLB.scala 243:54]
  assign _GEN_324 = _T_2 ? sectored_entries_0_5_valid_1 : _GEN_196; // @[TLB.scala 243:54]
  assign _GEN_325 = _T_2 ? sectored_entries_0_5_valid_2 : _GEN_197; // @[TLB.scala 243:54]
  assign _GEN_326 = _T_2 ? sectored_entries_0_5_valid_3 : _GEN_198; // @[TLB.scala 243:54]
  assign _GEN_333 = _T_2 ? sectored_entries_0_6_valid_0 : _GEN_221; // @[TLB.scala 243:54]
  assign _GEN_334 = _T_2 ? sectored_entries_0_6_valid_1 : _GEN_222; // @[TLB.scala 243:54]
  assign _GEN_335 = _T_2 ? sectored_entries_0_6_valid_2 : _GEN_223; // @[TLB.scala 243:54]
  assign _GEN_336 = _T_2 ? sectored_entries_0_6_valid_3 : _GEN_224; // @[TLB.scala 243:54]
  assign _GEN_343 = _T_2 ? sectored_entries_0_7_valid_0 : _GEN_247; // @[TLB.scala 243:54]
  assign _GEN_344 = _T_2 ? sectored_entries_0_7_valid_1 : _GEN_248; // @[TLB.scala 243:54]
  assign _GEN_345 = _T_2 ? sectored_entries_0_7_valid_2 : _GEN_249; // @[TLB.scala 243:54]
  assign _GEN_346 = _T_2 ? sectored_entries_0_7_valid_3 : _GEN_250; // @[TLB.scala 243:54]
  assign _GEN_355 = io_ptw_resp_bits_homogeneous ? special_entry_valid_0 : _GEN_32; // @[TLB.scala 238:68]
  assign _GEN_359 = io_ptw_resp_bits_homogeneous ? _GEN_259 : superpage_entries_0_valid_0; // @[TLB.scala 238:68]
  assign _GEN_363 = io_ptw_resp_bits_homogeneous ? _GEN_263 : superpage_entries_1_valid_0; // @[TLB.scala 238:68]
  assign _GEN_367 = io_ptw_resp_bits_homogeneous ? _GEN_267 : superpage_entries_2_valid_0; // @[TLB.scala 238:68]
  assign _GEN_371 = io_ptw_resp_bits_homogeneous ? _GEN_271 : superpage_entries_3_valid_0; // @[TLB.scala 238:68]
  assign _GEN_373 = io_ptw_resp_bits_homogeneous ? _GEN_273 : sectored_entries_0_0_valid_0; // @[TLB.scala 238:68]
  assign _GEN_374 = io_ptw_resp_bits_homogeneous ? _GEN_274 : sectored_entries_0_0_valid_1; // @[TLB.scala 238:68]
  assign _GEN_375 = io_ptw_resp_bits_homogeneous ? _GEN_275 : sectored_entries_0_0_valid_2; // @[TLB.scala 238:68]
  assign _GEN_376 = io_ptw_resp_bits_homogeneous ? _GEN_276 : sectored_entries_0_0_valid_3; // @[TLB.scala 238:68]
  assign _GEN_383 = io_ptw_resp_bits_homogeneous ? _GEN_283 : sectored_entries_0_1_valid_0; // @[TLB.scala 238:68]
  assign _GEN_384 = io_ptw_resp_bits_homogeneous ? _GEN_284 : sectored_entries_0_1_valid_1; // @[TLB.scala 238:68]
  assign _GEN_385 = io_ptw_resp_bits_homogeneous ? _GEN_285 : sectored_entries_0_1_valid_2; // @[TLB.scala 238:68]
  assign _GEN_386 = io_ptw_resp_bits_homogeneous ? _GEN_286 : sectored_entries_0_1_valid_3; // @[TLB.scala 238:68]
  assign _GEN_393 = io_ptw_resp_bits_homogeneous ? _GEN_293 : sectored_entries_0_2_valid_0; // @[TLB.scala 238:68]
  assign _GEN_394 = io_ptw_resp_bits_homogeneous ? _GEN_294 : sectored_entries_0_2_valid_1; // @[TLB.scala 238:68]
  assign _GEN_395 = io_ptw_resp_bits_homogeneous ? _GEN_295 : sectored_entries_0_2_valid_2; // @[TLB.scala 238:68]
  assign _GEN_396 = io_ptw_resp_bits_homogeneous ? _GEN_296 : sectored_entries_0_2_valid_3; // @[TLB.scala 238:68]
  assign _GEN_403 = io_ptw_resp_bits_homogeneous ? _GEN_303 : sectored_entries_0_3_valid_0; // @[TLB.scala 238:68]
  assign _GEN_404 = io_ptw_resp_bits_homogeneous ? _GEN_304 : sectored_entries_0_3_valid_1; // @[TLB.scala 238:68]
  assign _GEN_405 = io_ptw_resp_bits_homogeneous ? _GEN_305 : sectored_entries_0_3_valid_2; // @[TLB.scala 238:68]
  assign _GEN_406 = io_ptw_resp_bits_homogeneous ? _GEN_306 : sectored_entries_0_3_valid_3; // @[TLB.scala 238:68]
  assign _GEN_413 = io_ptw_resp_bits_homogeneous ? _GEN_313 : sectored_entries_0_4_valid_0; // @[TLB.scala 238:68]
  assign _GEN_414 = io_ptw_resp_bits_homogeneous ? _GEN_314 : sectored_entries_0_4_valid_1; // @[TLB.scala 238:68]
  assign _GEN_415 = io_ptw_resp_bits_homogeneous ? _GEN_315 : sectored_entries_0_4_valid_2; // @[TLB.scala 238:68]
  assign _GEN_416 = io_ptw_resp_bits_homogeneous ? _GEN_316 : sectored_entries_0_4_valid_3; // @[TLB.scala 238:68]
  assign _GEN_423 = io_ptw_resp_bits_homogeneous ? _GEN_323 : sectored_entries_0_5_valid_0; // @[TLB.scala 238:68]
  assign _GEN_424 = io_ptw_resp_bits_homogeneous ? _GEN_324 : sectored_entries_0_5_valid_1; // @[TLB.scala 238:68]
  assign _GEN_425 = io_ptw_resp_bits_homogeneous ? _GEN_325 : sectored_entries_0_5_valid_2; // @[TLB.scala 238:68]
  assign _GEN_426 = io_ptw_resp_bits_homogeneous ? _GEN_326 : sectored_entries_0_5_valid_3; // @[TLB.scala 238:68]
  assign _GEN_433 = io_ptw_resp_bits_homogeneous ? _GEN_333 : sectored_entries_0_6_valid_0; // @[TLB.scala 238:68]
  assign _GEN_434 = io_ptw_resp_bits_homogeneous ? _GEN_334 : sectored_entries_0_6_valid_1; // @[TLB.scala 238:68]
  assign _GEN_435 = io_ptw_resp_bits_homogeneous ? _GEN_335 : sectored_entries_0_6_valid_2; // @[TLB.scala 238:68]
  assign _GEN_436 = io_ptw_resp_bits_homogeneous ? _GEN_336 : sectored_entries_0_6_valid_3; // @[TLB.scala 238:68]
  assign _GEN_443 = io_ptw_resp_bits_homogeneous ? _GEN_343 : sectored_entries_0_7_valid_0; // @[TLB.scala 238:68]
  assign _GEN_444 = io_ptw_resp_bits_homogeneous ? _GEN_344 : sectored_entries_0_7_valid_1; // @[TLB.scala 238:68]
  assign _GEN_445 = io_ptw_resp_bits_homogeneous ? _GEN_345 : sectored_entries_0_7_valid_2; // @[TLB.scala 238:68]
  assign _GEN_446 = io_ptw_resp_bits_homogeneous ? _GEN_346 : sectored_entries_0_7_valid_3; // @[TLB.scala 238:68]
  assign _GEN_455 = io_ptw_resp_valid ? _GEN_355 : special_entry_valid_0; // @[TLB.scala 218:20]
  assign _GEN_459 = io_ptw_resp_valid ? _GEN_359 : superpage_entries_0_valid_0; // @[TLB.scala 218:20]
  assign _GEN_463 = io_ptw_resp_valid ? _GEN_363 : superpage_entries_1_valid_0; // @[TLB.scala 218:20]
  assign _GEN_467 = io_ptw_resp_valid ? _GEN_367 : superpage_entries_2_valid_0; // @[TLB.scala 218:20]
  assign _GEN_471 = io_ptw_resp_valid ? _GEN_371 : superpage_entries_3_valid_0; // @[TLB.scala 218:20]
  assign _GEN_473 = io_ptw_resp_valid ? _GEN_373 : sectored_entries_0_0_valid_0; // @[TLB.scala 218:20]
  assign _GEN_474 = io_ptw_resp_valid ? _GEN_374 : sectored_entries_0_0_valid_1; // @[TLB.scala 218:20]
  assign _GEN_475 = io_ptw_resp_valid ? _GEN_375 : sectored_entries_0_0_valid_2; // @[TLB.scala 218:20]
  assign _GEN_476 = io_ptw_resp_valid ? _GEN_376 : sectored_entries_0_0_valid_3; // @[TLB.scala 218:20]
  assign _GEN_483 = io_ptw_resp_valid ? _GEN_383 : sectored_entries_0_1_valid_0; // @[TLB.scala 218:20]
  assign _GEN_484 = io_ptw_resp_valid ? _GEN_384 : sectored_entries_0_1_valid_1; // @[TLB.scala 218:20]
  assign _GEN_485 = io_ptw_resp_valid ? _GEN_385 : sectored_entries_0_1_valid_2; // @[TLB.scala 218:20]
  assign _GEN_486 = io_ptw_resp_valid ? _GEN_386 : sectored_entries_0_1_valid_3; // @[TLB.scala 218:20]
  assign _GEN_493 = io_ptw_resp_valid ? _GEN_393 : sectored_entries_0_2_valid_0; // @[TLB.scala 218:20]
  assign _GEN_494 = io_ptw_resp_valid ? _GEN_394 : sectored_entries_0_2_valid_1; // @[TLB.scala 218:20]
  assign _GEN_495 = io_ptw_resp_valid ? _GEN_395 : sectored_entries_0_2_valid_2; // @[TLB.scala 218:20]
  assign _GEN_496 = io_ptw_resp_valid ? _GEN_396 : sectored_entries_0_2_valid_3; // @[TLB.scala 218:20]
  assign _GEN_503 = io_ptw_resp_valid ? _GEN_403 : sectored_entries_0_3_valid_0; // @[TLB.scala 218:20]
  assign _GEN_504 = io_ptw_resp_valid ? _GEN_404 : sectored_entries_0_3_valid_1; // @[TLB.scala 218:20]
  assign _GEN_505 = io_ptw_resp_valid ? _GEN_405 : sectored_entries_0_3_valid_2; // @[TLB.scala 218:20]
  assign _GEN_506 = io_ptw_resp_valid ? _GEN_406 : sectored_entries_0_3_valid_3; // @[TLB.scala 218:20]
  assign _GEN_513 = io_ptw_resp_valid ? _GEN_413 : sectored_entries_0_4_valid_0; // @[TLB.scala 218:20]
  assign _GEN_514 = io_ptw_resp_valid ? _GEN_414 : sectored_entries_0_4_valid_1; // @[TLB.scala 218:20]
  assign _GEN_515 = io_ptw_resp_valid ? _GEN_415 : sectored_entries_0_4_valid_2; // @[TLB.scala 218:20]
  assign _GEN_516 = io_ptw_resp_valid ? _GEN_416 : sectored_entries_0_4_valid_3; // @[TLB.scala 218:20]
  assign _GEN_523 = io_ptw_resp_valid ? _GEN_423 : sectored_entries_0_5_valid_0; // @[TLB.scala 218:20]
  assign _GEN_524 = io_ptw_resp_valid ? _GEN_424 : sectored_entries_0_5_valid_1; // @[TLB.scala 218:20]
  assign _GEN_525 = io_ptw_resp_valid ? _GEN_425 : sectored_entries_0_5_valid_2; // @[TLB.scala 218:20]
  assign _GEN_526 = io_ptw_resp_valid ? _GEN_426 : sectored_entries_0_5_valid_3; // @[TLB.scala 218:20]
  assign _GEN_533 = io_ptw_resp_valid ? _GEN_433 : sectored_entries_0_6_valid_0; // @[TLB.scala 218:20]
  assign _GEN_534 = io_ptw_resp_valid ? _GEN_434 : sectored_entries_0_6_valid_1; // @[TLB.scala 218:20]
  assign _GEN_535 = io_ptw_resp_valid ? _GEN_435 : sectored_entries_0_6_valid_2; // @[TLB.scala 218:20]
  assign _GEN_536 = io_ptw_resp_valid ? _GEN_436 : sectored_entries_0_6_valid_3; // @[TLB.scala 218:20]
  assign _GEN_543 = io_ptw_resp_valid ? _GEN_443 : sectored_entries_0_7_valid_0; // @[TLB.scala 218:20]
  assign _GEN_544 = io_ptw_resp_valid ? _GEN_444 : sectored_entries_0_7_valid_1; // @[TLB.scala 218:20]
  assign _GEN_545 = io_ptw_resp_valid ? _GEN_445 : sectored_entries_0_7_valid_2; // @[TLB.scala 218:20]
  assign _GEN_546 = io_ptw_resp_valid ? _GEN_446 : sectored_entries_0_7_valid_3; // @[TLB.scala 218:20]
  assign _GEN_554 = 2'h1 == hitsVec_idx ? sectored_entries_0_0_data_1 : sectored_entries_0_0_data_0;
  assign _GEN_555 = 2'h2 == hitsVec_idx ? sectored_entries_0_0_data_2 : _GEN_554;
  assign _GEN_556 = 2'h3 == hitsVec_idx ? sectored_entries_0_0_data_3 : _GEN_555;
  assign _GEN_558 = 2'h1 == hitsVec_idx ? sectored_entries_0_1_data_1 : sectored_entries_0_1_data_0;
  assign _GEN_559 = 2'h2 == hitsVec_idx ? sectored_entries_0_1_data_2 : _GEN_558;
  assign _GEN_560 = 2'h3 == hitsVec_idx ? sectored_entries_0_1_data_3 : _GEN_559;
  assign _GEN_562 = 2'h1 == hitsVec_idx ? sectored_entries_0_2_data_1 : sectored_entries_0_2_data_0;
  assign _GEN_563 = 2'h2 == hitsVec_idx ? sectored_entries_0_2_data_2 : _GEN_562;
  assign _GEN_564 = 2'h3 == hitsVec_idx ? sectored_entries_0_2_data_3 : _GEN_563;
  assign _GEN_566 = 2'h1 == hitsVec_idx ? sectored_entries_0_3_data_1 : sectored_entries_0_3_data_0;
  assign _GEN_567 = 2'h2 == hitsVec_idx ? sectored_entries_0_3_data_2 : _GEN_566;
  assign _GEN_568 = 2'h3 == hitsVec_idx ? sectored_entries_0_3_data_3 : _GEN_567;
  assign _GEN_570 = 2'h1 == hitsVec_idx ? sectored_entries_0_4_data_1 : sectored_entries_0_4_data_0;
  assign _GEN_571 = 2'h2 == hitsVec_idx ? sectored_entries_0_4_data_2 : _GEN_570;
  assign _GEN_572 = 2'h3 == hitsVec_idx ? sectored_entries_0_4_data_3 : _GEN_571;
  assign _GEN_574 = 2'h1 == hitsVec_idx ? sectored_entries_0_5_data_1 : sectored_entries_0_5_data_0;
  assign _GEN_575 = 2'h2 == hitsVec_idx ? sectored_entries_0_5_data_2 : _GEN_574;
  assign _GEN_576 = 2'h3 == hitsVec_idx ? sectored_entries_0_5_data_3 : _GEN_575;
  assign _GEN_578 = 2'h1 == hitsVec_idx ? sectored_entries_0_6_data_1 : sectored_entries_0_6_data_0;
  assign _GEN_579 = 2'h2 == hitsVec_idx ? sectored_entries_0_6_data_2 : _GEN_578;
  assign _GEN_580 = 2'h3 == hitsVec_idx ? sectored_entries_0_6_data_3 : _GEN_579;
  assign _GEN_582 = 2'h1 == hitsVec_idx ? sectored_entries_0_7_data_1 : sectored_entries_0_7_data_0;
  assign _GEN_583 = 2'h2 == hitsVec_idx ? sectored_entries_0_7_data_2 : _GEN_582;
  assign _GEN_584 = 2'h3 == hitsVec_idx ? sectored_entries_0_7_data_3 : _GEN_583;
  assign ppn_hi = entries_barrier_8_io_y_ppn[19:18]; // @[TLB.scala 105:26]
  assign _ppn_T_1 = superpage_hits_ignore_1 ? vpn : 27'h0; // @[TLB.scala 108:28]
  assign _GEN_953 = {{7'd0}, entries_barrier_8_io_y_ppn}; // @[TLB.scala 108:47]
  assign _ppn_T_2 = _ppn_T_1 | _GEN_953; // @[TLB.scala 108:47]
  assign ppn_lo = _ppn_T_2[17:9]; // @[TLB.scala 108:58]
  assign _ppn_T_4 = vpn | _GEN_953; // @[TLB.scala 108:47]
  assign ppn_lo_1 = _ppn_T_4[8:0]; // @[TLB.scala 108:58]
  assign _ppn_T_5 = {ppn_hi,ppn_lo,ppn_lo_1}; // @[Cat.scala 30:58]
  assign ppn_hi_2 = entries_barrier_9_io_y_ppn[19:18]; // @[TLB.scala 105:26]
  assign _ppn_T_6 = superpage_hits_ignore_4 ? vpn : 27'h0; // @[TLB.scala 108:28]
  assign _GEN_955 = {{7'd0}, entries_barrier_9_io_y_ppn}; // @[TLB.scala 108:47]
  assign _ppn_T_7 = _ppn_T_6 | _GEN_955; // @[TLB.scala 108:47]
  assign ppn_lo_2 = _ppn_T_7[17:9]; // @[TLB.scala 108:58]
  assign _ppn_T_9 = vpn | _GEN_955; // @[TLB.scala 108:47]
  assign ppn_lo_3 = _ppn_T_9[8:0]; // @[TLB.scala 108:58]
  assign _ppn_T_10 = {ppn_hi_2,ppn_lo_2,ppn_lo_3}; // @[Cat.scala 30:58]
  assign ppn_hi_4 = entries_barrier_10_io_y_ppn[19:18]; // @[TLB.scala 105:26]
  assign _ppn_T_11 = superpage_hits_ignore_7 ? vpn : 27'h0; // @[TLB.scala 108:28]
  assign _GEN_957 = {{7'd0}, entries_barrier_10_io_y_ppn}; // @[TLB.scala 108:47]
  assign _ppn_T_12 = _ppn_T_11 | _GEN_957; // @[TLB.scala 108:47]
  assign ppn_lo_4 = _ppn_T_12[17:9]; // @[TLB.scala 108:58]
  assign _ppn_T_14 = vpn | _GEN_957; // @[TLB.scala 108:47]
  assign ppn_lo_5 = _ppn_T_14[8:0]; // @[TLB.scala 108:58]
  assign _ppn_T_15 = {ppn_hi_4,ppn_lo_4,ppn_lo_5}; // @[Cat.scala 30:58]
  assign ppn_hi_6 = entries_barrier_11_io_y_ppn[19:18]; // @[TLB.scala 105:26]
  assign _ppn_T_16 = superpage_hits_ignore_10 ? vpn : 27'h0; // @[TLB.scala 108:28]
  assign _GEN_959 = {{7'd0}, entries_barrier_11_io_y_ppn}; // @[TLB.scala 108:47]
  assign _ppn_T_17 = _ppn_T_16 | _GEN_959; // @[TLB.scala 108:47]
  assign ppn_lo_6 = _ppn_T_17[17:9]; // @[TLB.scala 108:58]
  assign _ppn_T_19 = vpn | _GEN_959; // @[TLB.scala 108:47]
  assign ppn_lo_7 = _ppn_T_19[8:0]; // @[TLB.scala 108:58]
  assign _ppn_T_20 = {ppn_hi_6,ppn_lo_6,ppn_lo_7}; // @[Cat.scala 30:58]
  assign ppn_hi_8 = entries_barrier_12_io_y_ppn[19:18]; // @[TLB.scala 105:26]
  assign _GEN_961 = {{7'd0}, entries_barrier_12_io_y_ppn}; // @[TLB.scala 108:47]
  assign _ppn_T_22 = _mpu_ppn_T_17 | _GEN_961; // @[TLB.scala 108:47]
  assign ppn_lo_8 = _ppn_T_22[17:9]; // @[TLB.scala 108:58]
  assign _ppn_T_24 = _mpu_ppn_T_19 | _GEN_961; // @[TLB.scala 108:47]
  assign ppn_lo_9 = _ppn_T_24[8:0]; // @[TLB.scala 108:58]
  assign _ppn_T_25 = {ppn_hi_8,ppn_lo_8,ppn_lo_9}; // @[Cat.scala 30:58]
  assign _ppn_T_27 = hitsVec_0 ? entries_barrier_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  assign _ppn_T_28 = hitsVec_1 ? entries_barrier_1_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  assign _ppn_T_29 = hitsVec_2 ? entries_barrier_2_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  assign _ppn_T_30 = hitsVec_3 ? entries_barrier_3_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  assign _ppn_T_31 = hitsVec_4 ? entries_barrier_4_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  assign _ppn_T_32 = hitsVec_5 ? entries_barrier_5_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  assign _ppn_T_33 = hitsVec_6 ? entries_barrier_6_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  assign _ppn_T_34 = hitsVec_7 ? entries_barrier_7_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  assign _ppn_T_35 = hitsVec_8 ? _ppn_T_5 : 20'h0; // @[Mux.scala 27:72]
  assign _ppn_T_36 = hitsVec_9 ? _ppn_T_10 : 20'h0; // @[Mux.scala 27:72]
  assign _ppn_T_37 = hitsVec_10 ? _ppn_T_15 : 20'h0; // @[Mux.scala 27:72]
  assign _ppn_T_38 = hitsVec_11 ? _ppn_T_20 : 20'h0; // @[Mux.scala 27:72]
  assign _ppn_T_39 = hitsVec_12 ? _ppn_T_25 : 20'h0; // @[Mux.scala 27:72]
  assign _ppn_T_40 = hits_hi ? vpn[19:0] : 20'h0; // @[Mux.scala 27:72]
  assign _ppn_T_41 = _ppn_T_27 | _ppn_T_28; // @[Mux.scala 27:72]
  assign _ppn_T_42 = _ppn_T_41 | _ppn_T_29; // @[Mux.scala 27:72]
  assign _ppn_T_43 = _ppn_T_42 | _ppn_T_30; // @[Mux.scala 27:72]
  assign _ppn_T_44 = _ppn_T_43 | _ppn_T_31; // @[Mux.scala 27:72]
  assign _ppn_T_45 = _ppn_T_44 | _ppn_T_32; // @[Mux.scala 27:72]
  assign _ppn_T_46 = _ppn_T_45 | _ppn_T_33; // @[Mux.scala 27:72]
  assign _ppn_T_47 = _ppn_T_46 | _ppn_T_34; // @[Mux.scala 27:72]
  assign _ppn_T_48 = _ppn_T_47 | _ppn_T_35; // @[Mux.scala 27:72]
  assign _ppn_T_49 = _ppn_T_48 | _ppn_T_36; // @[Mux.scala 27:72]
  assign _ppn_T_50 = _ppn_T_49 | _ppn_T_37; // @[Mux.scala 27:72]
  assign _ppn_T_51 = _ppn_T_50 | _ppn_T_38; // @[Mux.scala 27:72]
  assign _ppn_T_52 = _ppn_T_51 | _ppn_T_39; // @[Mux.scala 27:72]
  assign ppn = _ppn_T_52 | _ppn_T_40; // @[Mux.scala 27:72]
  assign ptw_ae_array_lo = {entries_barrier_5_io_y_ae,entries_barrier_4_io_y_ae,entries_barrier_3_io_y_ae,entries_barrier_2_io_y_ae,entries_barrier_1_io_y_ae,entries_barrier_io_y_ae}; // @[Cat.scala 30:58]
  assign ptw_ae_array = {1'h0,entries_barrier_12_io_y_ae,entries_barrier_11_io_y_ae,entries_barrier_10_io_y_ae,entries_barrier_9_io_y_ae,entries_barrier_8_io_y_ae,entries_barrier_7_io_y_ae,entries_barrier_6_io_y_ae,ptw_ae_array_lo}; // @[Cat.scala 30:58]
  assign _priv_rw_ok_T_1 = ~priv_s | io_ptw_status_sum; // @[TLB.scala 265:32]
  assign priv_rw_ok_lo = {entries_barrier_5_io_y_u,entries_barrier_4_io_y_u,entries_barrier_3_io_y_u,entries_barrier_2_io_y_u,entries_barrier_1_io_y_u,entries_barrier_io_y_u}; // @[Cat.scala 30:58]
  assign _priv_rw_ok_T_2 = {entries_barrier_12_io_y_u,entries_barrier_11_io_y_u,entries_barrier_10_io_y_u,entries_barrier_9_io_y_u,entries_barrier_8_io_y_u,entries_barrier_7_io_y_u,entries_barrier_6_io_y_u,priv_rw_ok_lo}; // @[Cat.scala 30:58]
  assign _priv_rw_ok_T_3 = _priv_rw_ok_T_1 ? _priv_rw_ok_T_2 : 13'h0; // @[TLB.scala 265:23]
  assign _priv_rw_ok_T_6 = priv_s ? ~_priv_rw_ok_T_2 : 13'h0; // @[TLB.scala 265:89]
  assign priv_rw_ok = _priv_rw_ok_T_3 | _priv_rw_ok_T_6; // @[TLB.scala 265:84]
  assign r_array_lo = {entries_barrier_5_io_y_sr,entries_barrier_4_io_y_sr,entries_barrier_3_io_y_sr,entries_barrier_2_io_y_sr,entries_barrier_1_io_y_sr,entries_barrier_io_y_sr}; // @[Cat.scala 30:58]
  assign _r_array_T = {entries_barrier_12_io_y_sr,entries_barrier_11_io_y_sr,entries_barrier_10_io_y_sr,entries_barrier_9_io_y_sr,entries_barrier_8_io_y_sr,entries_barrier_7_io_y_sr,entries_barrier_6_io_y_sr,r_array_lo}; // @[Cat.scala 30:58]
  assign r_array_lo_1 = {entries_barrier_5_io_y_sx,entries_barrier_4_io_y_sx,entries_barrier_3_io_y_sx,entries_barrier_2_io_y_sx,entries_barrier_1_io_y_sx,entries_barrier_io_y_sx}; // @[Cat.scala 30:58]
  assign _r_array_T_1 = {entries_barrier_12_io_y_sx,entries_barrier_11_io_y_sx,entries_barrier_10_io_y_sx,entries_barrier_9_io_y_sx,entries_barrier_8_io_y_sx,entries_barrier_7_io_y_sx,entries_barrier_6_io_y_sx,r_array_lo_1}; // @[Cat.scala 30:58]
  assign _r_array_T_2 = io_ptw_status_mxr ? _r_array_T_1 : 13'h0; // @[TLB.scala 267:73]
  assign _r_array_T_3 = _r_array_T | _r_array_T_2; // @[TLB.scala 267:68]
  assign r_array_lo_2 = priv_rw_ok & _r_array_T_3; // @[TLB.scala 267:40]
  assign r_array = {1'h1,r_array_lo_2}; // @[Cat.scala 30:58]
  assign w_array_lo = {entries_barrier_5_io_y_sw,entries_barrier_4_io_y_sw,entries_barrier_3_io_y_sw,entries_barrier_2_io_y_sw,entries_barrier_1_io_y_sw,entries_barrier_io_y_sw}; // @[Cat.scala 30:58]
  assign _w_array_T = {entries_barrier_12_io_y_sw,entries_barrier_11_io_y_sw,entries_barrier_10_io_y_sw,entries_barrier_9_io_y_sw,entries_barrier_8_io_y_sw,entries_barrier_7_io_y_sw,entries_barrier_6_io_y_sw,w_array_lo}; // @[Cat.scala 30:58]
  assign w_array_lo_1 = priv_rw_ok & _w_array_T; // @[TLB.scala 268:40]
  assign w_array = {1'h1,w_array_lo_1}; // @[Cat.scala 30:58]
  assign pr_array_hi = prot_r ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  assign pr_array_lo = {entries_barrier_5_io_y_pr,entries_barrier_4_io_y_pr,entries_barrier_3_io_y_pr,entries_barrier_2_io_y_pr,entries_barrier_1_io_y_pr,entries_barrier_io_y_pr}; // @[Cat.scala 30:58]
  assign _pr_array_T_1 = {pr_array_hi,entries_barrier_11_io_y_pr,entries_barrier_10_io_y_pr,entries_barrier_9_io_y_pr,entries_barrier_8_io_y_pr,entries_barrier_7_io_y_pr,entries_barrier_6_io_y_pr,pr_array_lo}; // @[Cat.scala 30:58]
  assign pr_array = _pr_array_T_1 & ~ptw_ae_array; // @[TLB.scala 270:87]
  assign pw_array_hi = prot_w ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  assign pw_array_lo = {entries_barrier_5_io_y_pw,entries_barrier_4_io_y_pw,entries_barrier_3_io_y_pw,entries_barrier_2_io_y_pw,entries_barrier_1_io_y_pw,entries_barrier_io_y_pw}; // @[Cat.scala 30:58]
  assign _pw_array_T_1 = {pw_array_hi,entries_barrier_11_io_y_pw,entries_barrier_10_io_y_pw,entries_barrier_9_io_y_pw,entries_barrier_8_io_y_pw,entries_barrier_7_io_y_pw,entries_barrier_6_io_y_pw,pw_array_lo}; // @[Cat.scala 30:58]
  assign pw_array = _pw_array_T_1 & ~ptw_ae_array; // @[TLB.scala 271:87]
  assign eff_array_hi = prot_eff ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  assign eff_array_lo = {entries_barrier_5_io_y_eff,entries_barrier_4_io_y_eff,entries_barrier_3_io_y_eff,entries_barrier_2_io_y_eff,entries_barrier_1_io_y_eff,entries_barrier_io_y_eff}; // @[Cat.scala 30:58]
  assign eff_array = {eff_array_hi,entries_barrier_11_io_y_eff,entries_barrier_10_io_y_eff,entries_barrier_9_io_y_eff,entries_barrier_8_io_y_eff,entries_barrier_7_io_y_eff,entries_barrier_6_io_y_eff,eff_array_lo}; // @[Cat.scala 30:58]
  assign c_array_hi = cacheable ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  assign c_array_lo = {entries_barrier_5_io_y_c,entries_barrier_4_io_y_c,entries_barrier_3_io_y_c,entries_barrier_2_io_y_c,entries_barrier_1_io_y_c,entries_barrier_io_y_c}; // @[Cat.scala 30:58]
  assign c_array = {c_array_hi,entries_barrier_11_io_y_c,entries_barrier_10_io_y_c,entries_barrier_9_io_y_c,entries_barrier_8_io_y_c,entries_barrier_7_io_y_c,entries_barrier_6_io_y_c,c_array_lo}; // @[Cat.scala 30:58]
  assign ppp_array_hi = _prot_w_T_31 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  assign ppp_array_lo = {entries_barrier_5_io_y_ppp,entries_barrier_4_io_y_ppp,entries_barrier_3_io_y_ppp,entries_barrier_2_io_y_ppp,entries_barrier_1_io_y_ppp,entries_barrier_io_y_ppp}; // @[Cat.scala 30:58]
  assign ppp_array = {ppp_array_hi,entries_barrier_11_io_y_ppp,entries_barrier_10_io_y_ppp,entries_barrier_9_io_y_ppp,entries_barrier_8_io_y_ppp,entries_barrier_7_io_y_ppp,entries_barrier_6_io_y_ppp,ppp_array_lo}; // @[Cat.scala 30:58]
  assign paa_array_hi = prot_al ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  assign paa_array_lo = {entries_barrier_5_io_y_paa,entries_barrier_4_io_y_paa,entries_barrier_3_io_y_paa,entries_barrier_2_io_y_paa,entries_barrier_1_io_y_paa,entries_barrier_io_y_paa}; // @[Cat.scala 30:58]
  assign paa_array = {paa_array_hi,entries_barrier_11_io_y_paa,entries_barrier_10_io_y_paa,entries_barrier_9_io_y_paa,entries_barrier_8_io_y_paa,entries_barrier_7_io_y_paa,entries_barrier_6_io_y_paa,paa_array_lo}; // @[Cat.scala 30:58]
  assign pal_array_lo = {entries_barrier_5_io_y_pal,entries_barrier_4_io_y_pal,entries_barrier_3_io_y_pal,entries_barrier_2_io_y_pal,entries_barrier_1_io_y_pal,entries_barrier_io_y_pal}; // @[Cat.scala 30:58]
  assign pal_array = {paa_array_hi,entries_barrier_11_io_y_pal,entries_barrier_10_io_y_pal,entries_barrier_9_io_y_pal,entries_barrier_8_io_y_pal,entries_barrier_7_io_y_pal,entries_barrier_6_io_y_pal,pal_array_lo}; // @[Cat.scala 30:58]
  assign ppp_array_if_cached = ppp_array | c_array; // @[TLB.scala 278:39]
  assign paa_array_if_cached = paa_array | c_array; // @[TLB.scala 279:39]
  assign pal_array_if_cached = pal_array | c_array; // @[TLB.scala 280:39]
  assign _misaligned_T = 4'h1 << io_req_bits_size; // @[OneHot.scala 58:35]
  assign _misaligned_T_2 = _misaligned_T - 4'h1; // @[TLB.scala 283:69]
  assign _GEN_963 = {{36'd0}, _misaligned_T_2}; // @[TLB.scala 283:39]
  assign _misaligned_T_3 = io_req_bits_vaddr & _GEN_963; // @[TLB.scala 283:39]
  assign misaligned = |_misaligned_T_3; // @[TLB.scala 283:75]
  assign bad_va_maskedVAddr = io_req_bits_vaddr & 40'hc000000000; // @[TLB.scala 289:43]
  assign _bad_va_T_1 = bad_va_maskedVAddr == 40'h0; // @[TLB.scala 290:61]
  assign _bad_va_T_2 = bad_va_maskedVAddr == 40'hc000000000; // @[TLB.scala 290:82]
  assign _bad_va_T_3 = _bad_va_T_1 | _bad_va_T_2; // @[TLB.scala 290:67]
  assign bad_va = vm_enabled & ~_bad_va_T_3; // @[TLB.scala 284:117]
  assign _cmd_lrsc_T = io_req_bits_cmd == 5'h6; // @[package.scala 15:47]
  assign _cmd_lrsc_T_1 = io_req_bits_cmd == 5'h7; // @[package.scala 15:47]
  assign cmd_lrsc = _cmd_lrsc_T | _cmd_lrsc_T_1; // @[package.scala 72:59]
  assign _cmd_amo_logical_T = io_req_bits_cmd == 5'h4; // @[package.scala 15:47]
  assign _cmd_amo_logical_T_1 = io_req_bits_cmd == 5'h9; // @[package.scala 15:47]
  assign _cmd_amo_logical_T_2 = io_req_bits_cmd == 5'ha; // @[package.scala 15:47]
  assign _cmd_amo_logical_T_3 = io_req_bits_cmd == 5'hb; // @[package.scala 15:47]
  assign _cmd_amo_logical_T_4 = _cmd_amo_logical_T | _cmd_amo_logical_T_1; // @[package.scala 72:59]
  assign _cmd_amo_logical_T_5 = _cmd_amo_logical_T_4 | _cmd_amo_logical_T_2; // @[package.scala 72:59]
  assign cmd_amo_logical = _cmd_amo_logical_T_5 | _cmd_amo_logical_T_3; // @[package.scala 72:59]
  assign _cmd_amo_arithmetic_T = io_req_bits_cmd == 5'h8; // @[package.scala 15:47]
  assign _cmd_amo_arithmetic_T_1 = io_req_bits_cmd == 5'hc; // @[package.scala 15:47]
  assign _cmd_amo_arithmetic_T_2 = io_req_bits_cmd == 5'hd; // @[package.scala 15:47]
  assign _cmd_amo_arithmetic_T_3 = io_req_bits_cmd == 5'he; // @[package.scala 15:47]
  assign _cmd_amo_arithmetic_T_4 = io_req_bits_cmd == 5'hf; // @[package.scala 15:47]
  assign _cmd_amo_arithmetic_T_5 = _cmd_amo_arithmetic_T | _cmd_amo_arithmetic_T_1; // @[package.scala 72:59]
  assign _cmd_amo_arithmetic_T_6 = _cmd_amo_arithmetic_T_5 | _cmd_amo_arithmetic_T_2; // @[package.scala 72:59]
  assign _cmd_amo_arithmetic_T_7 = _cmd_amo_arithmetic_T_6 | _cmd_amo_arithmetic_T_3; // @[package.scala 72:59]
  assign cmd_amo_arithmetic = _cmd_amo_arithmetic_T_7 | _cmd_amo_arithmetic_T_4; // @[package.scala 72:59]
  assign cmd_put_partial = io_req_bits_cmd == 5'h11; // @[TLB.scala 297:41]
  assign _cmd_read_T = io_req_bits_cmd == 5'h0; // @[Consts.scala 81:31]
  assign _cmd_read_T_2 = _cmd_read_T | _cmd_lrsc_T; // @[Consts.scala 81:41]
  assign _cmd_read_T_4 = _cmd_read_T_2 | _cmd_lrsc_T_1; // @[Consts.scala 81:58]
  assign _cmd_read_T_21 = cmd_amo_logical | cmd_amo_arithmetic; // @[Consts.scala 79:44]
  assign cmd_read = _cmd_read_T_4 | _cmd_read_T_21; // @[Consts.scala 81:75]
  assign _cmd_write_T = io_req_bits_cmd == 5'h1; // @[Consts.scala 82:32]
  assign _cmd_write_T_2 = _cmd_write_T | cmd_put_partial; // @[Consts.scala 82:42]
  assign _cmd_write_T_4 = _cmd_write_T_2 | _cmd_lrsc_T_1; // @[Consts.scala 82:59]
  assign cmd_write = _cmd_write_T_4 | _cmd_read_T_21; // @[Consts.scala 82:76]
  assign _cmd_write_perms_T = io_req_bits_cmd == 5'h5; // @[package.scala 15:47]
  assign _cmd_write_perms_T_1 = io_req_bits_cmd == 5'h17; // @[package.scala 15:47]
  assign _cmd_write_perms_T_2 = _cmd_write_perms_T | _cmd_write_perms_T_1; // @[package.scala 72:59]
  assign cmd_write_perms = cmd_write | _cmd_write_perms_T_2; // @[TLB.scala 300:35]
  assign _ae_array_T = misaligned ? eff_array : 14'h0; // @[TLB.scala 305:8]
  assign _ae_array_T_2 = cmd_lrsc ? ~c_array : 14'h0; // @[TLB.scala 306:8]
  assign ae_array = _ae_array_T | _ae_array_T_2; // @[TLB.scala 305:37]
  assign _ae_ld_array_T_1 = ae_array | ~pr_array; // @[TLB.scala 307:44]
  assign ae_ld_array = cmd_read ? _ae_ld_array_T_1 : 14'h0; // @[TLB.scala 307:24]
  assign _ae_st_array_T_1 = ae_array | ~pw_array; // @[TLB.scala 309:35]
  assign _ae_st_array_T_2 = cmd_write_perms ? _ae_st_array_T_1 : 14'h0; // @[TLB.scala 309:8]
  assign _ae_st_array_T_4 = cmd_put_partial ? ~ppp_array_if_cached : 14'h0; // @[TLB.scala 310:8]
  assign _ae_st_array_T_5 = _ae_st_array_T_2 | _ae_st_array_T_4; // @[TLB.scala 309:53]
  assign _ae_st_array_T_7 = cmd_amo_logical ? ~pal_array_if_cached : 14'h0; // @[TLB.scala 311:8]
  assign _ae_st_array_T_8 = _ae_st_array_T_5 | _ae_st_array_T_7; // @[TLB.scala 310:53]
  assign _ae_st_array_T_10 = cmd_amo_arithmetic ? ~paa_array_if_cached : 14'h0; // @[TLB.scala 312:8]
  assign ae_st_array = _ae_st_array_T_8 | _ae_st_array_T_10; // @[TLB.scala 311:53]
  assign _ma_ld_array_T = misaligned & cmd_read; // @[TLB.scala 318:36]
  assign ma_ld_array = _ma_ld_array_T ? ~eff_array : 14'h0; // @[TLB.scala 318:24]
  assign _ma_st_array_T = misaligned & cmd_write; // @[TLB.scala 319:36]
  assign ma_st_array = _ma_st_array_T ? ~eff_array : 14'h0; // @[TLB.scala 319:24]
  assign _pf_ld_array_T = r_array | ptw_ae_array; // @[TLB.scala 320:45]
  assign pf_ld_array = cmd_read ? ~_pf_ld_array_T : 14'h0; // @[TLB.scala 320:24]
  assign _pf_st_array_T = w_array | ptw_ae_array; // @[TLB.scala 321:52]
  assign pf_st_array = cmd_write_perms ? ~_pf_st_array_T : 14'h0; // @[TLB.scala 321:24]
  assign tlb_hit = |real_hits; // @[TLB.scala 324:27]
  assign _tlb_miss_T_1 = vm_enabled & ~bad_va; // @[TLB.scala 325:29]
  assign tlb_miss = _tlb_miss_T_1 & ~tlb_hit; // @[TLB.scala 325:40]
  assign _T_23 = io_req_valid & vm_enabled; // @[TLB.scala 329:22]
  assign _T_24 = sector_hits_0 | sector_hits_1; // @[package.scala 72:59]
  assign _T_25 = _T_24 | sector_hits_2; // @[package.scala 72:59]
  assign _T_26 = _T_25 | sector_hits_3; // @[package.scala 72:59]
  assign _T_27 = _T_26 | sector_hits_4; // @[package.scala 72:59]
  assign _T_28 = _T_27 | sector_hits_5; // @[package.scala 72:59]
  assign _T_29 = _T_28 | sector_hits_6; // @[package.scala 72:59]
  assign _T_30 = _T_29 | sector_hits_7; // @[package.scala 72:59]
  assign _T_31 = {sector_hits_7,sector_hits_6,sector_hits_5,sector_hits_4,sector_hits_3,sector_hits_2,sector_hits_1,sector_hits_0}; // @[Cat.scala 30:58]
  assign hi_1 = _T_31[7:4]; // @[OneHot.scala 30:18]
  assign lo_1 = _T_31[3:0]; // @[OneHot.scala 31:18]
  assign hi_2 = |hi_1; // @[OneHot.scala 32:14]
  assign _T_32 = hi_1 | lo_1; // @[OneHot.scala 32:28]
  assign hi_3 = _T_32[3:2]; // @[OneHot.scala 30:18]
  assign lo_2 = _T_32[1:0]; // @[OneHot.scala 31:18]
  assign hi_4 = |hi_3; // @[OneHot.scala 32:14]
  assign _T_33 = hi_3 | lo_2; // @[OneHot.scala 32:28]
  assign lo_3 = _T_33[1]; // @[CircuitMath.scala 30:8]
  assign state_vec_0_touch_way_sized = {hi_2,hi_4,lo_3}; // @[Cat.scala 30:58]
  assign state_vec_0_hi_hi = ~state_vec_0_touch_way_sized[2]; // @[Replacement.scala 196:33]
  assign state_vec_0_left_subtree_state = state_vec_0[5:3]; // @[package.scala 154:13]
  assign state_vec_0_right_subtree_state = state_vec_0[2:0]; // @[Replacement.scala 198:38]
  assign state_vec_0_hi_hi_1 = ~state_vec_0_touch_way_sized[1]; // @[Replacement.scala 196:33]
  assign state_vec_0_left_subtree_state_1 = state_vec_0_left_subtree_state[1]; // @[package.scala 154:13]
  assign state_vec_0_right_subtree_state_1 = state_vec_0_left_subtree_state[0]; // @[Replacement.scala 198:38]
  assign state_vec_0_hi_lo = state_vec_0_hi_hi_1 ? state_vec_0_left_subtree_state_1 : ~state_vec_0_touch_way_sized[0]; // @[Replacement.scala 203:16]
  assign state_vec_0_lo = state_vec_0_hi_hi_1 ? ~state_vec_0_touch_way_sized[0] : state_vec_0_right_subtree_state_1; // @[Replacement.scala 206:16]
  assign _state_vec_0_T_7 = {state_vec_0_hi_hi_1,state_vec_0_hi_lo,state_vec_0_lo}; // @[Cat.scala 30:58]
  assign state_vec_0_hi_lo_1 = state_vec_0_hi_hi ? state_vec_0_left_subtree_state : _state_vec_0_T_7; // @[Replacement.scala 203:16]
  assign state_vec_0_left_subtree_state_2 = state_vec_0_right_subtree_state[1]; // @[package.scala 154:13]
  assign state_vec_0_right_subtree_state_2 = state_vec_0_right_subtree_state[0]; // @[Replacement.scala 198:38]
  assign state_vec_0_hi_lo_2 = state_vec_0_hi_hi_1 ? state_vec_0_left_subtree_state_2 : ~state_vec_0_touch_way_sized[0]; // @[Replacement.scala 203:16]
  assign state_vec_0_lo_1 = state_vec_0_hi_hi_1 ? ~state_vec_0_touch_way_sized[0] : state_vec_0_right_subtree_state_2; // @[Replacement.scala 206:16]
  assign _state_vec_0_T_15 = {state_vec_0_hi_hi_1,state_vec_0_hi_lo_2,state_vec_0_lo_1}; // @[Cat.scala 30:58]
  assign state_vec_0_lo_2 = state_vec_0_hi_hi ? _state_vec_0_T_15 : state_vec_0_right_subtree_state; // @[Replacement.scala 206:16]
  assign _state_vec_0_T_16 = {state_vec_0_hi_hi,state_vec_0_hi_lo_1,state_vec_0_lo_2}; // @[Cat.scala 30:58]
  assign _T_35 = superpage_hits_0 | superpage_hits_1; // @[package.scala 72:59]
  assign _T_36 = _T_35 | superpage_hits_2; // @[package.scala 72:59]
  assign _T_37 = _T_36 | superpage_hits_3; // @[package.scala 72:59]
  assign _T_38 = {superpage_hits_3,superpage_hits_2,superpage_hits_1,superpage_hits_0}; // @[Cat.scala 30:58]
  assign hi_6 = _T_38[3:2]; // @[OneHot.scala 30:18]
  assign lo_6 = _T_38[1:0]; // @[OneHot.scala 31:18]
  assign hi_7 = |hi_6; // @[OneHot.scala 32:14]
  assign _T_39 = hi_6 | lo_6; // @[OneHot.scala 32:28]
  assign lo_7 = _T_39[1]; // @[CircuitMath.scala 30:8]
  assign state_reg_touch_way_sized = {hi_7,lo_7}; // @[Cat.scala 30:58]
  assign state_reg_hi_hi = ~state_reg_touch_way_sized[1]; // @[Replacement.scala 196:33]
  assign state_reg_left_subtree_state = state_reg_1[1]; // @[package.scala 154:13]
  assign state_reg_right_subtree_state = state_reg_1[0]; // @[Replacement.scala 198:38]
  assign state_reg_hi_lo = state_reg_hi_hi ? state_reg_left_subtree_state : ~state_reg_touch_way_sized[0]; // @[Replacement.scala 203:16]
  assign state_reg_lo = state_reg_hi_hi ? ~state_reg_touch_way_sized[0] : state_reg_right_subtree_state; // @[Replacement.scala 206:16]
  assign _state_reg_T_6 = {state_reg_hi_hi,state_reg_hi_lo,state_reg_lo}; // @[Cat.scala 30:58]
  assign multipleHits_leftOne = real_hits[0]; // @[Misc.scala 180:37]
  assign multipleHits_leftOne_1 = real_hits[1]; // @[Misc.scala 180:37]
  assign multipleHits_rightOne = real_hits[2]; // @[Misc.scala 181:39]
  assign multipleHits_rightOne_1 = multipleHits_leftOne_1 | multipleHits_rightOne; // @[Misc.scala 182:16]
  assign multipleHits_rightTwo = multipleHits_leftOne_1 & multipleHits_rightOne; // @[Misc.scala 182:61]
  assign multipleHits_leftOne_2 = multipleHits_leftOne | multipleHits_rightOne_1; // @[Misc.scala 182:16]
  assign _multipleHits_T_9 = multipleHits_leftOne & multipleHits_rightOne_1; // @[Misc.scala 182:61]
  assign multipleHits_leftTwo = multipleHits_rightTwo | _multipleHits_T_9; // @[Misc.scala 182:49]
  assign multipleHits_leftOne_3 = real_hits[3]; // @[Misc.scala 180:37]
  assign multipleHits_leftOne_4 = real_hits[4]; // @[Misc.scala 180:37]
  assign multipleHits_rightOne_2 = real_hits[5]; // @[Misc.scala 181:39]
  assign multipleHits_rightOne_3 = multipleHits_leftOne_4 | multipleHits_rightOne_2; // @[Misc.scala 182:16]
  assign multipleHits_rightTwo_1 = multipleHits_leftOne_4 & multipleHits_rightOne_2; // @[Misc.scala 182:61]
  assign multipleHits_rightOne_4 = multipleHits_leftOne_3 | multipleHits_rightOne_3; // @[Misc.scala 182:16]
  assign _multipleHits_T_18 = multipleHits_leftOne_3 & multipleHits_rightOne_3; // @[Misc.scala 182:61]
  assign multipleHits_rightTwo_2 = multipleHits_rightTwo_1 | _multipleHits_T_18; // @[Misc.scala 182:49]
  assign multipleHits_leftOne_5 = multipleHits_leftOne_2 | multipleHits_rightOne_4; // @[Misc.scala 182:16]
  assign _multipleHits_T_19 = multipleHits_leftTwo | multipleHits_rightTwo_2; // @[Misc.scala 182:37]
  assign _multipleHits_T_20 = multipleHits_leftOne_2 & multipleHits_rightOne_4; // @[Misc.scala 182:61]
  assign multipleHits_leftTwo_1 = _multipleHits_T_19 | _multipleHits_T_20; // @[Misc.scala 182:49]
  assign multipleHits_leftOne_6 = real_hits[6]; // @[Misc.scala 180:37]
  assign multipleHits_leftOne_7 = real_hits[7]; // @[Misc.scala 180:37]
  assign multipleHits_rightOne_5 = real_hits[8]; // @[Misc.scala 181:39]
  assign multipleHits_rightOne_6 = multipleHits_leftOne_7 | multipleHits_rightOne_5; // @[Misc.scala 182:16]
  assign multipleHits_rightTwo_3 = multipleHits_leftOne_7 & multipleHits_rightOne_5; // @[Misc.scala 182:61]
  assign multipleHits_leftOne_8 = multipleHits_leftOne_6 | multipleHits_rightOne_6; // @[Misc.scala 182:16]
  assign _multipleHits_T_30 = multipleHits_leftOne_6 & multipleHits_rightOne_6; // @[Misc.scala 182:61]
  assign multipleHits_leftTwo_2 = multipleHits_rightTwo_3 | _multipleHits_T_30; // @[Misc.scala 182:49]
  assign multipleHits_leftOne_9 = real_hits[9]; // @[Misc.scala 180:37]
  assign multipleHits_rightOne_7 = real_hits[10]; // @[Misc.scala 181:39]
  assign multipleHits_leftOne_10 = multipleHits_leftOne_9 | multipleHits_rightOne_7; // @[Misc.scala 182:16]
  assign multipleHits_leftTwo_3 = multipleHits_leftOne_9 & multipleHits_rightOne_7; // @[Misc.scala 182:61]
  assign multipleHits_leftOne_11 = real_hits[11]; // @[Misc.scala 180:37]
  assign multipleHits_rightOne_8 = real_hits[12]; // @[Misc.scala 181:39]
  assign multipleHits_rightOne_9 = multipleHits_leftOne_11 | multipleHits_rightOne_8; // @[Misc.scala 182:16]
  assign multipleHits_rightTwo_4 = multipleHits_leftOne_11 & multipleHits_rightOne_8; // @[Misc.scala 182:61]
  assign multipleHits_rightOne_10 = multipleHits_leftOne_10 | multipleHits_rightOne_9; // @[Misc.scala 182:16]
  assign _multipleHits_T_42 = multipleHits_leftTwo_3 | multipleHits_rightTwo_4; // @[Misc.scala 182:37]
  assign _multipleHits_T_43 = multipleHits_leftOne_10 & multipleHits_rightOne_9; // @[Misc.scala 182:61]
  assign multipleHits_rightTwo_5 = _multipleHits_T_42 | _multipleHits_T_43; // @[Misc.scala 182:49]
  assign multipleHits_rightOne_11 = multipleHits_leftOne_8 | multipleHits_rightOne_10; // @[Misc.scala 182:16]
  assign _multipleHits_T_44 = multipleHits_leftTwo_2 | multipleHits_rightTwo_5; // @[Misc.scala 182:37]
  assign _multipleHits_T_45 = multipleHits_leftOne_8 & multipleHits_rightOne_10; // @[Misc.scala 182:61]
  assign multipleHits_rightTwo_6 = _multipleHits_T_44 | _multipleHits_T_45; // @[Misc.scala 182:49]
  assign _multipleHits_T_47 = multipleHits_leftTwo_1 | multipleHits_rightTwo_6; // @[Misc.scala 182:37]
  assign _multipleHits_T_48 = multipleHits_leftOne_5 & multipleHits_rightOne_11; // @[Misc.scala 182:61]
  assign multipleHits = _multipleHits_T_47 | _multipleHits_T_48; // @[Misc.scala 182:49]
  assign _io_resp_pf_ld_T = bad_va & cmd_read; // @[TLB.scala 342:28]
  assign _io_resp_pf_ld_T_1 = pf_ld_array & hits; // @[TLB.scala 342:57]
  assign _io_resp_pf_ld_T_2 = |_io_resp_pf_ld_T_1; // @[TLB.scala 342:65]
  assign _io_resp_pf_st_T = bad_va & cmd_write_perms; // @[TLB.scala 343:28]
  assign _io_resp_pf_st_T_1 = pf_st_array & hits; // @[TLB.scala 343:64]
  assign _io_resp_pf_st_T_2 = |_io_resp_pf_st_T_1; // @[TLB.scala 343:72]
  assign _io_resp_ae_ld_T = ae_ld_array & hits; // @[TLB.scala 345:33]
  assign _io_resp_ae_st_T = ae_st_array & hits; // @[TLB.scala 346:33]
  assign _io_resp_ma_ld_T = ma_ld_array & hits; // @[TLB.scala 348:33]
  assign _io_resp_ma_st_T = ma_st_array & hits; // @[TLB.scala 349:33]
  assign _io_resp_cacheable_T = c_array & hits; // @[TLB.scala 351:33]
  assign _io_resp_miss_T = io_ptw_resp_valid | tlb_miss; // @[TLB.scala 354:29]
  assign _T_41 = io_req_ready & io_req_valid; // @[Decoupled.scala 40:37]
  assign _T_42 = _T_41 & tlb_miss; // @[TLB.scala 363:25]
  assign r_superpage_repl_addr_hi = state_reg_1[2]; // @[Replacement.scala 243:38]
  assign r_superpage_repl_addr_lo = r_superpage_repl_addr_hi ? state_reg_left_subtree_state : state_reg_right_subtree_state; // @[Replacement.scala 250:16]
  assign _r_superpage_repl_addr_T_2 = {r_superpage_repl_addr_hi,r_superpage_repl_addr_lo}; // @[Cat.scala 30:58]
  assign r_superpage_repl_addr_valids = {superpage_entries_3_valid_0,superpage_entries_2_valid_0,superpage_entries_1_valid_0,superpage_entries_0_valid_0}; // @[Cat.scala 30:58]
  assign _r_superpage_repl_addr_T_3 = &r_superpage_repl_addr_valids; // @[TLB.scala 411:16]
  assign _r_superpage_repl_addr_T_5 = ~r_superpage_repl_addr_valids[0]; // @[OneHot.scala 47:40]
  assign _r_superpage_repl_addr_T_6 = ~r_superpage_repl_addr_valids[1]; // @[OneHot.scala 47:40]
  assign _r_superpage_repl_addr_T_7 = ~r_superpage_repl_addr_valids[2]; // @[OneHot.scala 47:40]
  assign r_sectored_repl_addr_hi = state_vec_0[6]; // @[Replacement.scala 243:38]
  assign r_sectored_repl_addr_hi_1 = state_vec_0_left_subtree_state[2]; // @[Replacement.scala 243:38]
  assign r_sectored_repl_addr_lo = r_sectored_repl_addr_hi_1 ? state_vec_0_left_subtree_state_1 : state_vec_0_right_subtree_state_1; // @[Replacement.scala 250:16]
  assign _r_sectored_repl_addr_T_2 = {r_sectored_repl_addr_hi_1,r_sectored_repl_addr_lo}; // @[Cat.scala 30:58]
  assign r_sectored_repl_addr_hi_2 = state_vec_0_right_subtree_state[2]; // @[Replacement.scala 243:38]
  assign r_sectored_repl_addr_lo_1 = r_sectored_repl_addr_hi_2 ? state_vec_0_left_subtree_state_2 : state_vec_0_right_subtree_state_2; // @[Replacement.scala 250:16]
  assign _r_sectored_repl_addr_T_5 = {r_sectored_repl_addr_hi_2,r_sectored_repl_addr_lo_1}; // @[Cat.scala 30:58]
  assign r_sectored_repl_addr_lo_2 = r_sectored_repl_addr_hi ? _r_sectored_repl_addr_T_2 : _r_sectored_repl_addr_T_5; // @[Replacement.scala 250:16]
  assign _r_sectored_repl_addr_T_6 = {r_sectored_repl_addr_hi,r_sectored_repl_addr_lo_2}; // @[Cat.scala 30:58]
  assign r_sectored_repl_addr_valids = {_sector_hits_T_44,_sector_hits_T_38,_sector_hits_T_32,_sector_hits_T_26,_sector_hits_T_20,_sector_hits_T_14,_sector_hits_T_8,_sector_hits_T_2}; // @[Cat.scala 30:58]
  assign _r_sectored_repl_addr_T_7 = &r_sectored_repl_addr_valids; // @[TLB.scala 411:16]
  assign _r_sectored_repl_addr_T_9 = ~r_sectored_repl_addr_valids[0]; // @[OneHot.scala 47:40]
  assign _r_sectored_repl_addr_T_10 = ~r_sectored_repl_addr_valids[1]; // @[OneHot.scala 47:40]
  assign _r_sectored_repl_addr_T_11 = ~r_sectored_repl_addr_valids[2]; // @[OneHot.scala 47:40]
  assign _r_sectored_repl_addr_T_12 = ~r_sectored_repl_addr_valids[3]; // @[OneHot.scala 47:40]
  assign _r_sectored_repl_addr_T_13 = ~r_sectored_repl_addr_valids[4]; // @[OneHot.scala 47:40]
  assign _r_sectored_repl_addr_T_14 = ~r_sectored_repl_addr_valids[5]; // @[OneHot.scala 47:40]
  assign _r_sectored_repl_addr_T_15 = ~r_sectored_repl_addr_valids[6]; // @[OneHot.scala 47:40]
  assign _T_44 = state == 2'h2; // @[TLB.scala 377:17]
  assign _T_45 = _T_44 & io_sfence_valid; // @[TLB.scala 377:28]
  assign _T_48 = io_sfence_bits_addr[38:12] == vpn; // @[TLB.scala 385:72]
  assign _T_49 = ~io_sfence_bits_rs1 | _T_48; // @[TLB.scala 385:34]
  assign _T_51 = _T_49 | reset; // @[TLB.scala 385:13]
  assign _T_59 = _sector_hits_T_3[26:18] == 9'h0; // @[TLB.scala 134:61]
  assign _GEN_617 = sectored_entries_0_0_data_0[13] ? _GEN_473 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_618 = sectored_entries_0_0_data_1[13] ? _GEN_474 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_619 = sectored_entries_0_0_data_2[13] ? _GEN_475 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_620 = sectored_entries_0_0_data_3[13] ? _GEN_476 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_621 = io_sfence_bits_rs2 & _GEN_617; // @[TLB.scala 388:40]
  assign _GEN_622 = io_sfence_bits_rs2 & _GEN_618; // @[TLB.scala 388:40]
  assign _GEN_623 = io_sfence_bits_rs2 & _GEN_619; // @[TLB.scala 388:40]
  assign _GEN_624 = io_sfence_bits_rs2 & _GEN_620; // @[TLB.scala 388:40]
  assign _T_198 = _sector_hits_T_9[26:18] == 9'h0; // @[TLB.scala 134:61]
  assign _GEN_645 = sectored_entries_0_1_data_0[13] ? _GEN_483 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_646 = sectored_entries_0_1_data_1[13] ? _GEN_484 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_647 = sectored_entries_0_1_data_2[13] ? _GEN_485 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_648 = sectored_entries_0_1_data_3[13] ? _GEN_486 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_649 = io_sfence_bits_rs2 & _GEN_645; // @[TLB.scala 388:40]
  assign _GEN_650 = io_sfence_bits_rs2 & _GEN_646; // @[TLB.scala 388:40]
  assign _GEN_651 = io_sfence_bits_rs2 & _GEN_647; // @[TLB.scala 388:40]
  assign _GEN_652 = io_sfence_bits_rs2 & _GEN_648; // @[TLB.scala 388:40]
  assign _T_337 = _sector_hits_T_15[26:18] == 9'h0; // @[TLB.scala 134:61]
  assign _GEN_673 = sectored_entries_0_2_data_0[13] ? _GEN_493 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_674 = sectored_entries_0_2_data_1[13] ? _GEN_494 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_675 = sectored_entries_0_2_data_2[13] ? _GEN_495 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_676 = sectored_entries_0_2_data_3[13] ? _GEN_496 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_677 = io_sfence_bits_rs2 & _GEN_673; // @[TLB.scala 388:40]
  assign _GEN_678 = io_sfence_bits_rs2 & _GEN_674; // @[TLB.scala 388:40]
  assign _GEN_679 = io_sfence_bits_rs2 & _GEN_675; // @[TLB.scala 388:40]
  assign _GEN_680 = io_sfence_bits_rs2 & _GEN_676; // @[TLB.scala 388:40]
  assign _T_476 = _sector_hits_T_21[26:18] == 9'h0; // @[TLB.scala 134:61]
  assign _GEN_701 = sectored_entries_0_3_data_0[13] ? _GEN_503 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_702 = sectored_entries_0_3_data_1[13] ? _GEN_504 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_703 = sectored_entries_0_3_data_2[13] ? _GEN_505 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_704 = sectored_entries_0_3_data_3[13] ? _GEN_506 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_705 = io_sfence_bits_rs2 & _GEN_701; // @[TLB.scala 388:40]
  assign _GEN_706 = io_sfence_bits_rs2 & _GEN_702; // @[TLB.scala 388:40]
  assign _GEN_707 = io_sfence_bits_rs2 & _GEN_703; // @[TLB.scala 388:40]
  assign _GEN_708 = io_sfence_bits_rs2 & _GEN_704; // @[TLB.scala 388:40]
  assign _T_615 = _sector_hits_T_27[26:18] == 9'h0; // @[TLB.scala 134:61]
  assign _GEN_729 = sectored_entries_0_4_data_0[13] ? _GEN_513 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_730 = sectored_entries_0_4_data_1[13] ? _GEN_514 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_731 = sectored_entries_0_4_data_2[13] ? _GEN_515 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_732 = sectored_entries_0_4_data_3[13] ? _GEN_516 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_733 = io_sfence_bits_rs2 & _GEN_729; // @[TLB.scala 388:40]
  assign _GEN_734 = io_sfence_bits_rs2 & _GEN_730; // @[TLB.scala 388:40]
  assign _GEN_735 = io_sfence_bits_rs2 & _GEN_731; // @[TLB.scala 388:40]
  assign _GEN_736 = io_sfence_bits_rs2 & _GEN_732; // @[TLB.scala 388:40]
  assign _T_754 = _sector_hits_T_33[26:18] == 9'h0; // @[TLB.scala 134:61]
  assign _GEN_757 = sectored_entries_0_5_data_0[13] ? _GEN_523 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_758 = sectored_entries_0_5_data_1[13] ? _GEN_524 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_759 = sectored_entries_0_5_data_2[13] ? _GEN_525 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_760 = sectored_entries_0_5_data_3[13] ? _GEN_526 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_761 = io_sfence_bits_rs2 & _GEN_757; // @[TLB.scala 388:40]
  assign _GEN_762 = io_sfence_bits_rs2 & _GEN_758; // @[TLB.scala 388:40]
  assign _GEN_763 = io_sfence_bits_rs2 & _GEN_759; // @[TLB.scala 388:40]
  assign _GEN_764 = io_sfence_bits_rs2 & _GEN_760; // @[TLB.scala 388:40]
  assign _T_893 = _sector_hits_T_39[26:18] == 9'h0; // @[TLB.scala 134:61]
  assign _GEN_785 = sectored_entries_0_6_data_0[13] ? _GEN_533 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_786 = sectored_entries_0_6_data_1[13] ? _GEN_534 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_787 = sectored_entries_0_6_data_2[13] ? _GEN_535 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_788 = sectored_entries_0_6_data_3[13] ? _GEN_536 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_789 = io_sfence_bits_rs2 & _GEN_785; // @[TLB.scala 388:40]
  assign _GEN_790 = io_sfence_bits_rs2 & _GEN_786; // @[TLB.scala 388:40]
  assign _GEN_791 = io_sfence_bits_rs2 & _GEN_787; // @[TLB.scala 388:40]
  assign _GEN_792 = io_sfence_bits_rs2 & _GEN_788; // @[TLB.scala 388:40]
  assign _T_1032 = _sector_hits_T_45[26:18] == 9'h0; // @[TLB.scala 134:61]
  assign _GEN_813 = sectored_entries_0_7_data_0[13] ? _GEN_543 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_814 = sectored_entries_0_7_data_1[13] ? _GEN_544 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_815 = sectored_entries_0_7_data_2[13] ? _GEN_545 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_816 = sectored_entries_0_7_data_3[13] ? _GEN_546 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_817 = io_sfence_bits_rs2 & _GEN_813; // @[TLB.scala 388:40]
  assign _GEN_818 = io_sfence_bits_rs2 & _GEN_814; // @[TLB.scala 388:40]
  assign _GEN_819 = io_sfence_bits_rs2 & _GEN_815; // @[TLB.scala 388:40]
  assign _GEN_820 = io_sfence_bits_rs2 & _GEN_816; // @[TLB.scala 388:40]
  assign _GEN_826 = superpage_entries_0_data_0[13] ? _GEN_459 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_827 = io_sfence_bits_rs2 & _GEN_826; // @[TLB.scala 388:40]
  assign _GEN_830 = superpage_entries_1_data_0[13] ? _GEN_463 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_831 = io_sfence_bits_rs2 & _GEN_830; // @[TLB.scala 388:40]
  assign _GEN_834 = superpage_entries_2_data_0[13] ? _GEN_467 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_835 = io_sfence_bits_rs2 & _GEN_834; // @[TLB.scala 388:40]
  assign _GEN_838 = superpage_entries_3_data_0[13] ? _GEN_471 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_839 = io_sfence_bits_rs2 & _GEN_838; // @[TLB.scala 388:40]
  assign _GEN_842 = special_entry_data_0[13] ? _GEN_455 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_843 = io_sfence_bits_rs2 & _GEN_842; // @[TLB.scala 388:40]
  assign _T_1326 = multipleHits | reset; // @[TLB.scala 392:24]
  assign io_req_ready = state == 2'h0; // @[TLB.scala 341:16]
  assign io_resp_miss = _io_resp_miss_T | multipleHits; // @[TLB.scala 354:16]
  assign io_resp_paddr = {ppn,mpu_physaddr_lo}; // @[TLB.scala 355:17]
  assign io_resp_pf_ld = _io_resp_pf_ld_T | _io_resp_pf_ld_T_2; // @[TLB.scala 342:17]
  assign io_resp_pf_st = _io_resp_pf_st_T | _io_resp_pf_st_T_2; // @[TLB.scala 343:17]
  assign io_resp_ae_ld = |_io_resp_ae_ld_T; // @[TLB.scala 345:17]
  assign io_resp_ae_st = |_io_resp_ae_st_T; // @[TLB.scala 346:17]
  assign io_resp_ma_ld = |_io_resp_ma_ld_T; // @[TLB.scala 348:17]
  assign io_resp_ma_st = |_io_resp_ma_st_T; // @[TLB.scala 349:17]
  assign io_resp_cacheable = |_io_resp_cacheable_T; // @[TLB.scala 351:21]
  assign io_ptw_req_valid = state == 2'h1; // @[TLB.scala 357:20]
  assign io_ptw_req_bits_bits_addr = r_refill_tag; // @[TLB.scala 359:29]
  assign mpu_ppn_barrier_io_x_ppn = special_entry_data_0[34:15]; // @[package.scala 266:18]
  assign mpu_ppn_barrier_io_x_u = special_entry_data_0[14]; // @[package.scala 266:18]
  assign mpu_ppn_barrier_io_x_ae = special_entry_data_0[12]; // @[package.scala 266:18]
  assign mpu_ppn_barrier_io_x_sw = special_entry_data_0[11]; // @[package.scala 266:18]
  assign mpu_ppn_barrier_io_x_sx = special_entry_data_0[10]; // @[package.scala 266:18]
  assign mpu_ppn_barrier_io_x_sr = special_entry_data_0[9]; // @[package.scala 266:18]
  assign mpu_ppn_barrier_io_x_pw = special_entry_data_0[8]; // @[package.scala 266:18]
  assign mpu_ppn_barrier_io_x_px = special_entry_data_0[7]; // @[package.scala 266:18]
  assign mpu_ppn_barrier_io_x_pr = special_entry_data_0[6]; // @[package.scala 266:18]
  assign mpu_ppn_barrier_io_x_ppp = special_entry_data_0[5]; // @[package.scala 266:18]
  assign mpu_ppn_barrier_io_x_pal = special_entry_data_0[4]; // @[package.scala 266:18]
  assign mpu_ppn_barrier_io_x_paa = special_entry_data_0[3]; // @[package.scala 266:18]
  assign mpu_ppn_barrier_io_x_eff = special_entry_data_0[2]; // @[package.scala 266:18]
  assign mpu_ppn_barrier_io_x_c = special_entry_data_0[1]; // @[package.scala 266:18]
  assign pmp_io_prv = mpu_priv[1:0]; // @[TLB.scala 196:14]
  assign pmp_io_pmp_0_cfg_l = io_ptw_pmp_0_cfg_l; // @[TLB.scala 195:14]
  assign pmp_io_pmp_0_cfg_a = io_ptw_pmp_0_cfg_a; // @[TLB.scala 195:14]
  assign pmp_io_pmp_0_cfg_x = io_ptw_pmp_0_cfg_x; // @[TLB.scala 195:14]
  assign pmp_io_pmp_0_cfg_w = io_ptw_pmp_0_cfg_w; // @[TLB.scala 195:14]
  assign pmp_io_pmp_0_cfg_r = io_ptw_pmp_0_cfg_r; // @[TLB.scala 195:14]
  assign pmp_io_pmp_0_addr = io_ptw_pmp_0_addr; // @[TLB.scala 195:14]
  assign pmp_io_pmp_0_mask = io_ptw_pmp_0_mask; // @[TLB.scala 195:14]
  assign pmp_io_pmp_1_cfg_l = io_ptw_pmp_1_cfg_l; // @[TLB.scala 195:14]
  assign pmp_io_pmp_1_cfg_a = io_ptw_pmp_1_cfg_a; // @[TLB.scala 195:14]
  assign pmp_io_pmp_1_cfg_x = io_ptw_pmp_1_cfg_x; // @[TLB.scala 195:14]
  assign pmp_io_pmp_1_cfg_w = io_ptw_pmp_1_cfg_w; // @[TLB.scala 195:14]
  assign pmp_io_pmp_1_cfg_r = io_ptw_pmp_1_cfg_r; // @[TLB.scala 195:14]
  assign pmp_io_pmp_1_addr = io_ptw_pmp_1_addr; // @[TLB.scala 195:14]
  assign pmp_io_pmp_1_mask = io_ptw_pmp_1_mask; // @[TLB.scala 195:14]
  assign pmp_io_pmp_2_cfg_l = io_ptw_pmp_2_cfg_l; // @[TLB.scala 195:14]
  assign pmp_io_pmp_2_cfg_a = io_ptw_pmp_2_cfg_a; // @[TLB.scala 195:14]
  assign pmp_io_pmp_2_cfg_x = io_ptw_pmp_2_cfg_x; // @[TLB.scala 195:14]
  assign pmp_io_pmp_2_cfg_w = io_ptw_pmp_2_cfg_w; // @[TLB.scala 195:14]
  assign pmp_io_pmp_2_cfg_r = io_ptw_pmp_2_cfg_r; // @[TLB.scala 195:14]
  assign pmp_io_pmp_2_addr = io_ptw_pmp_2_addr; // @[TLB.scala 195:14]
  assign pmp_io_pmp_2_mask = io_ptw_pmp_2_mask; // @[TLB.scala 195:14]
  assign pmp_io_pmp_3_cfg_l = io_ptw_pmp_3_cfg_l; // @[TLB.scala 195:14]
  assign pmp_io_pmp_3_cfg_a = io_ptw_pmp_3_cfg_a; // @[TLB.scala 195:14]
  assign pmp_io_pmp_3_cfg_x = io_ptw_pmp_3_cfg_x; // @[TLB.scala 195:14]
  assign pmp_io_pmp_3_cfg_w = io_ptw_pmp_3_cfg_w; // @[TLB.scala 195:14]
  assign pmp_io_pmp_3_cfg_r = io_ptw_pmp_3_cfg_r; // @[TLB.scala 195:14]
  assign pmp_io_pmp_3_addr = io_ptw_pmp_3_addr; // @[TLB.scala 195:14]
  assign pmp_io_pmp_3_mask = io_ptw_pmp_3_mask; // @[TLB.scala 195:14]
  assign pmp_io_pmp_4_cfg_l = io_ptw_pmp_4_cfg_l; // @[TLB.scala 195:14]
  assign pmp_io_pmp_4_cfg_a = io_ptw_pmp_4_cfg_a; // @[TLB.scala 195:14]
  assign pmp_io_pmp_4_cfg_x = io_ptw_pmp_4_cfg_x; // @[TLB.scala 195:14]
  assign pmp_io_pmp_4_cfg_w = io_ptw_pmp_4_cfg_w; // @[TLB.scala 195:14]
  assign pmp_io_pmp_4_cfg_r = io_ptw_pmp_4_cfg_r; // @[TLB.scala 195:14]
  assign pmp_io_pmp_4_addr = io_ptw_pmp_4_addr; // @[TLB.scala 195:14]
  assign pmp_io_pmp_4_mask = io_ptw_pmp_4_mask; // @[TLB.scala 195:14]
  assign pmp_io_pmp_5_cfg_l = io_ptw_pmp_5_cfg_l; // @[TLB.scala 195:14]
  assign pmp_io_pmp_5_cfg_a = io_ptw_pmp_5_cfg_a; // @[TLB.scala 195:14]
  assign pmp_io_pmp_5_cfg_x = io_ptw_pmp_5_cfg_x; // @[TLB.scala 195:14]
  assign pmp_io_pmp_5_cfg_w = io_ptw_pmp_5_cfg_w; // @[TLB.scala 195:14]
  assign pmp_io_pmp_5_cfg_r = io_ptw_pmp_5_cfg_r; // @[TLB.scala 195:14]
  assign pmp_io_pmp_5_addr = io_ptw_pmp_5_addr; // @[TLB.scala 195:14]
  assign pmp_io_pmp_5_mask = io_ptw_pmp_5_mask; // @[TLB.scala 195:14]
  assign pmp_io_pmp_6_cfg_l = io_ptw_pmp_6_cfg_l; // @[TLB.scala 195:14]
  assign pmp_io_pmp_6_cfg_a = io_ptw_pmp_6_cfg_a; // @[TLB.scala 195:14]
  assign pmp_io_pmp_6_cfg_x = io_ptw_pmp_6_cfg_x; // @[TLB.scala 195:14]
  assign pmp_io_pmp_6_cfg_w = io_ptw_pmp_6_cfg_w; // @[TLB.scala 195:14]
  assign pmp_io_pmp_6_cfg_r = io_ptw_pmp_6_cfg_r; // @[TLB.scala 195:14]
  assign pmp_io_pmp_6_addr = io_ptw_pmp_6_addr; // @[TLB.scala 195:14]
  assign pmp_io_pmp_6_mask = io_ptw_pmp_6_mask; // @[TLB.scala 195:14]
  assign pmp_io_pmp_7_cfg_l = io_ptw_pmp_7_cfg_l; // @[TLB.scala 195:14]
  assign pmp_io_pmp_7_cfg_a = io_ptw_pmp_7_cfg_a; // @[TLB.scala 195:14]
  assign pmp_io_pmp_7_cfg_x = io_ptw_pmp_7_cfg_x; // @[TLB.scala 195:14]
  assign pmp_io_pmp_7_cfg_w = io_ptw_pmp_7_cfg_w; // @[TLB.scala 195:14]
  assign pmp_io_pmp_7_cfg_r = io_ptw_pmp_7_cfg_r; // @[TLB.scala 195:14]
  assign pmp_io_pmp_7_addr = io_ptw_pmp_7_addr; // @[TLB.scala 195:14]
  assign pmp_io_pmp_7_mask = io_ptw_pmp_7_mask; // @[TLB.scala 195:14]
  assign pmp_io_addr = mpu_physaddr[31:0]; // @[TLB.scala 193:15]
  assign pmp_io_size = io_req_bits_size; // @[TLB.scala 194:15]
  assign entries_barrier_io_x_ppn = _GEN_556[34:15]; // @[package.scala 266:18]
  assign entries_barrier_io_x_u = _GEN_556[14]; // @[package.scala 266:18]
  assign entries_barrier_io_x_ae = _GEN_556[12]; // @[package.scala 266:18]
  assign entries_barrier_io_x_sw = _GEN_556[11]; // @[package.scala 266:18]
  assign entries_barrier_io_x_sx = _GEN_556[10]; // @[package.scala 266:18]
  assign entries_barrier_io_x_sr = _GEN_556[9]; // @[package.scala 266:18]
  assign entries_barrier_io_x_pw = _GEN_556[8]; // @[package.scala 266:18]
  assign entries_barrier_io_x_px = _GEN_556[7]; // @[package.scala 266:18]
  assign entries_barrier_io_x_pr = _GEN_556[6]; // @[package.scala 266:18]
  assign entries_barrier_io_x_ppp = _GEN_556[5]; // @[package.scala 266:18]
  assign entries_barrier_io_x_pal = _GEN_556[4]; // @[package.scala 266:18]
  assign entries_barrier_io_x_paa = _GEN_556[3]; // @[package.scala 266:18]
  assign entries_barrier_io_x_eff = _GEN_556[2]; // @[package.scala 266:18]
  assign entries_barrier_io_x_c = _GEN_556[1]; // @[package.scala 266:18]
  assign entries_barrier_1_io_x_ppn = _GEN_560[34:15]; // @[package.scala 266:18]
  assign entries_barrier_1_io_x_u = _GEN_560[14]; // @[package.scala 266:18]
  assign entries_barrier_1_io_x_ae = _GEN_560[12]; // @[package.scala 266:18]
  assign entries_barrier_1_io_x_sw = _GEN_560[11]; // @[package.scala 266:18]
  assign entries_barrier_1_io_x_sx = _GEN_560[10]; // @[package.scala 266:18]
  assign entries_barrier_1_io_x_sr = _GEN_560[9]; // @[package.scala 266:18]
  assign entries_barrier_1_io_x_pw = _GEN_560[8]; // @[package.scala 266:18]
  assign entries_barrier_1_io_x_px = _GEN_560[7]; // @[package.scala 266:18]
  assign entries_barrier_1_io_x_pr = _GEN_560[6]; // @[package.scala 266:18]
  assign entries_barrier_1_io_x_ppp = _GEN_560[5]; // @[package.scala 266:18]
  assign entries_barrier_1_io_x_pal = _GEN_560[4]; // @[package.scala 266:18]
  assign entries_barrier_1_io_x_paa = _GEN_560[3]; // @[package.scala 266:18]
  assign entries_barrier_1_io_x_eff = _GEN_560[2]; // @[package.scala 266:18]
  assign entries_barrier_1_io_x_c = _GEN_560[1]; // @[package.scala 266:18]
  assign entries_barrier_2_io_x_ppn = _GEN_564[34:15]; // @[package.scala 266:18]
  assign entries_barrier_2_io_x_u = _GEN_564[14]; // @[package.scala 266:18]
  assign entries_barrier_2_io_x_ae = _GEN_564[12]; // @[package.scala 266:18]
  assign entries_barrier_2_io_x_sw = _GEN_564[11]; // @[package.scala 266:18]
  assign entries_barrier_2_io_x_sx = _GEN_564[10]; // @[package.scala 266:18]
  assign entries_barrier_2_io_x_sr = _GEN_564[9]; // @[package.scala 266:18]
  assign entries_barrier_2_io_x_pw = _GEN_564[8]; // @[package.scala 266:18]
  assign entries_barrier_2_io_x_px = _GEN_564[7]; // @[package.scala 266:18]
  assign entries_barrier_2_io_x_pr = _GEN_564[6]; // @[package.scala 266:18]
  assign entries_barrier_2_io_x_ppp = _GEN_564[5]; // @[package.scala 266:18]
  assign entries_barrier_2_io_x_pal = _GEN_564[4]; // @[package.scala 266:18]
  assign entries_barrier_2_io_x_paa = _GEN_564[3]; // @[package.scala 266:18]
  assign entries_barrier_2_io_x_eff = _GEN_564[2]; // @[package.scala 266:18]
  assign entries_barrier_2_io_x_c = _GEN_564[1]; // @[package.scala 266:18]
  assign entries_barrier_3_io_x_ppn = _GEN_568[34:15]; // @[package.scala 266:18]
  assign entries_barrier_3_io_x_u = _GEN_568[14]; // @[package.scala 266:18]
  assign entries_barrier_3_io_x_ae = _GEN_568[12]; // @[package.scala 266:18]
  assign entries_barrier_3_io_x_sw = _GEN_568[11]; // @[package.scala 266:18]
  assign entries_barrier_3_io_x_sx = _GEN_568[10]; // @[package.scala 266:18]
  assign entries_barrier_3_io_x_sr = _GEN_568[9]; // @[package.scala 266:18]
  assign entries_barrier_3_io_x_pw = _GEN_568[8]; // @[package.scala 266:18]
  assign entries_barrier_3_io_x_px = _GEN_568[7]; // @[package.scala 266:18]
  assign entries_barrier_3_io_x_pr = _GEN_568[6]; // @[package.scala 266:18]
  assign entries_barrier_3_io_x_ppp = _GEN_568[5]; // @[package.scala 266:18]
  assign entries_barrier_3_io_x_pal = _GEN_568[4]; // @[package.scala 266:18]
  assign entries_barrier_3_io_x_paa = _GEN_568[3]; // @[package.scala 266:18]
  assign entries_barrier_3_io_x_eff = _GEN_568[2]; // @[package.scala 266:18]
  assign entries_barrier_3_io_x_c = _GEN_568[1]; // @[package.scala 266:18]
  assign entries_barrier_4_io_x_ppn = _GEN_572[34:15]; // @[package.scala 266:18]
  assign entries_barrier_4_io_x_u = _GEN_572[14]; // @[package.scala 266:18]
  assign entries_barrier_4_io_x_ae = _GEN_572[12]; // @[package.scala 266:18]
  assign entries_barrier_4_io_x_sw = _GEN_572[11]; // @[package.scala 266:18]
  assign entries_barrier_4_io_x_sx = _GEN_572[10]; // @[package.scala 266:18]
  assign entries_barrier_4_io_x_sr = _GEN_572[9]; // @[package.scala 266:18]
  assign entries_barrier_4_io_x_pw = _GEN_572[8]; // @[package.scala 266:18]
  assign entries_barrier_4_io_x_px = _GEN_572[7]; // @[package.scala 266:18]
  assign entries_barrier_4_io_x_pr = _GEN_572[6]; // @[package.scala 266:18]
  assign entries_barrier_4_io_x_ppp = _GEN_572[5]; // @[package.scala 266:18]
  assign entries_barrier_4_io_x_pal = _GEN_572[4]; // @[package.scala 266:18]
  assign entries_barrier_4_io_x_paa = _GEN_572[3]; // @[package.scala 266:18]
  assign entries_barrier_4_io_x_eff = _GEN_572[2]; // @[package.scala 266:18]
  assign entries_barrier_4_io_x_c = _GEN_572[1]; // @[package.scala 266:18]
  assign entries_barrier_5_io_x_ppn = _GEN_576[34:15]; // @[package.scala 266:18]
  assign entries_barrier_5_io_x_u = _GEN_576[14]; // @[package.scala 266:18]
  assign entries_barrier_5_io_x_ae = _GEN_576[12]; // @[package.scala 266:18]
  assign entries_barrier_5_io_x_sw = _GEN_576[11]; // @[package.scala 266:18]
  assign entries_barrier_5_io_x_sx = _GEN_576[10]; // @[package.scala 266:18]
  assign entries_barrier_5_io_x_sr = _GEN_576[9]; // @[package.scala 266:18]
  assign entries_barrier_5_io_x_pw = _GEN_576[8]; // @[package.scala 266:18]
  assign entries_barrier_5_io_x_px = _GEN_576[7]; // @[package.scala 266:18]
  assign entries_barrier_5_io_x_pr = _GEN_576[6]; // @[package.scala 266:18]
  assign entries_barrier_5_io_x_ppp = _GEN_576[5]; // @[package.scala 266:18]
  assign entries_barrier_5_io_x_pal = _GEN_576[4]; // @[package.scala 266:18]
  assign entries_barrier_5_io_x_paa = _GEN_576[3]; // @[package.scala 266:18]
  assign entries_barrier_5_io_x_eff = _GEN_576[2]; // @[package.scala 266:18]
  assign entries_barrier_5_io_x_c = _GEN_576[1]; // @[package.scala 266:18]
  assign entries_barrier_6_io_x_ppn = _GEN_580[34:15]; // @[package.scala 266:18]
  assign entries_barrier_6_io_x_u = _GEN_580[14]; // @[package.scala 266:18]
  assign entries_barrier_6_io_x_ae = _GEN_580[12]; // @[package.scala 266:18]
  assign entries_barrier_6_io_x_sw = _GEN_580[11]; // @[package.scala 266:18]
  assign entries_barrier_6_io_x_sx = _GEN_580[10]; // @[package.scala 266:18]
  assign entries_barrier_6_io_x_sr = _GEN_580[9]; // @[package.scala 266:18]
  assign entries_barrier_6_io_x_pw = _GEN_580[8]; // @[package.scala 266:18]
  assign entries_barrier_6_io_x_px = _GEN_580[7]; // @[package.scala 266:18]
  assign entries_barrier_6_io_x_pr = _GEN_580[6]; // @[package.scala 266:18]
  assign entries_barrier_6_io_x_ppp = _GEN_580[5]; // @[package.scala 266:18]
  assign entries_barrier_6_io_x_pal = _GEN_580[4]; // @[package.scala 266:18]
  assign entries_barrier_6_io_x_paa = _GEN_580[3]; // @[package.scala 266:18]
  assign entries_barrier_6_io_x_eff = _GEN_580[2]; // @[package.scala 266:18]
  assign entries_barrier_6_io_x_c = _GEN_580[1]; // @[package.scala 266:18]
  assign entries_barrier_7_io_x_ppn = _GEN_584[34:15]; // @[package.scala 266:18]
  assign entries_barrier_7_io_x_u = _GEN_584[14]; // @[package.scala 266:18]
  assign entries_barrier_7_io_x_ae = _GEN_584[12]; // @[package.scala 266:18]
  assign entries_barrier_7_io_x_sw = _GEN_584[11]; // @[package.scala 266:18]
  assign entries_barrier_7_io_x_sx = _GEN_584[10]; // @[package.scala 266:18]
  assign entries_barrier_7_io_x_sr = _GEN_584[9]; // @[package.scala 266:18]
  assign entries_barrier_7_io_x_pw = _GEN_584[8]; // @[package.scala 266:18]
  assign entries_barrier_7_io_x_px = _GEN_584[7]; // @[package.scala 266:18]
  assign entries_barrier_7_io_x_pr = _GEN_584[6]; // @[package.scala 266:18]
  assign entries_barrier_7_io_x_ppp = _GEN_584[5]; // @[package.scala 266:18]
  assign entries_barrier_7_io_x_pal = _GEN_584[4]; // @[package.scala 266:18]
  assign entries_barrier_7_io_x_paa = _GEN_584[3]; // @[package.scala 266:18]
  assign entries_barrier_7_io_x_eff = _GEN_584[2]; // @[package.scala 266:18]
  assign entries_barrier_7_io_x_c = _GEN_584[1]; // @[package.scala 266:18]
  assign entries_barrier_8_io_x_ppn = superpage_entries_0_data_0[34:15]; // @[package.scala 266:18]
  assign entries_barrier_8_io_x_u = superpage_entries_0_data_0[14]; // @[package.scala 266:18]
  assign entries_barrier_8_io_x_ae = superpage_entries_0_data_0[12]; // @[package.scala 266:18]
  assign entries_barrier_8_io_x_sw = superpage_entries_0_data_0[11]; // @[package.scala 266:18]
  assign entries_barrier_8_io_x_sx = superpage_entries_0_data_0[10]; // @[package.scala 266:18]
  assign entries_barrier_8_io_x_sr = superpage_entries_0_data_0[9]; // @[package.scala 266:18]
  assign entries_barrier_8_io_x_pw = superpage_entries_0_data_0[8]; // @[package.scala 266:18]
  assign entries_barrier_8_io_x_px = superpage_entries_0_data_0[7]; // @[package.scala 266:18]
  assign entries_barrier_8_io_x_pr = superpage_entries_0_data_0[6]; // @[package.scala 266:18]
  assign entries_barrier_8_io_x_ppp = superpage_entries_0_data_0[5]; // @[package.scala 266:18]
  assign entries_barrier_8_io_x_pal = superpage_entries_0_data_0[4]; // @[package.scala 266:18]
  assign entries_barrier_8_io_x_paa = superpage_entries_0_data_0[3]; // @[package.scala 266:18]
  assign entries_barrier_8_io_x_eff = superpage_entries_0_data_0[2]; // @[package.scala 266:18]
  assign entries_barrier_8_io_x_c = superpage_entries_0_data_0[1]; // @[package.scala 266:18]
  assign entries_barrier_9_io_x_ppn = superpage_entries_1_data_0[34:15]; // @[package.scala 266:18]
  assign entries_barrier_9_io_x_u = superpage_entries_1_data_0[14]; // @[package.scala 266:18]
  assign entries_barrier_9_io_x_ae = superpage_entries_1_data_0[12]; // @[package.scala 266:18]
  assign entries_barrier_9_io_x_sw = superpage_entries_1_data_0[11]; // @[package.scala 266:18]
  assign entries_barrier_9_io_x_sx = superpage_entries_1_data_0[10]; // @[package.scala 266:18]
  assign entries_barrier_9_io_x_sr = superpage_entries_1_data_0[9]; // @[package.scala 266:18]
  assign entries_barrier_9_io_x_pw = superpage_entries_1_data_0[8]; // @[package.scala 266:18]
  assign entries_barrier_9_io_x_px = superpage_entries_1_data_0[7]; // @[package.scala 266:18]
  assign entries_barrier_9_io_x_pr = superpage_entries_1_data_0[6]; // @[package.scala 266:18]
  assign entries_barrier_9_io_x_ppp = superpage_entries_1_data_0[5]; // @[package.scala 266:18]
  assign entries_barrier_9_io_x_pal = superpage_entries_1_data_0[4]; // @[package.scala 266:18]
  assign entries_barrier_9_io_x_paa = superpage_entries_1_data_0[3]; // @[package.scala 266:18]
  assign entries_barrier_9_io_x_eff = superpage_entries_1_data_0[2]; // @[package.scala 266:18]
  assign entries_barrier_9_io_x_c = superpage_entries_1_data_0[1]; // @[package.scala 266:18]
  assign entries_barrier_10_io_x_ppn = superpage_entries_2_data_0[34:15]; // @[package.scala 266:18]
  assign entries_barrier_10_io_x_u = superpage_entries_2_data_0[14]; // @[package.scala 266:18]
  assign entries_barrier_10_io_x_ae = superpage_entries_2_data_0[12]; // @[package.scala 266:18]
  assign entries_barrier_10_io_x_sw = superpage_entries_2_data_0[11]; // @[package.scala 266:18]
  assign entries_barrier_10_io_x_sx = superpage_entries_2_data_0[10]; // @[package.scala 266:18]
  assign entries_barrier_10_io_x_sr = superpage_entries_2_data_0[9]; // @[package.scala 266:18]
  assign entries_barrier_10_io_x_pw = superpage_entries_2_data_0[8]; // @[package.scala 266:18]
  assign entries_barrier_10_io_x_px = superpage_entries_2_data_0[7]; // @[package.scala 266:18]
  assign entries_barrier_10_io_x_pr = superpage_entries_2_data_0[6]; // @[package.scala 266:18]
  assign entries_barrier_10_io_x_ppp = superpage_entries_2_data_0[5]; // @[package.scala 266:18]
  assign entries_barrier_10_io_x_pal = superpage_entries_2_data_0[4]; // @[package.scala 266:18]
  assign entries_barrier_10_io_x_paa = superpage_entries_2_data_0[3]; // @[package.scala 266:18]
  assign entries_barrier_10_io_x_eff = superpage_entries_2_data_0[2]; // @[package.scala 266:18]
  assign entries_barrier_10_io_x_c = superpage_entries_2_data_0[1]; // @[package.scala 266:18]
  assign entries_barrier_11_io_x_ppn = superpage_entries_3_data_0[34:15]; // @[package.scala 266:18]
  assign entries_barrier_11_io_x_u = superpage_entries_3_data_0[14]; // @[package.scala 266:18]
  assign entries_barrier_11_io_x_ae = superpage_entries_3_data_0[12]; // @[package.scala 266:18]
  assign entries_barrier_11_io_x_sw = superpage_entries_3_data_0[11]; // @[package.scala 266:18]
  assign entries_barrier_11_io_x_sx = superpage_entries_3_data_0[10]; // @[package.scala 266:18]
  assign entries_barrier_11_io_x_sr = superpage_entries_3_data_0[9]; // @[package.scala 266:18]
  assign entries_barrier_11_io_x_pw = superpage_entries_3_data_0[8]; // @[package.scala 266:18]
  assign entries_barrier_11_io_x_px = superpage_entries_3_data_0[7]; // @[package.scala 266:18]
  assign entries_barrier_11_io_x_pr = superpage_entries_3_data_0[6]; // @[package.scala 266:18]
  assign entries_barrier_11_io_x_ppp = superpage_entries_3_data_0[5]; // @[package.scala 266:18]
  assign entries_barrier_11_io_x_pal = superpage_entries_3_data_0[4]; // @[package.scala 266:18]
  assign entries_barrier_11_io_x_paa = superpage_entries_3_data_0[3]; // @[package.scala 266:18]
  assign entries_barrier_11_io_x_eff = superpage_entries_3_data_0[2]; // @[package.scala 266:18]
  assign entries_barrier_11_io_x_c = superpage_entries_3_data_0[1]; // @[package.scala 266:18]
  assign entries_barrier_12_io_x_ppn = special_entry_data_0[34:15]; // @[package.scala 266:18]
  assign entries_barrier_12_io_x_u = special_entry_data_0[14]; // @[package.scala 266:18]
  assign entries_barrier_12_io_x_ae = special_entry_data_0[12]; // @[package.scala 266:18]
  assign entries_barrier_12_io_x_sw = special_entry_data_0[11]; // @[package.scala 266:18]
  assign entries_barrier_12_io_x_sx = special_entry_data_0[10]; // @[package.scala 266:18]
  assign entries_barrier_12_io_x_sr = special_entry_data_0[9]; // @[package.scala 266:18]
  assign entries_barrier_12_io_x_pw = special_entry_data_0[8]; // @[package.scala 266:18]
  assign entries_barrier_12_io_x_px = special_entry_data_0[7]; // @[package.scala 266:18]
  assign entries_barrier_12_io_x_pr = special_entry_data_0[6]; // @[package.scala 266:18]
  assign entries_barrier_12_io_x_ppp = special_entry_data_0[5]; // @[package.scala 266:18]
  assign entries_barrier_12_io_x_pal = special_entry_data_0[4]; // @[package.scala 266:18]
  assign entries_barrier_12_io_x_paa = special_entry_data_0[3]; // @[package.scala 266:18]
  assign entries_barrier_12_io_x_eff = special_entry_data_0[2]; // @[package.scala 266:18]
  assign entries_barrier_12_io_x_c = special_entry_data_0[1]; // @[package.scala 266:18]
  assign TLB_cov_read_addr = TLB_state;
  assign TLB_cov_read_data = TLB_cov[TLB_cov_read_addr]; // @[Coverage map for TLB]
  assign TLB_cov_write_data = 1'h1;
  assign TLB_cov_write_addr = TLB_state;
  assign TLB_cov_write_mask = 1'h1;
  assign TLB_cov_write_en = 1'h1;
  assign mux_cond_0 = sectored_entries_0_6_data_1[0];
  assign mux_cond_1 = sectored_entries_0_7_data_1[0];
  assign mux_cond_2 = ~sectored_entries_0_2_data_0[13];
  assign mux_cond_3 = ~sectored_entries_0_7_data_1[13];
  assign mux_cond_4 = sectored_entries_0_7_data_3[0];
  assign mux_cond_5 = sectored_entries_0_4_data_0[0];
  assign mux_cond_6 = sectored_entries_0_3_data_3[0];
  assign mux_cond_7 = sectored_entries_0_2_data_3[0];
  assign mux_cond_8 = sectored_entries_0_2_data_0[0];
  assign mux_cond_9 = ~sectored_entries_0_6_data_1[13];
  assign mux_cond_10 = ~sectored_entries_0_2_data_2[13];
  assign mux_cond_11 = ~superpage_entries_0_data_0[13];
  assign mux_cond_12 = sectored_entries_0_3_data_1[0];
  assign mux_cond_13 = sectored_entries_0_4_data_3[0];
  assign mux_cond_14 = ~sectored_entries_0_3_data_3[13];
  assign mux_cond_15 = sectored_entries_0_3_data_2[0];
  assign mux_cond_16 = ~sectored_entries_0_4_data_3[13];
  assign mux_cond_17 = ~sectored_entries_0_4_data_0[13];
  assign mux_cond_18 = ~sectored_entries_0_4_data_1[13];
  assign mux_cond_19 = sectored_entries_0_6_data_0[0];
  assign mux_cond_20 = sectored_entries_0_5_data_0[0];
  assign mux_cond_21 = sectored_entries_0_6_data_2[0];
  assign mux_cond_22 = sectored_entries_0_0_data_3[0];
  assign mux_cond_23 = ~sectored_entries_0_3_data_1[13];
  assign mux_cond_24 = ~sectored_entries_0_7_data_0[13];
  assign mux_cond_25 = sectored_entries_0_7_data_0[0];
  assign mux_cond_26 = ~sectored_entries_0_7_data_3[13];
  assign mux_cond_27 = ~sectored_entries_0_0_data_3[13];
  assign mux_cond_28 = ~superpage_entries_1_data_0[13];
  assign mux_cond_29 = ~sectored_entries_0_7_data_2[13];
  assign mux_cond_30 = ~sectored_entries_0_6_data_0[13];
  assign mux_cond_31 = ~sectored_entries_0_6_data_3[13];
  assign mux_cond_32 = sectored_entries_0_2_data_2[0];
  assign mux_cond_33 = sectored_entries_0_1_data_1[0];
  assign mux_cond_34 = ~sectored_entries_0_2_data_1[13];
  assign mux_cond_35 = ~sectored_entries_0_4_data_2[13];
  assign mux_cond_36 = ~sectored_entries_0_1_data_3[13];
  assign mux_cond_37 = ~sectored_entries_0_0_data_2[13];
  assign mux_cond_38 = ~sectored_entries_0_0_data_0[13];
  assign mux_cond_39 = ~sectored_entries_0_2_data_3[13];
  assign mux_cond_40 = sectored_entries_0_7_data_2[0];
  assign mux_cond_41 = sectored_entries_0_0_data_0[0];
  assign mux_cond_42 = ~sectored_entries_0_5_data_0[13];
  assign mux_cond_43 = sectored_entries_0_4_data_1[0];
  assign mux_cond_44 = sectored_entries_0_5_data_1[0];
  assign mux_cond_45 = ~sectored_entries_0_5_data_3[13];
  assign mux_cond_46 = sectored_entries_0_1_data_0[0];
  assign mux_cond_47 = sectored_entries_0_5_data_3[0];
  assign mux_cond_48 = ~sectored_entries_0_0_data_1[13];
  assign mux_cond_49 = ~special_entry_data_0[13];
  assign mux_cond_50 = ~superpage_entries_2_data_0[13];
  assign mux_cond_51 = sectored_entries_0_0_data_2[0];
  assign mux_cond_52 = sectored_entries_0_6_data_3[0];
  assign mux_cond_53 = ~sectored_entries_0_3_data_0[13];
  assign mux_cond_54 = ~sectored_entries_0_1_data_0[13];
  assign mux_cond_55 = sectored_entries_0_1_data_2[0];
  assign mux_cond_56 = ~sectored_entries_0_5_data_2[13];
  assign mux_cond_57 = ~sectored_entries_0_6_data_2[13];
  assign mux_cond_58 = sectored_entries_0_1_data_3[0];
  assign mux_cond_59 = ~sectored_entries_0_3_data_2[13];
  assign mux_cond_60 = ~sectored_entries_0_1_data_1[13];
  assign mux_cond_61 = ~sectored_entries_0_1_data_2[13];
  assign mux_cond_62 = sectored_entries_0_3_data_0[0];
  assign mux_cond_63 = sectored_entries_0_5_data_2[0];
  assign mux_cond_64 = sectored_entries_0_0_data_1[0];
  assign mux_cond_65 = sectored_entries_0_2_data_1[0];
  assign mux_cond_66 = ~sectored_entries_0_5_data_1[13];
  assign mux_cond_67 = ~superpage_entries_3_data_0[13];
  assign mux_cond_68 = sectored_entries_0_4_data_2[0];
  assign r_sectored_hit_shl = r_sectored_hit;
  assign r_sectored_hit_pad = {19'h0,r_sectored_hit_shl};
  assign r_sectored_repl_addr_shl = {r_sectored_repl_addr, 7'h0};
  assign r_sectored_repl_addr_pad = {10'h0,r_sectored_repl_addr_shl};
  assign r_superpage_repl_addr_shl = {r_superpage_repl_addr, 18'h0};
  assign r_superpage_repl_addr_pad = r_superpage_repl_addr_shl;
  assign special_entry_valid_0_shl = {special_entry_valid_0, 7'h0};
  assign special_entry_valid_0_pad = {12'h0,special_entry_valid_0_shl};
  assign special_entry_level_shl = {special_entry_level, 18'h0};
  assign special_entry_level_pad = special_entry_level_shl;
  assign state_shl = {state, 6'h0};
  assign state_pad = {12'h0,state_shl};
  assign r_sectored_hit_addr_shl = {r_sectored_hit_addr, 12'h0};
  assign r_sectored_hit_addr_pad = {5'h0,r_sectored_hit_addr_shl};
  assign mux_cond_0_shl = {mux_cond_0, 5'h0};
  assign mux_cond_0_pad = {14'h0,mux_cond_0_shl};
  assign mux_cond_1_shl = {mux_cond_1, 11'h0};
  assign mux_cond_1_pad = {8'h0,mux_cond_1_shl};
  assign mux_cond_2_shl = {mux_cond_2, 2'h0};
  assign mux_cond_2_pad = {17'h0,mux_cond_2_shl};
  assign mux_cond_3_shl = {mux_cond_3, 12'h0};
  assign mux_cond_3_pad = {7'h0,mux_cond_3_shl};
  assign mux_cond_4_shl = {mux_cond_4, 11'h0};
  assign mux_cond_4_pad = {8'h0,mux_cond_4_shl};
  assign mux_cond_5_shl = {mux_cond_5, 1'h0};
  assign mux_cond_5_pad = {18'h0,mux_cond_5_shl};
  assign mux_cond_6_shl = {mux_cond_6, 13'h0};
  assign mux_cond_6_pad = {6'h0,mux_cond_6_shl};
  assign mux_cond_7_shl = {mux_cond_7, 6'h0};
  assign mux_cond_7_pad = {13'h0,mux_cond_7_shl};
  assign mux_cond_8_shl = {mux_cond_8, 4'h0};
  assign mux_cond_8_pad = {15'h0,mux_cond_8_shl};
  assign mux_cond_9_shl = {mux_cond_9, 17'h0};
  assign mux_cond_9_pad = {2'h0,mux_cond_9_shl};
  assign mux_cond_10_shl = {mux_cond_10, 5'h0};
  assign mux_cond_10_pad = {14'h0,mux_cond_10_shl};
  assign mux_cond_11_shl = {mux_cond_11, 9'h0};
  assign mux_cond_11_pad = {10'h0,mux_cond_11_shl};
  assign mux_cond_12_shl = {mux_cond_12, 1'h0};
  assign mux_cond_12_pad = {18'h0,mux_cond_12_shl};
  assign mux_cond_13_shl = {mux_cond_13, 9'h0};
  assign mux_cond_13_pad = {10'h0,mux_cond_13_shl};
  assign mux_cond_14_shl = {mux_cond_14, 12'h0};
  assign mux_cond_14_pad = {7'h0,mux_cond_14_shl};
  assign mux_cond_15_shl = {mux_cond_15, 7'h0};
  assign mux_cond_15_pad = {12'h0,mux_cond_15_shl};
  assign mux_cond_16_shl = {mux_cond_16, 6'h0};
  assign mux_cond_16_pad = {13'h0,mux_cond_16_shl};
  assign mux_cond_17_shl = {mux_cond_17, 7'h0};
  assign mux_cond_17_pad = {12'h0,mux_cond_17_shl};
  assign mux_cond_18_shl = {mux_cond_18, 16'h0};
  assign mux_cond_18_pad = {3'h0,mux_cond_18_shl};
  assign mux_cond_19_shl = {mux_cond_19, 8'h0};
  assign mux_cond_19_pad = {11'h0,mux_cond_19_shl};
  assign mux_cond_20_shl = {mux_cond_20, 1'h0};
  assign mux_cond_20_pad = {18'h0,mux_cond_20_shl};
  assign mux_cond_21_shl = {mux_cond_21, 5'h0};
  assign mux_cond_21_pad = {14'h0,mux_cond_21_shl};
  assign mux_cond_22_shl = {mux_cond_22, 11'h0};
  assign mux_cond_22_pad = {8'h0,mux_cond_22_shl};
  assign mux_cond_23_shl = {mux_cond_23, 2'h0};
  assign mux_cond_23_pad = {17'h0,mux_cond_23_shl};
  assign mux_cond_24_shl = {mux_cond_24, 14'h0};
  assign mux_cond_24_pad = {5'h0,mux_cond_24_shl};
  assign mux_cond_25_shl = {mux_cond_25, 3'h0};
  assign mux_cond_25_pad = {16'h0,mux_cond_25_shl};
  assign mux_cond_26_shl = {mux_cond_26, 11'h0};
  assign mux_cond_26_pad = {8'h0,mux_cond_26_shl};
  assign mux_cond_27_shl = mux_cond_27;
  assign mux_cond_27_pad = {19'h0,mux_cond_27_shl};
  assign mux_cond_28_shl = {mux_cond_28, 18'h0};
  assign mux_cond_28_pad = {1'h0,mux_cond_28_shl};
  assign mux_cond_29_shl = {mux_cond_29, 14'h0};
  assign mux_cond_29_pad = {5'h0,mux_cond_29_shl};
  assign mux_cond_30_shl = {mux_cond_30, 8'h0};
  assign mux_cond_30_pad = {11'h0,mux_cond_30_shl};
  assign mux_cond_31_shl = {mux_cond_31, 3'h0};
  assign mux_cond_31_pad = {16'h0,mux_cond_31_shl};
  assign mux_cond_32_shl = {mux_cond_32, 2'h0};
  assign mux_cond_32_pad = {17'h0,mux_cond_32_shl};
  assign mux_cond_33_shl = mux_cond_33;
  assign mux_cond_33_pad = {19'h0,mux_cond_33_shl};
  assign mux_cond_34_shl = {mux_cond_34, 7'h0};
  assign mux_cond_34_pad = {12'h0,mux_cond_34_shl};
  assign mux_cond_35_shl = {mux_cond_35, 4'h0};
  assign mux_cond_35_pad = {15'h0,mux_cond_35_shl};
  assign mux_cond_36_shl = {mux_cond_36, 3'h0};
  assign mux_cond_36_pad = {16'h0,mux_cond_36_shl};
  assign mux_cond_37_shl = {mux_cond_37, 4'h0};
  assign mux_cond_37_pad = {15'h0,mux_cond_37_shl};
  assign mux_cond_38_shl = {mux_cond_38, 12'h0};
  assign mux_cond_38_pad = {7'h0,mux_cond_38_shl};
  assign mux_cond_39_shl = {mux_cond_39, 9'h0};
  assign mux_cond_39_pad = {10'h0,mux_cond_39_shl};
  assign mux_cond_40_shl = mux_cond_40;
  assign mux_cond_40_pad = {19'h0,mux_cond_40_shl};
  assign mux_cond_41_shl = {mux_cond_41, 16'h0};
  assign mux_cond_41_pad = {3'h0,mux_cond_41_shl};
  assign mux_cond_42_shl = {mux_cond_42, 4'h0};
  assign mux_cond_42_pad = {15'h0,mux_cond_42_shl};
  assign mux_cond_43_shl = {mux_cond_43, 18'h0};
  assign mux_cond_43_pad = {1'h0,mux_cond_43_shl};
  assign mux_cond_44_shl = {mux_cond_44, 8'h0};
  assign mux_cond_44_pad = {11'h0,mux_cond_44_shl};
  assign mux_cond_45_shl = {mux_cond_45, 17'h0};
  assign mux_cond_45_pad = {2'h0,mux_cond_45_shl};
  assign mux_cond_46_shl = {mux_cond_46, 5'h0};
  assign mux_cond_46_pad = {14'h0,mux_cond_46_shl};
  assign mux_cond_47_shl = {mux_cond_47, 8'h0};
  assign mux_cond_47_pad = {11'h0,mux_cond_47_shl};
  assign mux_cond_48_shl = {mux_cond_48, 7'h0};
  assign mux_cond_48_pad = {12'h0,mux_cond_48_shl};
  assign mux_cond_49_shl = {mux_cond_49, 16'h0};
  assign mux_cond_49_pad = {3'h0,mux_cond_49_shl};
  assign mux_cond_50_shl = {mux_cond_50, 8'h0};
  assign mux_cond_50_pad = {11'h0,mux_cond_50_shl};
  assign mux_cond_51_shl = {mux_cond_51, 4'h0};
  assign mux_cond_51_pad = {15'h0,mux_cond_51_shl};
  assign mux_cond_52_shl = {mux_cond_52, 3'h0};
  assign mux_cond_52_pad = {16'h0,mux_cond_52_shl};
  assign mux_cond_53_shl = {mux_cond_53, 6'h0};
  assign mux_cond_53_pad = {13'h0,mux_cond_53_shl};
  assign mux_cond_54_shl = {mux_cond_54, 18'h0};
  assign mux_cond_54_pad = {1'h0,mux_cond_54_shl};
  assign mux_cond_55_shl = {mux_cond_55, 15'h0};
  assign mux_cond_55_pad = {4'h0,mux_cond_55_shl};
  assign mux_cond_56_shl = {mux_cond_56, 16'h0};
  assign mux_cond_56_pad = {3'h0,mux_cond_56_shl};
  assign mux_cond_57_shl = {mux_cond_57, 7'h0};
  assign mux_cond_57_pad = {12'h0,mux_cond_57_shl};
  assign mux_cond_58_shl = {mux_cond_58, 11'h0};
  assign mux_cond_58_pad = {8'h0,mux_cond_58_shl};
  assign mux_cond_59_shl = {mux_cond_59, 14'h0};
  assign mux_cond_59_pad = {5'h0,mux_cond_59_shl};
  assign mux_cond_60_shl = {mux_cond_60, 13'h0};
  assign mux_cond_60_pad = {6'h0,mux_cond_60_shl};
  assign mux_cond_61_shl = {mux_cond_61, 8'h0};
  assign mux_cond_61_pad = {11'h0,mux_cond_61_shl};
  assign mux_cond_62_shl = {mux_cond_62, 7'h0};
  assign mux_cond_62_pad = {12'h0,mux_cond_62_shl};
  assign mux_cond_63_shl = {mux_cond_63, 6'h0};
  assign mux_cond_63_pad = {13'h0,mux_cond_63_shl};
  assign mux_cond_64_shl = {mux_cond_64, 19'h0};
  assign mux_cond_64_pad = mux_cond_64_shl;
  assign mux_cond_65_shl = {mux_cond_65, 11'h0};
  assign mux_cond_65_pad = {8'h0,mux_cond_65_shl};
  assign mux_cond_66_shl = {mux_cond_66, 6'h0};
  assign mux_cond_66_pad = {13'h0,mux_cond_66_shl};
  assign mux_cond_67_shl = {mux_cond_67, 10'h0};
  assign mux_cond_67_pad = {9'h0,mux_cond_67_shl};
  assign mux_cond_68_shl = {mux_cond_68, 13'h0};
  assign mux_cond_68_pad = {6'h0,mux_cond_68_shl};
  assign sectored_entries_0_0_valid_3_shl = {sectored_entries_0_0_valid_3, 16'h0};
  assign sectored_entries_0_0_valid_3_pad = {3'h0,sectored_entries_0_0_valid_3_shl};
  assign sectored_entries_0_0_valid_2_shl = {sectored_entries_0_0_valid_2, 8'h0};
  assign sectored_entries_0_0_valid_2_pad = {11'h0,sectored_entries_0_0_valid_2_shl};
  assign sectored_entries_0_2_valid_0_shl = {sectored_entries_0_2_valid_0, 8'h0};
  assign sectored_entries_0_2_valid_0_pad = {11'h0,sectored_entries_0_2_valid_0_shl};
  assign sectored_entries_0_3_valid_0_shl = {sectored_entries_0_3_valid_0, 8'h0};
  assign sectored_entries_0_3_valid_0_pad = {11'h0,sectored_entries_0_3_valid_0_shl};
  assign superpage_entries_2_level_shl = superpage_entries_2_level;
  assign superpage_entries_2_level_pad = {18'h0,superpage_entries_2_level_shl};
  assign sectored_entries_0_7_valid_1_shl = sectored_entries_0_7_valid_1;
  assign sectored_entries_0_7_valid_1_pad = {19'h0,sectored_entries_0_7_valid_1_shl};
  assign sectored_entries_0_4_valid_0_shl = {sectored_entries_0_4_valid_0, 8'h0};
  assign sectored_entries_0_4_valid_0_pad = {11'h0,sectored_entries_0_4_valid_0_shl};
  assign sectored_entries_0_1_valid_3_shl = {sectored_entries_0_1_valid_3, 16'h0};
  assign sectored_entries_0_1_valid_3_pad = {3'h0,sectored_entries_0_1_valid_3_shl};
  assign sectored_entries_0_1_valid_1_shl = sectored_entries_0_1_valid_1;
  assign sectored_entries_0_1_valid_1_pad = {19'h0,sectored_entries_0_1_valid_1_shl};
  assign sectored_entries_0_2_valid_3_shl = {sectored_entries_0_2_valid_3, 16'h0};
  assign sectored_entries_0_2_valid_3_pad = {3'h0,sectored_entries_0_2_valid_3_shl};
  assign sectored_entries_0_2_valid_1_shl = sectored_entries_0_2_valid_1;
  assign sectored_entries_0_2_valid_1_pad = {19'h0,sectored_entries_0_2_valid_1_shl};
  assign superpage_entries_1_valid_0_shl = {superpage_entries_1_valid_0, 11'h0};
  assign superpage_entries_1_valid_0_pad = {8'h0,superpage_entries_1_valid_0_shl};
  assign sectored_entries_0_7_valid_0_shl = {sectored_entries_0_7_valid_0, 8'h0};
  assign sectored_entries_0_7_valid_0_pad = {11'h0,sectored_entries_0_7_valid_0_shl};
  assign superpage_entries_3_valid_0_shl = {superpage_entries_3_valid_0, 11'h0};
  assign superpage_entries_3_valid_0_pad = {8'h0,superpage_entries_3_valid_0_shl};
  assign sectored_entries_0_5_valid_3_shl = {sectored_entries_0_5_valid_3, 16'h0};
  assign sectored_entries_0_5_valid_3_pad = {3'h0,sectored_entries_0_5_valid_3_shl};
  assign sectored_entries_0_5_valid_1_shl = sectored_entries_0_5_valid_1;
  assign sectored_entries_0_5_valid_1_pad = {19'h0,sectored_entries_0_5_valid_1_shl};
  assign sectored_entries_0_4_valid_3_shl = {sectored_entries_0_4_valid_3, 16'h0};
  assign sectored_entries_0_4_valid_3_pad = {3'h0,sectored_entries_0_4_valid_3_shl};
  assign sectored_entries_0_5_valid_2_shl = {sectored_entries_0_5_valid_2, 8'h0};
  assign sectored_entries_0_5_valid_2_pad = {11'h0,sectored_entries_0_5_valid_2_shl};
  assign sectored_entries_0_1_valid_2_shl = {sectored_entries_0_1_valid_2, 8'h0};
  assign sectored_entries_0_1_valid_2_pad = {11'h0,sectored_entries_0_1_valid_2_shl};
  assign sectored_entries_0_3_valid_1_shl = sectored_entries_0_3_valid_1;
  assign sectored_entries_0_3_valid_1_pad = {19'h0,sectored_entries_0_3_valid_1_shl};
  assign sectored_entries_0_1_valid_0_shl = {sectored_entries_0_1_valid_0, 8'h0};
  assign sectored_entries_0_1_valid_0_pad = {11'h0,sectored_entries_0_1_valid_0_shl};
  assign sectored_entries_0_4_valid_2_shl = {sectored_entries_0_4_valid_2, 8'h0};
  assign sectored_entries_0_4_valid_2_pad = {11'h0,sectored_entries_0_4_valid_2_shl};
  assign sectored_entries_0_4_valid_1_shl = sectored_entries_0_4_valid_1;
  assign sectored_entries_0_4_valid_1_pad = {19'h0,sectored_entries_0_4_valid_1_shl};
  assign superpage_entries_3_level_shl = superpage_entries_3_level;
  assign superpage_entries_3_level_pad = {18'h0,superpage_entries_3_level_shl};
  assign sectored_entries_0_0_valid_1_shl = sectored_entries_0_0_valid_1;
  assign sectored_entries_0_0_valid_1_pad = {19'h0,sectored_entries_0_0_valid_1_shl};
  assign sectored_entries_0_3_valid_2_shl = {sectored_entries_0_3_valid_2, 8'h0};
  assign sectored_entries_0_3_valid_2_pad = {11'h0,sectored_entries_0_3_valid_2_shl};
  assign sectored_entries_0_6_valid_1_shl = sectored_entries_0_6_valid_1;
  assign sectored_entries_0_6_valid_1_pad = {19'h0,sectored_entries_0_6_valid_1_shl};
  assign sectored_entries_0_7_valid_3_shl = {sectored_entries_0_7_valid_3, 16'h0};
  assign sectored_entries_0_7_valid_3_pad = {3'h0,sectored_entries_0_7_valid_3_shl};
  assign sectored_entries_0_3_valid_3_shl = {sectored_entries_0_3_valid_3, 16'h0};
  assign sectored_entries_0_3_valid_3_pad = {3'h0,sectored_entries_0_3_valid_3_shl};
  assign sectored_entries_0_0_valid_0_shl = {sectored_entries_0_0_valid_0, 8'h0};
  assign sectored_entries_0_0_valid_0_pad = {11'h0,sectored_entries_0_0_valid_0_shl};
  assign superpage_entries_0_valid_0_shl = {superpage_entries_0_valid_0, 11'h0};
  assign superpage_entries_0_valid_0_pad = {8'h0,superpage_entries_0_valid_0_shl};
  assign sectored_entries_0_2_valid_2_shl = {sectored_entries_0_2_valid_2, 8'h0};
  assign sectored_entries_0_2_valid_2_pad = {11'h0,sectored_entries_0_2_valid_2_shl};
  assign sectored_entries_0_6_valid_2_shl = {sectored_entries_0_6_valid_2, 8'h0};
  assign sectored_entries_0_6_valid_2_pad = {11'h0,sectored_entries_0_6_valid_2_shl};
  assign superpage_entries_2_valid_0_shl = {superpage_entries_2_valid_0, 11'h0};
  assign superpage_entries_2_valid_0_pad = {8'h0,superpage_entries_2_valid_0_shl};
  assign sectored_entries_0_6_valid_3_shl = {sectored_entries_0_6_valid_3, 16'h0};
  assign sectored_entries_0_6_valid_3_pad = {3'h0,sectored_entries_0_6_valid_3_shl};
  assign sectored_entries_0_6_valid_0_shl = {sectored_entries_0_6_valid_0, 8'h0};
  assign sectored_entries_0_6_valid_0_pad = {11'h0,sectored_entries_0_6_valid_0_shl};
  assign sectored_entries_0_7_valid_2_shl = {sectored_entries_0_7_valid_2, 8'h0};
  assign sectored_entries_0_7_valid_2_pad = {11'h0,sectored_entries_0_7_valid_2_shl};
  assign superpage_entries_0_level_shl = superpage_entries_0_level;
  assign superpage_entries_0_level_pad = {18'h0,superpage_entries_0_level_shl};
  assign superpage_entries_1_level_shl = superpage_entries_1_level;
  assign superpage_entries_1_level_pad = {18'h0,superpage_entries_1_level_shl};
  assign sectored_entries_0_5_valid_0_shl = {sectored_entries_0_5_valid_0, 8'h0};
  assign sectored_entries_0_5_valid_0_pad = {11'h0,sectored_entries_0_5_valid_0_shl};
  assign TLB_xor64 = r_sectored_repl_addr_pad ^ r_superpage_repl_addr_pad;
  assign TLB_xor31 = r_sectored_hit_pad ^ TLB_xor64;
  assign TLB_xor65 = special_entry_valid_0_pad ^ special_entry_level_pad;
  assign TLB_xor66 = state_pad ^ r_sectored_hit_addr_pad;
  assign TLB_xor32 = TLB_xor65 ^ TLB_xor66;
  assign TLB_xor15 = TLB_xor31 ^ TLB_xor32;
  assign TLB_xor68 = mux_cond_1_pad ^ mux_cond_2_pad;
  assign TLB_xor33 = mux_cond_0_pad ^ TLB_xor68;
  assign TLB_xor69 = mux_cond_3_pad ^ mux_cond_4_pad;
  assign TLB_xor70 = mux_cond_5_pad ^ mux_cond_6_pad;
  assign TLB_xor34 = TLB_xor69 ^ TLB_xor70;
  assign TLB_xor16 = TLB_xor33 ^ TLB_xor34;
  assign TLB_xor7 = TLB_xor15 ^ TLB_xor16;
  assign TLB_xor72 = mux_cond_8_pad ^ mux_cond_9_pad;
  assign TLB_xor35 = mux_cond_7_pad ^ TLB_xor72;
  assign TLB_xor73 = mux_cond_10_pad ^ mux_cond_11_pad;
  assign TLB_xor74 = mux_cond_12_pad ^ mux_cond_13_pad;
  assign TLB_xor36 = TLB_xor73 ^ TLB_xor74;
  assign TLB_xor17 = TLB_xor35 ^ TLB_xor36;
  assign TLB_xor75 = mux_cond_14_pad ^ mux_cond_15_pad;
  assign TLB_xor76 = mux_cond_16_pad ^ mux_cond_17_pad;
  assign TLB_xor37 = TLB_xor75 ^ TLB_xor76;
  assign TLB_xor77 = mux_cond_18_pad ^ mux_cond_19_pad;
  assign TLB_xor78 = mux_cond_20_pad ^ mux_cond_21_pad;
  assign TLB_xor38 = TLB_xor77 ^ TLB_xor78;
  assign TLB_xor18 = TLB_xor37 ^ TLB_xor38;
  assign TLB_xor8 = TLB_xor17 ^ TLB_xor18;
  assign TLB_xor3 = TLB_xor7 ^ TLB_xor8;
  assign TLB_xor80 = mux_cond_23_pad ^ mux_cond_24_pad;
  assign TLB_xor39 = mux_cond_22_pad ^ TLB_xor80;
  assign TLB_xor81 = mux_cond_25_pad ^ mux_cond_26_pad;
  assign TLB_xor82 = mux_cond_27_pad ^ mux_cond_28_pad;
  assign TLB_xor40 = TLB_xor81 ^ TLB_xor82;
  assign TLB_xor19 = TLB_xor39 ^ TLB_xor40;
  assign TLB_xor84 = mux_cond_30_pad ^ mux_cond_31_pad;
  assign TLB_xor41 = mux_cond_29_pad ^ TLB_xor84;
  assign TLB_xor85 = mux_cond_32_pad ^ mux_cond_33_pad;
  assign TLB_xor86 = mux_cond_34_pad ^ mux_cond_35_pad;
  assign TLB_xor42 = TLB_xor85 ^ TLB_xor86;
  assign TLB_xor20 = TLB_xor41 ^ TLB_xor42;
  assign TLB_xor9 = TLB_xor19 ^ TLB_xor20;
  assign TLB_xor88 = mux_cond_37_pad ^ mux_cond_38_pad;
  assign TLB_xor43 = mux_cond_36_pad ^ TLB_xor88;
  assign TLB_xor89 = mux_cond_39_pad ^ mux_cond_40_pad;
  assign TLB_xor90 = mux_cond_41_pad ^ mux_cond_42_pad;
  assign TLB_xor44 = TLB_xor89 ^ TLB_xor90;
  assign TLB_xor21 = TLB_xor43 ^ TLB_xor44;
  assign TLB_xor91 = mux_cond_43_pad ^ mux_cond_44_pad;
  assign TLB_xor92 = mux_cond_45_pad ^ mux_cond_46_pad;
  assign TLB_xor45 = TLB_xor91 ^ TLB_xor92;
  assign TLB_xor93 = mux_cond_47_pad ^ mux_cond_48_pad;
  assign TLB_xor94 = mux_cond_49_pad ^ mux_cond_50_pad;
  assign TLB_xor46 = TLB_xor93 ^ TLB_xor94;
  assign TLB_xor22 = TLB_xor45 ^ TLB_xor46;
  assign TLB_xor10 = TLB_xor21 ^ TLB_xor22;
  assign TLB_xor4 = TLB_xor9 ^ TLB_xor10;
  assign TLB_xor1 = TLB_xor3 ^ TLB_xor4;
  assign TLB_xor96 = mux_cond_52_pad ^ mux_cond_53_pad;
  assign TLB_xor47 = mux_cond_51_pad ^ TLB_xor96;
  assign TLB_xor97 = mux_cond_54_pad ^ mux_cond_55_pad;
  assign TLB_xor98 = mux_cond_56_pad ^ mux_cond_57_pad;
  assign TLB_xor48 = TLB_xor97 ^ TLB_xor98;
  assign TLB_xor23 = TLB_xor47 ^ TLB_xor48;
  assign TLB_xor100 = mux_cond_59_pad ^ mux_cond_60_pad;
  assign TLB_xor49 = mux_cond_58_pad ^ TLB_xor100;
  assign TLB_xor101 = mux_cond_61_pad ^ mux_cond_62_pad;
  assign TLB_xor102 = mux_cond_63_pad ^ mux_cond_64_pad;
  assign TLB_xor50 = TLB_xor101 ^ TLB_xor102;
  assign TLB_xor24 = TLB_xor49 ^ TLB_xor50;
  assign TLB_xor11 = TLB_xor23 ^ TLB_xor24;
  assign TLB_xor104 = mux_cond_66_pad ^ mux_cond_67_pad;
  assign TLB_xor51 = mux_cond_65_pad ^ TLB_xor104;
  assign TLB_xor105 = mux_cond_68_pad ^ sectored_entries_0_0_valid_3_pad;
  assign TLB_xor106 = sectored_entries_0_0_valid_2_pad ^ sectored_entries_0_2_valid_0_pad;
  assign TLB_xor52 = TLB_xor105 ^ TLB_xor106;
  assign TLB_xor25 = TLB_xor51 ^ TLB_xor52;
  assign TLB_xor107 = sectored_entries_0_3_valid_0_pad ^ superpage_entries_2_level_pad;
  assign TLB_xor108 = sectored_entries_0_7_valid_1_pad ^ sectored_entries_0_4_valid_0_pad;
  assign TLB_xor53 = TLB_xor107 ^ TLB_xor108;
  assign TLB_xor109 = sectored_entries_0_1_valid_3_pad ^ sectored_entries_0_1_valid_1_pad;
  assign TLB_xor110 = sectored_entries_0_2_valid_3_pad ^ sectored_entries_0_2_valid_1_pad;
  assign TLB_xor54 = TLB_xor109 ^ TLB_xor110;
  assign TLB_xor26 = TLB_xor53 ^ TLB_xor54;
  assign TLB_xor12 = TLB_xor25 ^ TLB_xor26;
  assign TLB_xor5 = TLB_xor11 ^ TLB_xor12;
  assign TLB_xor112 = sectored_entries_0_7_valid_0_pad ^ superpage_entries_3_valid_0_pad;
  assign TLB_xor55 = superpage_entries_1_valid_0_pad ^ TLB_xor112;
  assign TLB_xor113 = sectored_entries_0_5_valid_3_pad ^ sectored_entries_0_5_valid_1_pad;
  assign TLB_xor114 = sectored_entries_0_4_valid_3_pad ^ sectored_entries_0_5_valid_2_pad;
  assign TLB_xor56 = TLB_xor113 ^ TLB_xor114;
  assign TLB_xor27 = TLB_xor55 ^ TLB_xor56;
  assign TLB_xor116 = sectored_entries_0_3_valid_1_pad ^ sectored_entries_0_1_valid_0_pad;
  assign TLB_xor57 = sectored_entries_0_1_valid_2_pad ^ TLB_xor116;
  assign TLB_xor117 = sectored_entries_0_4_valid_2_pad ^ sectored_entries_0_4_valid_1_pad;
  assign TLB_xor118 = superpage_entries_3_level_pad ^ sectored_entries_0_0_valid_1_pad;
  assign TLB_xor58 = TLB_xor117 ^ TLB_xor118;
  assign TLB_xor28 = TLB_xor57 ^ TLB_xor58;
  assign TLB_xor13 = TLB_xor27 ^ TLB_xor28;
  assign TLB_xor120 = sectored_entries_0_6_valid_1_pad ^ sectored_entries_0_7_valid_3_pad;
  assign TLB_xor59 = sectored_entries_0_3_valid_2_pad ^ TLB_xor120;
  assign TLB_xor121 = sectored_entries_0_3_valid_3_pad ^ sectored_entries_0_0_valid_0_pad;
  assign TLB_xor122 = superpage_entries_0_valid_0_pad ^ sectored_entries_0_2_valid_2_pad;
  assign TLB_xor60 = TLB_xor121 ^ TLB_xor122;
  assign TLB_xor29 = TLB_xor59 ^ TLB_xor60;
  assign TLB_xor123 = sectored_entries_0_6_valid_2_pad ^ superpage_entries_2_valid_0_pad;
  assign TLB_xor124 = sectored_entries_0_6_valid_3_pad ^ sectored_entries_0_6_valid_0_pad;
  assign TLB_xor61 = TLB_xor123 ^ TLB_xor124;
  assign TLB_xor125 = sectored_entries_0_7_valid_2_pad ^ superpage_entries_0_level_pad;
  assign TLB_xor126 = superpage_entries_1_level_pad ^ sectored_entries_0_5_valid_0_pad;
  assign TLB_xor62 = TLB_xor125 ^ TLB_xor126;
  assign TLB_xor30 = TLB_xor61 ^ TLB_xor62;
  assign TLB_xor14 = TLB_xor29 ^ TLB_xor30;
  assign TLB_xor6 = TLB_xor13 ^ TLB_xor14;
  assign TLB_xor2 = TLB_xor5 ^ TLB_xor6;
  assign TLB_xor0 = TLB_xor1 ^ TLB_xor2;
  assign mpu_ppn_barrier_sum = TLB_covSum + mpu_ppn_barrier_io_covSum;
  assign entries_barrier_10_sum = mpu_ppn_barrier_sum + entries_barrier_10_io_covSum;
  assign entries_barrier_9_sum = entries_barrier_10_sum + entries_barrier_9_io_covSum;
  assign entries_barrier_7_sum = entries_barrier_9_sum + entries_barrier_7_io_covSum;
  assign entries_barrier_sum = entries_barrier_7_sum + entries_barrier_io_covSum;
  assign entries_barrier_6_sum = entries_barrier_sum + entries_barrier_6_io_covSum;
  assign entries_barrier_12_sum = entries_barrier_6_sum + entries_barrier_12_io_covSum;
  assign entries_barrier_1_sum = entries_barrier_12_sum + entries_barrier_1_io_covSum;
  assign entries_barrier_11_sum = entries_barrier_1_sum + entries_barrier_11_io_covSum;
  assign entries_barrier_8_sum = entries_barrier_11_sum + entries_barrier_8_io_covSum;
  assign pmp_sum = entries_barrier_8_sum + pmp_io_covSum;
  assign entries_barrier_2_sum = pmp_sum + entries_barrier_2_io_covSum;
  assign entries_barrier_4_sum = entries_barrier_2_sum + entries_barrier_4_io_covSum;
  assign entries_barrier_5_sum = entries_barrier_4_sum + entries_barrier_5_io_covSum;
  assign entries_barrier_3_sum = entries_barrier_5_sum + entries_barrier_3_io_covSum;
  assign io_covSum = entries_barrier_3_sum;
  assign stopEn0 = io_sfence_valid & ~_T_51;
  assign entries_barrier_12_metaAssert_wire = entries_barrier_12_metaAssert;
  assign entries_barrier_metaAssert_wire = entries_barrier_metaAssert;
  assign entries_barrier_10_metaAssert_wire = entries_barrier_10_metaAssert;
  assign entries_barrier_5_metaAssert_wire = entries_barrier_5_metaAssert;
  assign entries_barrier_11_metaAssert_wire = entries_barrier_11_metaAssert;
  assign entries_barrier_9_metaAssert_wire = entries_barrier_9_metaAssert;
  assign entries_barrier_8_metaAssert_wire = entries_barrier_8_metaAssert;
  assign entries_barrier_1_metaAssert_wire = entries_barrier_1_metaAssert;
  assign mpu_ppn_barrier_metaAssert_wire = mpu_ppn_barrier_metaAssert;
  assign entries_barrier_4_metaAssert_wire = entries_barrier_4_metaAssert;
  assign entries_barrier_6_metaAssert_wire = entries_barrier_6_metaAssert;
  assign entries_barrier_3_metaAssert_wire = entries_barrier_3_metaAssert;
  assign pmp_metaAssert_wire = pmp_metaAssert;
  assign entries_barrier_7_metaAssert_wire = entries_barrier_7_metaAssert;
  assign entries_barrier_2_metaAssert_wire = entries_barrier_2_metaAssert;
  assign TLB_or7 = stopEn0 | entries_barrier_6_metaAssert_wire;
  assign TLB_or8 = entries_barrier_10_metaAssert_wire | entries_barrier_7_metaAssert_wire;
  assign TLB_or3 = TLB_or7 | TLB_or8;
  assign TLB_or9 = entries_barrier_4_metaAssert_wire | entries_barrier_11_metaAssert_wire;
  assign TLB_or10 = entries_barrier_8_metaAssert_wire | entries_barrier_9_metaAssert_wire;
  assign TLB_or4 = TLB_or9 | TLB_or10;
  assign TLB_or1 = TLB_or3 | TLB_or4;
  assign TLB_or11 = entries_barrier_metaAssert_wire | entries_barrier_3_metaAssert_wire;
  assign TLB_or12 = pmp_metaAssert_wire | mpu_ppn_barrier_metaAssert_wire;
  assign TLB_or5 = TLB_or11 | TLB_or12;
  assign TLB_or13 = entries_barrier_12_metaAssert_wire | entries_barrier_5_metaAssert_wire;
  assign TLB_or14 = entries_barrier_2_metaAssert_wire | entries_barrier_1_metaAssert_wire;
  assign TLB_or6 = TLB_or13 | TLB_or14;
  assign TLB_or2 = TLB_or5 | TLB_or6;
  assign TLB_or0 = TLB_or1 | TLB_or2;
  assign metaAssert = TLB_metaAssert;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sectored_entries_0_0_tag = _RAND_0[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {2{`RANDOM}};
  sectored_entries_0_0_data_0 = _RAND_1[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {2{`RANDOM}};
  sectored_entries_0_0_data_1 = _RAND_2[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {2{`RANDOM}};
  sectored_entries_0_0_data_2 = _RAND_3[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {2{`RANDOM}};
  sectored_entries_0_0_data_3 = _RAND_4[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  sectored_entries_0_0_valid_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  sectored_entries_0_0_valid_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  sectored_entries_0_0_valid_2 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  sectored_entries_0_0_valid_3 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  sectored_entries_0_1_tag = _RAND_9[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {2{`RANDOM}};
  sectored_entries_0_1_data_0 = _RAND_10[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {2{`RANDOM}};
  sectored_entries_0_1_data_1 = _RAND_11[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {2{`RANDOM}};
  sectored_entries_0_1_data_2 = _RAND_12[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {2{`RANDOM}};
  sectored_entries_0_1_data_3 = _RAND_13[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  sectored_entries_0_1_valid_0 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  sectored_entries_0_1_valid_1 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  sectored_entries_0_1_valid_2 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  sectored_entries_0_1_valid_3 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  sectored_entries_0_2_tag = _RAND_18[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {2{`RANDOM}};
  sectored_entries_0_2_data_0 = _RAND_19[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {2{`RANDOM}};
  sectored_entries_0_2_data_1 = _RAND_20[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {2{`RANDOM}};
  sectored_entries_0_2_data_2 = _RAND_21[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {2{`RANDOM}};
  sectored_entries_0_2_data_3 = _RAND_22[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  sectored_entries_0_2_valid_0 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  sectored_entries_0_2_valid_1 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  sectored_entries_0_2_valid_2 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  sectored_entries_0_2_valid_3 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  sectored_entries_0_3_tag = _RAND_27[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {2{`RANDOM}};
  sectored_entries_0_3_data_0 = _RAND_28[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {2{`RANDOM}};
  sectored_entries_0_3_data_1 = _RAND_29[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {2{`RANDOM}};
  sectored_entries_0_3_data_2 = _RAND_30[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {2{`RANDOM}};
  sectored_entries_0_3_data_3 = _RAND_31[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  sectored_entries_0_3_valid_0 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  sectored_entries_0_3_valid_1 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  sectored_entries_0_3_valid_2 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  sectored_entries_0_3_valid_3 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  sectored_entries_0_4_tag = _RAND_36[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {2{`RANDOM}};
  sectored_entries_0_4_data_0 = _RAND_37[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {2{`RANDOM}};
  sectored_entries_0_4_data_1 = _RAND_38[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {2{`RANDOM}};
  sectored_entries_0_4_data_2 = _RAND_39[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {2{`RANDOM}};
  sectored_entries_0_4_data_3 = _RAND_40[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  sectored_entries_0_4_valid_0 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  sectored_entries_0_4_valid_1 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  sectored_entries_0_4_valid_2 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  sectored_entries_0_4_valid_3 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  sectored_entries_0_5_tag = _RAND_45[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {2{`RANDOM}};
  sectored_entries_0_5_data_0 = _RAND_46[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {2{`RANDOM}};
  sectored_entries_0_5_data_1 = _RAND_47[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {2{`RANDOM}};
  sectored_entries_0_5_data_2 = _RAND_48[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {2{`RANDOM}};
  sectored_entries_0_5_data_3 = _RAND_49[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  sectored_entries_0_5_valid_0 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  sectored_entries_0_5_valid_1 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  sectored_entries_0_5_valid_2 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  sectored_entries_0_5_valid_3 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  sectored_entries_0_6_tag = _RAND_54[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {2{`RANDOM}};
  sectored_entries_0_6_data_0 = _RAND_55[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {2{`RANDOM}};
  sectored_entries_0_6_data_1 = _RAND_56[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {2{`RANDOM}};
  sectored_entries_0_6_data_2 = _RAND_57[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {2{`RANDOM}};
  sectored_entries_0_6_data_3 = _RAND_58[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  sectored_entries_0_6_valid_0 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  sectored_entries_0_6_valid_1 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  sectored_entries_0_6_valid_2 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  sectored_entries_0_6_valid_3 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  sectored_entries_0_7_tag = _RAND_63[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {2{`RANDOM}};
  sectored_entries_0_7_data_0 = _RAND_64[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {2{`RANDOM}};
  sectored_entries_0_7_data_1 = _RAND_65[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {2{`RANDOM}};
  sectored_entries_0_7_data_2 = _RAND_66[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {2{`RANDOM}};
  sectored_entries_0_7_data_3 = _RAND_67[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  sectored_entries_0_7_valid_0 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  sectored_entries_0_7_valid_1 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  sectored_entries_0_7_valid_2 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  sectored_entries_0_7_valid_3 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  superpage_entries_0_level = _RAND_72[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  superpage_entries_0_tag = _RAND_73[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {2{`RANDOM}};
  superpage_entries_0_data_0 = _RAND_74[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  superpage_entries_0_valid_0 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  superpage_entries_1_level = _RAND_76[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  superpage_entries_1_tag = _RAND_77[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {2{`RANDOM}};
  superpage_entries_1_data_0 = _RAND_78[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  superpage_entries_1_valid_0 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  superpage_entries_2_level = _RAND_80[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  superpage_entries_2_tag = _RAND_81[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {2{`RANDOM}};
  superpage_entries_2_data_0 = _RAND_82[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  superpage_entries_2_valid_0 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  superpage_entries_3_level = _RAND_84[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  superpage_entries_3_tag = _RAND_85[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {2{`RANDOM}};
  superpage_entries_3_data_0 = _RAND_86[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  superpage_entries_3_valid_0 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  special_entry_level = _RAND_88[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  special_entry_tag = _RAND_89[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {2{`RANDOM}};
  special_entry_data_0 = _RAND_90[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  special_entry_valid_0 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  state = _RAND_92[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  r_refill_tag = _RAND_93[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  r_superpage_repl_addr = _RAND_94[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  r_sectored_repl_addr = _RAND_95[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  r_sectored_hit_addr = _RAND_96[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  r_sectored_hit = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  state_vec_0 = _RAND_98[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  state_reg_1 = _RAND_99[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  TLB_state = _RAND_100[19:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1048576; initvar = initvar+1)
    TLB_cov[initvar] = _RAND_101[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  TLB_covSum = _RAND_102[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  TLB_metaAssert = _RAND_103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      sectored_entries_0_0_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_7) begin
            sectored_entries_0_0_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_0_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_7) begin
            if (2'h0 == idx) begin
              sectored_entries_0_0_data_0 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_0_data_1 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_7) begin
            if (2'h1 == idx) begin
              sectored_entries_0_0_data_1 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_0_data_2 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_7) begin
            if (2'h2 == idx) begin
              sectored_entries_0_0_data_2 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_0_data_3 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_7) begin
            if (2'h3 == idx) begin
              sectored_entries_0_0_data_3 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_0_valid_0 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_0_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_59) begin
          if (sectored_entries_0_0_data_0[0]) begin
            sectored_entries_0_0_valid_0 <= 1'h0;
          end else if (_sector_hits_T_5) begin
            if (2'h0 == hitsVec_idx) begin
              sectored_entries_0_0_valid_0 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_7) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_0_valid_0 <= 1'h0;
                    end else begin
                      sectored_entries_0_0_valid_0 <= _GEN_53;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_7) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_0_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_0_0_valid_0 <= _GEN_53;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_5) begin
          if (2'h0 == hitsVec_idx) begin
            sectored_entries_0_0_valid_0 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_7) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_0_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_0_0_valid_0 <= _GEN_53;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_7) begin
                if (invalidate_refill) begin
                  sectored_entries_0_0_valid_0 <= 1'h0;
                end else begin
                  sectored_entries_0_0_valid_0 <= _GEN_53;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_0_valid_0 <= _GEN_621;
      end
    end else begin
      sectored_entries_0_0_valid_0 <= _GEN_473;
    end
    if (metaReset) begin
      sectored_entries_0_0_valid_1 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_0_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_59) begin
          if (sectored_entries_0_0_data_1[0]) begin
            sectored_entries_0_0_valid_1 <= 1'h0;
          end else if (_sector_hits_T_5) begin
            if (2'h1 == hitsVec_idx) begin
              sectored_entries_0_0_valid_1 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_7) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_0_valid_1 <= 1'h0;
                    end else begin
                      sectored_entries_0_0_valid_1 <= _GEN_54;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_7) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_0_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_0_0_valid_1 <= _GEN_54;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_5) begin
          if (2'h1 == hitsVec_idx) begin
            sectored_entries_0_0_valid_1 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_7) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_0_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_0_0_valid_1 <= _GEN_54;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_7) begin
                if (invalidate_refill) begin
                  sectored_entries_0_0_valid_1 <= 1'h0;
                end else begin
                  sectored_entries_0_0_valid_1 <= _GEN_54;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_0_valid_1 <= _GEN_622;
      end
    end else begin
      sectored_entries_0_0_valid_1 <= _GEN_474;
    end
    if (metaReset) begin
      sectored_entries_0_0_valid_2 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_0_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_59) begin
          if (sectored_entries_0_0_data_2[0]) begin
            sectored_entries_0_0_valid_2 <= 1'h0;
          end else if (_sector_hits_T_5) begin
            if (2'h2 == hitsVec_idx) begin
              sectored_entries_0_0_valid_2 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_7) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_0_valid_2 <= 1'h0;
                    end else begin
                      sectored_entries_0_0_valid_2 <= _GEN_55;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_7) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_0_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_0_0_valid_2 <= _GEN_55;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_5) begin
          if (2'h2 == hitsVec_idx) begin
            sectored_entries_0_0_valid_2 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_7) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_0_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_0_0_valid_2 <= _GEN_55;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_7) begin
                if (invalidate_refill) begin
                  sectored_entries_0_0_valid_2 <= 1'h0;
                end else begin
                  sectored_entries_0_0_valid_2 <= _GEN_55;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_0_valid_2 <= _GEN_623;
      end
    end else begin
      sectored_entries_0_0_valid_2 <= _GEN_475;
    end
    if (metaReset) begin
      sectored_entries_0_0_valid_3 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_0_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_59) begin
          if (sectored_entries_0_0_data_3[0]) begin
            sectored_entries_0_0_valid_3 <= 1'h0;
          end else if (_sector_hits_T_5) begin
            if (2'h3 == hitsVec_idx) begin
              sectored_entries_0_0_valid_3 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_7) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_0_valid_3 <= 1'h0;
                    end else begin
                      sectored_entries_0_0_valid_3 <= _GEN_56;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_7) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_0_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_0_0_valid_3 <= _GEN_56;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_5) begin
          if (2'h3 == hitsVec_idx) begin
            sectored_entries_0_0_valid_3 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_7) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_0_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_0_0_valid_3 <= _GEN_56;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_7) begin
                if (invalidate_refill) begin
                  sectored_entries_0_0_valid_3 <= 1'h0;
                end else begin
                  sectored_entries_0_0_valid_3 <= _GEN_56;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_0_valid_3 <= _GEN_624;
      end
    end else begin
      sectored_entries_0_0_valid_3 <= _GEN_476;
    end
    if (metaReset) begin
      sectored_entries_0_1_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_9) begin
            sectored_entries_0_1_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_1_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_9) begin
            if (2'h0 == idx) begin
              sectored_entries_0_1_data_0 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_1_data_1 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_9) begin
            if (2'h1 == idx) begin
              sectored_entries_0_1_data_1 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_1_data_2 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_9) begin
            if (2'h2 == idx) begin
              sectored_entries_0_1_data_2 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_1_data_3 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_9) begin
            if (2'h3 == idx) begin
              sectored_entries_0_1_data_3 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_1_valid_0 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_1_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_198) begin
          if (sectored_entries_0_1_data_0[0]) begin
            sectored_entries_0_1_valid_0 <= 1'h0;
          end else if (_sector_hits_T_11) begin
            if (2'h0 == hitsVec_idx) begin
              sectored_entries_0_1_valid_0 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_9) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_1_valid_0 <= 1'h0;
                    end else begin
                      sectored_entries_0_1_valid_0 <= _GEN_79;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_9) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_1_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_0_1_valid_0 <= _GEN_79;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_11) begin
          if (2'h0 == hitsVec_idx) begin
            sectored_entries_0_1_valid_0 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_9) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_1_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_0_1_valid_0 <= _GEN_79;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_9) begin
                if (invalidate_refill) begin
                  sectored_entries_0_1_valid_0 <= 1'h0;
                end else begin
                  sectored_entries_0_1_valid_0 <= _GEN_79;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_1_valid_0 <= _GEN_649;
      end
    end else begin
      sectored_entries_0_1_valid_0 <= _GEN_483;
    end
    if (metaReset) begin
      sectored_entries_0_1_valid_1 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_1_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_198) begin
          if (sectored_entries_0_1_data_1[0]) begin
            sectored_entries_0_1_valid_1 <= 1'h0;
          end else if (_sector_hits_T_11) begin
            if (2'h1 == hitsVec_idx) begin
              sectored_entries_0_1_valid_1 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_9) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_1_valid_1 <= 1'h0;
                    end else begin
                      sectored_entries_0_1_valid_1 <= _GEN_80;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_9) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_1_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_0_1_valid_1 <= _GEN_80;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_11) begin
          if (2'h1 == hitsVec_idx) begin
            sectored_entries_0_1_valid_1 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_9) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_1_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_0_1_valid_1 <= _GEN_80;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_9) begin
                if (invalidate_refill) begin
                  sectored_entries_0_1_valid_1 <= 1'h0;
                end else begin
                  sectored_entries_0_1_valid_1 <= _GEN_80;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_1_valid_1 <= _GEN_650;
      end
    end else begin
      sectored_entries_0_1_valid_1 <= _GEN_484;
    end
    if (metaReset) begin
      sectored_entries_0_1_valid_2 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_1_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_198) begin
          if (sectored_entries_0_1_data_2[0]) begin
            sectored_entries_0_1_valid_2 <= 1'h0;
          end else if (_sector_hits_T_11) begin
            if (2'h2 == hitsVec_idx) begin
              sectored_entries_0_1_valid_2 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_9) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_1_valid_2 <= 1'h0;
                    end else begin
                      sectored_entries_0_1_valid_2 <= _GEN_81;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_9) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_1_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_0_1_valid_2 <= _GEN_81;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_11) begin
          if (2'h2 == hitsVec_idx) begin
            sectored_entries_0_1_valid_2 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_9) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_1_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_0_1_valid_2 <= _GEN_81;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_9) begin
                if (invalidate_refill) begin
                  sectored_entries_0_1_valid_2 <= 1'h0;
                end else begin
                  sectored_entries_0_1_valid_2 <= _GEN_81;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_1_valid_2 <= _GEN_651;
      end
    end else begin
      sectored_entries_0_1_valid_2 <= _GEN_485;
    end
    if (metaReset) begin
      sectored_entries_0_1_valid_3 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_1_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_198) begin
          if (sectored_entries_0_1_data_3[0]) begin
            sectored_entries_0_1_valid_3 <= 1'h0;
          end else if (_sector_hits_T_11) begin
            if (2'h3 == hitsVec_idx) begin
              sectored_entries_0_1_valid_3 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_9) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_1_valid_3 <= 1'h0;
                    end else begin
                      sectored_entries_0_1_valid_3 <= _GEN_82;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_9) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_1_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_0_1_valid_3 <= _GEN_82;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_11) begin
          if (2'h3 == hitsVec_idx) begin
            sectored_entries_0_1_valid_3 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_9) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_1_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_0_1_valid_3 <= _GEN_82;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_9) begin
                if (invalidate_refill) begin
                  sectored_entries_0_1_valid_3 <= 1'h0;
                end else begin
                  sectored_entries_0_1_valid_3 <= _GEN_82;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_1_valid_3 <= _GEN_652;
      end
    end else begin
      sectored_entries_0_1_valid_3 <= _GEN_486;
    end
    if (metaReset) begin
      sectored_entries_0_2_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_11) begin
            sectored_entries_0_2_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_2_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_11) begin
            if (2'h0 == idx) begin
              sectored_entries_0_2_data_0 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_2_data_1 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_11) begin
            if (2'h1 == idx) begin
              sectored_entries_0_2_data_1 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_2_data_2 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_11) begin
            if (2'h2 == idx) begin
              sectored_entries_0_2_data_2 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_2_data_3 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_11) begin
            if (2'h3 == idx) begin
              sectored_entries_0_2_data_3 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_2_valid_0 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_2_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_337) begin
          if (sectored_entries_0_2_data_0[0]) begin
            sectored_entries_0_2_valid_0 <= 1'h0;
          end else if (_sector_hits_T_17) begin
            if (2'h0 == hitsVec_idx) begin
              sectored_entries_0_2_valid_0 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_11) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_2_valid_0 <= 1'h0;
                    end else begin
                      sectored_entries_0_2_valid_0 <= _GEN_105;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_11) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_2_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_0_2_valid_0 <= _GEN_105;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_17) begin
          if (2'h0 == hitsVec_idx) begin
            sectored_entries_0_2_valid_0 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_11) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_2_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_0_2_valid_0 <= _GEN_105;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_11) begin
                if (invalidate_refill) begin
                  sectored_entries_0_2_valid_0 <= 1'h0;
                end else begin
                  sectored_entries_0_2_valid_0 <= _GEN_105;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_2_valid_0 <= _GEN_677;
      end
    end else begin
      sectored_entries_0_2_valid_0 <= _GEN_493;
    end
    if (metaReset) begin
      sectored_entries_0_2_valid_1 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_2_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_337) begin
          if (sectored_entries_0_2_data_1[0]) begin
            sectored_entries_0_2_valid_1 <= 1'h0;
          end else if (_sector_hits_T_17) begin
            if (2'h1 == hitsVec_idx) begin
              sectored_entries_0_2_valid_1 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_11) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_2_valid_1 <= 1'h0;
                    end else begin
                      sectored_entries_0_2_valid_1 <= _GEN_106;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_11) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_2_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_0_2_valid_1 <= _GEN_106;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_17) begin
          if (2'h1 == hitsVec_idx) begin
            sectored_entries_0_2_valid_1 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_11) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_2_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_0_2_valid_1 <= _GEN_106;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_11) begin
                if (invalidate_refill) begin
                  sectored_entries_0_2_valid_1 <= 1'h0;
                end else begin
                  sectored_entries_0_2_valid_1 <= _GEN_106;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_2_valid_1 <= _GEN_678;
      end
    end else begin
      sectored_entries_0_2_valid_1 <= _GEN_494;
    end
    if (metaReset) begin
      sectored_entries_0_2_valid_2 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_2_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_337) begin
          if (sectored_entries_0_2_data_2[0]) begin
            sectored_entries_0_2_valid_2 <= 1'h0;
          end else if (_sector_hits_T_17) begin
            if (2'h2 == hitsVec_idx) begin
              sectored_entries_0_2_valid_2 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_11) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_2_valid_2 <= 1'h0;
                    end else begin
                      sectored_entries_0_2_valid_2 <= _GEN_107;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_11) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_2_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_0_2_valid_2 <= _GEN_107;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_17) begin
          if (2'h2 == hitsVec_idx) begin
            sectored_entries_0_2_valid_2 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_11) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_2_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_0_2_valid_2 <= _GEN_107;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_11) begin
                if (invalidate_refill) begin
                  sectored_entries_0_2_valid_2 <= 1'h0;
                end else begin
                  sectored_entries_0_2_valid_2 <= _GEN_107;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_2_valid_2 <= _GEN_679;
      end
    end else begin
      sectored_entries_0_2_valid_2 <= _GEN_495;
    end
    if (metaReset) begin
      sectored_entries_0_2_valid_3 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_2_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_337) begin
          if (sectored_entries_0_2_data_3[0]) begin
            sectored_entries_0_2_valid_3 <= 1'h0;
          end else if (_sector_hits_T_17) begin
            if (2'h3 == hitsVec_idx) begin
              sectored_entries_0_2_valid_3 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_11) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_2_valid_3 <= 1'h0;
                    end else begin
                      sectored_entries_0_2_valid_3 <= _GEN_108;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_11) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_2_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_0_2_valid_3 <= _GEN_108;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_17) begin
          if (2'h3 == hitsVec_idx) begin
            sectored_entries_0_2_valid_3 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_11) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_2_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_0_2_valid_3 <= _GEN_108;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_11) begin
                if (invalidate_refill) begin
                  sectored_entries_0_2_valid_3 <= 1'h0;
                end else begin
                  sectored_entries_0_2_valid_3 <= _GEN_108;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_2_valid_3 <= _GEN_680;
      end
    end else begin
      sectored_entries_0_2_valid_3 <= _GEN_496;
    end
    if (metaReset) begin
      sectored_entries_0_3_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_13) begin
            sectored_entries_0_3_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_3_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_13) begin
            if (2'h0 == idx) begin
              sectored_entries_0_3_data_0 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_3_data_1 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_13) begin
            if (2'h1 == idx) begin
              sectored_entries_0_3_data_1 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_3_data_2 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_13) begin
            if (2'h2 == idx) begin
              sectored_entries_0_3_data_2 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_3_data_3 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_13) begin
            if (2'h3 == idx) begin
              sectored_entries_0_3_data_3 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_3_valid_0 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_3_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_476) begin
          if (sectored_entries_0_3_data_0[0]) begin
            sectored_entries_0_3_valid_0 <= 1'h0;
          end else if (_sector_hits_T_23) begin
            if (2'h0 == hitsVec_idx) begin
              sectored_entries_0_3_valid_0 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_13) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_3_valid_0 <= 1'h0;
                    end else begin
                      sectored_entries_0_3_valid_0 <= _GEN_131;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_13) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_3_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_0_3_valid_0 <= _GEN_131;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_23) begin
          if (2'h0 == hitsVec_idx) begin
            sectored_entries_0_3_valid_0 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_13) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_3_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_0_3_valid_0 <= _GEN_131;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_13) begin
                if (invalidate_refill) begin
                  sectored_entries_0_3_valid_0 <= 1'h0;
                end else begin
                  sectored_entries_0_3_valid_0 <= _GEN_131;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_3_valid_0 <= _GEN_705;
      end
    end else begin
      sectored_entries_0_3_valid_0 <= _GEN_503;
    end
    if (metaReset) begin
      sectored_entries_0_3_valid_1 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_3_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_476) begin
          if (sectored_entries_0_3_data_1[0]) begin
            sectored_entries_0_3_valid_1 <= 1'h0;
          end else if (_sector_hits_T_23) begin
            if (2'h1 == hitsVec_idx) begin
              sectored_entries_0_3_valid_1 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_13) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_3_valid_1 <= 1'h0;
                    end else begin
                      sectored_entries_0_3_valid_1 <= _GEN_132;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_13) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_3_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_0_3_valid_1 <= _GEN_132;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_23) begin
          if (2'h1 == hitsVec_idx) begin
            sectored_entries_0_3_valid_1 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_13) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_3_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_0_3_valid_1 <= _GEN_132;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_13) begin
                if (invalidate_refill) begin
                  sectored_entries_0_3_valid_1 <= 1'h0;
                end else begin
                  sectored_entries_0_3_valid_1 <= _GEN_132;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_3_valid_1 <= _GEN_706;
      end
    end else begin
      sectored_entries_0_3_valid_1 <= _GEN_504;
    end
    if (metaReset) begin
      sectored_entries_0_3_valid_2 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_3_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_476) begin
          if (sectored_entries_0_3_data_2[0]) begin
            sectored_entries_0_3_valid_2 <= 1'h0;
          end else if (_sector_hits_T_23) begin
            if (2'h2 == hitsVec_idx) begin
              sectored_entries_0_3_valid_2 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_13) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_3_valid_2 <= 1'h0;
                    end else begin
                      sectored_entries_0_3_valid_2 <= _GEN_133;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_13) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_3_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_0_3_valid_2 <= _GEN_133;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_23) begin
          if (2'h2 == hitsVec_idx) begin
            sectored_entries_0_3_valid_2 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_13) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_3_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_0_3_valid_2 <= _GEN_133;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_13) begin
                if (invalidate_refill) begin
                  sectored_entries_0_3_valid_2 <= 1'h0;
                end else begin
                  sectored_entries_0_3_valid_2 <= _GEN_133;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_3_valid_2 <= _GEN_707;
      end
    end else begin
      sectored_entries_0_3_valid_2 <= _GEN_505;
    end
    if (metaReset) begin
      sectored_entries_0_3_valid_3 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_3_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_476) begin
          if (sectored_entries_0_3_data_3[0]) begin
            sectored_entries_0_3_valid_3 <= 1'h0;
          end else if (_sector_hits_T_23) begin
            if (2'h3 == hitsVec_idx) begin
              sectored_entries_0_3_valid_3 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_13) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_3_valid_3 <= 1'h0;
                    end else begin
                      sectored_entries_0_3_valid_3 <= _GEN_134;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_13) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_3_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_0_3_valid_3 <= _GEN_134;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_23) begin
          if (2'h3 == hitsVec_idx) begin
            sectored_entries_0_3_valid_3 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_13) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_3_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_0_3_valid_3 <= _GEN_134;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_13) begin
                if (invalidate_refill) begin
                  sectored_entries_0_3_valid_3 <= 1'h0;
                end else begin
                  sectored_entries_0_3_valid_3 <= _GEN_134;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_3_valid_3 <= _GEN_708;
      end
    end else begin
      sectored_entries_0_3_valid_3 <= _GEN_506;
    end
    if (metaReset) begin
      sectored_entries_0_4_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_15) begin
            sectored_entries_0_4_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_4_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_15) begin
            if (2'h0 == idx) begin
              sectored_entries_0_4_data_0 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_4_data_1 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_15) begin
            if (2'h1 == idx) begin
              sectored_entries_0_4_data_1 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_4_data_2 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_15) begin
            if (2'h2 == idx) begin
              sectored_entries_0_4_data_2 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_4_data_3 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_15) begin
            if (2'h3 == idx) begin
              sectored_entries_0_4_data_3 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_4_valid_0 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_4_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_615) begin
          if (sectored_entries_0_4_data_0[0]) begin
            sectored_entries_0_4_valid_0 <= 1'h0;
          end else if (_sector_hits_T_29) begin
            if (2'h0 == hitsVec_idx) begin
              sectored_entries_0_4_valid_0 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_15) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_4_valid_0 <= 1'h0;
                    end else begin
                      sectored_entries_0_4_valid_0 <= _GEN_157;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_15) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_4_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_0_4_valid_0 <= _GEN_157;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_29) begin
          if (2'h0 == hitsVec_idx) begin
            sectored_entries_0_4_valid_0 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_15) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_4_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_0_4_valid_0 <= _GEN_157;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_15) begin
                if (invalidate_refill) begin
                  sectored_entries_0_4_valid_0 <= 1'h0;
                end else begin
                  sectored_entries_0_4_valid_0 <= _GEN_157;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_4_valid_0 <= _GEN_733;
      end
    end else begin
      sectored_entries_0_4_valid_0 <= _GEN_513;
    end
    if (metaReset) begin
      sectored_entries_0_4_valid_1 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_4_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_615) begin
          if (sectored_entries_0_4_data_1[0]) begin
            sectored_entries_0_4_valid_1 <= 1'h0;
          end else if (_sector_hits_T_29) begin
            if (2'h1 == hitsVec_idx) begin
              sectored_entries_0_4_valid_1 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_15) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_4_valid_1 <= 1'h0;
                    end else begin
                      sectored_entries_0_4_valid_1 <= _GEN_158;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_15) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_4_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_0_4_valid_1 <= _GEN_158;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_29) begin
          if (2'h1 == hitsVec_idx) begin
            sectored_entries_0_4_valid_1 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_15) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_4_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_0_4_valid_1 <= _GEN_158;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_15) begin
                if (invalidate_refill) begin
                  sectored_entries_0_4_valid_1 <= 1'h0;
                end else begin
                  sectored_entries_0_4_valid_1 <= _GEN_158;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_4_valid_1 <= _GEN_734;
      end
    end else begin
      sectored_entries_0_4_valid_1 <= _GEN_514;
    end
    if (metaReset) begin
      sectored_entries_0_4_valid_2 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_4_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_615) begin
          if (sectored_entries_0_4_data_2[0]) begin
            sectored_entries_0_4_valid_2 <= 1'h0;
          end else if (_sector_hits_T_29) begin
            if (2'h2 == hitsVec_idx) begin
              sectored_entries_0_4_valid_2 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_15) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_4_valid_2 <= 1'h0;
                    end else begin
                      sectored_entries_0_4_valid_2 <= _GEN_159;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_15) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_4_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_0_4_valid_2 <= _GEN_159;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_29) begin
          if (2'h2 == hitsVec_idx) begin
            sectored_entries_0_4_valid_2 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_15) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_4_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_0_4_valid_2 <= _GEN_159;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_15) begin
                if (invalidate_refill) begin
                  sectored_entries_0_4_valid_2 <= 1'h0;
                end else begin
                  sectored_entries_0_4_valid_2 <= _GEN_159;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_4_valid_2 <= _GEN_735;
      end
    end else begin
      sectored_entries_0_4_valid_2 <= _GEN_515;
    end
    if (metaReset) begin
      sectored_entries_0_4_valid_3 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_4_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_615) begin
          if (sectored_entries_0_4_data_3[0]) begin
            sectored_entries_0_4_valid_3 <= 1'h0;
          end else if (_sector_hits_T_29) begin
            if (2'h3 == hitsVec_idx) begin
              sectored_entries_0_4_valid_3 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_15) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_4_valid_3 <= 1'h0;
                    end else begin
                      sectored_entries_0_4_valid_3 <= _GEN_160;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_15) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_4_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_0_4_valid_3 <= _GEN_160;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_29) begin
          if (2'h3 == hitsVec_idx) begin
            sectored_entries_0_4_valid_3 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_15) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_4_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_0_4_valid_3 <= _GEN_160;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_15) begin
                if (invalidate_refill) begin
                  sectored_entries_0_4_valid_3 <= 1'h0;
                end else begin
                  sectored_entries_0_4_valid_3 <= _GEN_160;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_4_valid_3 <= _GEN_736;
      end
    end else begin
      sectored_entries_0_4_valid_3 <= _GEN_516;
    end
    if (metaReset) begin
      sectored_entries_0_5_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_17) begin
            sectored_entries_0_5_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_5_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_17) begin
            if (2'h0 == idx) begin
              sectored_entries_0_5_data_0 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_5_data_1 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_17) begin
            if (2'h1 == idx) begin
              sectored_entries_0_5_data_1 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_5_data_2 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_17) begin
            if (2'h2 == idx) begin
              sectored_entries_0_5_data_2 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_5_data_3 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_17) begin
            if (2'h3 == idx) begin
              sectored_entries_0_5_data_3 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_5_valid_0 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_5_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_754) begin
          if (sectored_entries_0_5_data_0[0]) begin
            sectored_entries_0_5_valid_0 <= 1'h0;
          end else if (_sector_hits_T_35) begin
            if (2'h0 == hitsVec_idx) begin
              sectored_entries_0_5_valid_0 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_17) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_5_valid_0 <= 1'h0;
                    end else begin
                      sectored_entries_0_5_valid_0 <= _GEN_183;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_17) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_5_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_0_5_valid_0 <= _GEN_183;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_35) begin
          if (2'h0 == hitsVec_idx) begin
            sectored_entries_0_5_valid_0 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_17) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_5_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_0_5_valid_0 <= _GEN_183;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_17) begin
                if (invalidate_refill) begin
                  sectored_entries_0_5_valid_0 <= 1'h0;
                end else begin
                  sectored_entries_0_5_valid_0 <= _GEN_183;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_5_valid_0 <= _GEN_761;
      end
    end else begin
      sectored_entries_0_5_valid_0 <= _GEN_523;
    end
    if (metaReset) begin
      sectored_entries_0_5_valid_1 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_5_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_754) begin
          if (sectored_entries_0_5_data_1[0]) begin
            sectored_entries_0_5_valid_1 <= 1'h0;
          end else if (_sector_hits_T_35) begin
            if (2'h1 == hitsVec_idx) begin
              sectored_entries_0_5_valid_1 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_17) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_5_valid_1 <= 1'h0;
                    end else begin
                      sectored_entries_0_5_valid_1 <= _GEN_184;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_17) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_5_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_0_5_valid_1 <= _GEN_184;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_35) begin
          if (2'h1 == hitsVec_idx) begin
            sectored_entries_0_5_valid_1 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_17) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_5_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_0_5_valid_1 <= _GEN_184;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_17) begin
                if (invalidate_refill) begin
                  sectored_entries_0_5_valid_1 <= 1'h0;
                end else begin
                  sectored_entries_0_5_valid_1 <= _GEN_184;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_5_valid_1 <= _GEN_762;
      end
    end else begin
      sectored_entries_0_5_valid_1 <= _GEN_524;
    end
    if (metaReset) begin
      sectored_entries_0_5_valid_2 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_5_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_754) begin
          if (sectored_entries_0_5_data_2[0]) begin
            sectored_entries_0_5_valid_2 <= 1'h0;
          end else if (_sector_hits_T_35) begin
            if (2'h2 == hitsVec_idx) begin
              sectored_entries_0_5_valid_2 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_17) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_5_valid_2 <= 1'h0;
                    end else begin
                      sectored_entries_0_5_valid_2 <= _GEN_185;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_17) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_5_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_0_5_valid_2 <= _GEN_185;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_35) begin
          if (2'h2 == hitsVec_idx) begin
            sectored_entries_0_5_valid_2 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_17) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_5_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_0_5_valid_2 <= _GEN_185;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_17) begin
                if (invalidate_refill) begin
                  sectored_entries_0_5_valid_2 <= 1'h0;
                end else begin
                  sectored_entries_0_5_valid_2 <= _GEN_185;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_5_valid_2 <= _GEN_763;
      end
    end else begin
      sectored_entries_0_5_valid_2 <= _GEN_525;
    end
    if (metaReset) begin
      sectored_entries_0_5_valid_3 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_5_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_754) begin
          if (sectored_entries_0_5_data_3[0]) begin
            sectored_entries_0_5_valid_3 <= 1'h0;
          end else if (_sector_hits_T_35) begin
            if (2'h3 == hitsVec_idx) begin
              sectored_entries_0_5_valid_3 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_17) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_5_valid_3 <= 1'h0;
                    end else begin
                      sectored_entries_0_5_valid_3 <= _GEN_186;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_17) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_5_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_0_5_valid_3 <= _GEN_186;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_35) begin
          if (2'h3 == hitsVec_idx) begin
            sectored_entries_0_5_valid_3 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_17) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_5_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_0_5_valid_3 <= _GEN_186;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_17) begin
                if (invalidate_refill) begin
                  sectored_entries_0_5_valid_3 <= 1'h0;
                end else begin
                  sectored_entries_0_5_valid_3 <= _GEN_186;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_5_valid_3 <= _GEN_764;
      end
    end else begin
      sectored_entries_0_5_valid_3 <= _GEN_526;
    end
    if (metaReset) begin
      sectored_entries_0_6_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_19) begin
            sectored_entries_0_6_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_6_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_19) begin
            if (2'h0 == idx) begin
              sectored_entries_0_6_data_0 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_6_data_1 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_19) begin
            if (2'h1 == idx) begin
              sectored_entries_0_6_data_1 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_6_data_2 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_19) begin
            if (2'h2 == idx) begin
              sectored_entries_0_6_data_2 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_6_data_3 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_19) begin
            if (2'h3 == idx) begin
              sectored_entries_0_6_data_3 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_6_valid_0 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_6_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_893) begin
          if (sectored_entries_0_6_data_0[0]) begin
            sectored_entries_0_6_valid_0 <= 1'h0;
          end else if (_sector_hits_T_41) begin
            if (2'h0 == hitsVec_idx) begin
              sectored_entries_0_6_valid_0 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_19) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_6_valid_0 <= 1'h0;
                    end else begin
                      sectored_entries_0_6_valid_0 <= _GEN_209;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_19) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_6_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_0_6_valid_0 <= _GEN_209;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_41) begin
          if (2'h0 == hitsVec_idx) begin
            sectored_entries_0_6_valid_0 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_19) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_6_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_0_6_valid_0 <= _GEN_209;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_19) begin
                if (invalidate_refill) begin
                  sectored_entries_0_6_valid_0 <= 1'h0;
                end else begin
                  sectored_entries_0_6_valid_0 <= _GEN_209;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_6_valid_0 <= _GEN_789;
      end
    end else begin
      sectored_entries_0_6_valid_0 <= _GEN_533;
    end
    if (metaReset) begin
      sectored_entries_0_6_valid_1 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_6_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_893) begin
          if (sectored_entries_0_6_data_1[0]) begin
            sectored_entries_0_6_valid_1 <= 1'h0;
          end else if (_sector_hits_T_41) begin
            if (2'h1 == hitsVec_idx) begin
              sectored_entries_0_6_valid_1 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_19) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_6_valid_1 <= 1'h0;
                    end else begin
                      sectored_entries_0_6_valid_1 <= _GEN_210;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_19) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_6_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_0_6_valid_1 <= _GEN_210;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_41) begin
          if (2'h1 == hitsVec_idx) begin
            sectored_entries_0_6_valid_1 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_19) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_6_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_0_6_valid_1 <= _GEN_210;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_19) begin
                if (invalidate_refill) begin
                  sectored_entries_0_6_valid_1 <= 1'h0;
                end else begin
                  sectored_entries_0_6_valid_1 <= _GEN_210;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_6_valid_1 <= _GEN_790;
      end
    end else begin
      sectored_entries_0_6_valid_1 <= _GEN_534;
    end
    if (metaReset) begin
      sectored_entries_0_6_valid_2 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_6_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_893) begin
          if (sectored_entries_0_6_data_2[0]) begin
            sectored_entries_0_6_valid_2 <= 1'h0;
          end else if (_sector_hits_T_41) begin
            if (2'h2 == hitsVec_idx) begin
              sectored_entries_0_6_valid_2 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_19) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_6_valid_2 <= 1'h0;
                    end else begin
                      sectored_entries_0_6_valid_2 <= _GEN_211;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_19) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_6_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_0_6_valid_2 <= _GEN_211;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_41) begin
          if (2'h2 == hitsVec_idx) begin
            sectored_entries_0_6_valid_2 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_19) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_6_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_0_6_valid_2 <= _GEN_211;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_19) begin
                if (invalidate_refill) begin
                  sectored_entries_0_6_valid_2 <= 1'h0;
                end else begin
                  sectored_entries_0_6_valid_2 <= _GEN_211;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_6_valid_2 <= _GEN_791;
      end
    end else begin
      sectored_entries_0_6_valid_2 <= _GEN_535;
    end
    if (metaReset) begin
      sectored_entries_0_6_valid_3 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_6_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_893) begin
          if (sectored_entries_0_6_data_3[0]) begin
            sectored_entries_0_6_valid_3 <= 1'h0;
          end else if (_sector_hits_T_41) begin
            if (2'h3 == hitsVec_idx) begin
              sectored_entries_0_6_valid_3 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_19) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_6_valid_3 <= 1'h0;
                    end else begin
                      sectored_entries_0_6_valid_3 <= _GEN_212;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_19) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_6_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_0_6_valid_3 <= _GEN_212;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_41) begin
          if (2'h3 == hitsVec_idx) begin
            sectored_entries_0_6_valid_3 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_19) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_6_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_0_6_valid_3 <= _GEN_212;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_19) begin
                if (invalidate_refill) begin
                  sectored_entries_0_6_valid_3 <= 1'h0;
                end else begin
                  sectored_entries_0_6_valid_3 <= _GEN_212;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_6_valid_3 <= _GEN_792;
      end
    end else begin
      sectored_entries_0_6_valid_3 <= _GEN_536;
    end
    if (metaReset) begin
      sectored_entries_0_7_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_21) begin
            sectored_entries_0_7_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_7_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_21) begin
            if (2'h0 == idx) begin
              sectored_entries_0_7_data_0 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_7_data_1 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_21) begin
            if (2'h1 == idx) begin
              sectored_entries_0_7_data_1 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_7_data_2 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_21) begin
            if (2'h2 == idx) begin
              sectored_entries_0_7_data_2 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_7_data_3 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_21) begin
            if (2'h3 == idx) begin
              sectored_entries_0_7_data_3 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_7_valid_0 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_7_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_1032) begin
          if (sectored_entries_0_7_data_0[0]) begin
            sectored_entries_0_7_valid_0 <= 1'h0;
          end else if (_sector_hits_T_47) begin
            if (2'h0 == hitsVec_idx) begin
              sectored_entries_0_7_valid_0 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_21) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_7_valid_0 <= 1'h0;
                    end else begin
                      sectored_entries_0_7_valid_0 <= _GEN_235;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_21) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_7_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_0_7_valid_0 <= _GEN_235;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_47) begin
          if (2'h0 == hitsVec_idx) begin
            sectored_entries_0_7_valid_0 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_21) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_7_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_0_7_valid_0 <= _GEN_235;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_21) begin
                if (invalidate_refill) begin
                  sectored_entries_0_7_valid_0 <= 1'h0;
                end else begin
                  sectored_entries_0_7_valid_0 <= _GEN_235;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_7_valid_0 <= _GEN_817;
      end
    end else begin
      sectored_entries_0_7_valid_0 <= _GEN_543;
    end
    if (metaReset) begin
      sectored_entries_0_7_valid_1 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_7_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_1032) begin
          if (sectored_entries_0_7_data_1[0]) begin
            sectored_entries_0_7_valid_1 <= 1'h0;
          end else if (_sector_hits_T_47) begin
            if (2'h1 == hitsVec_idx) begin
              sectored_entries_0_7_valid_1 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_21) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_7_valid_1 <= 1'h0;
                    end else begin
                      sectored_entries_0_7_valid_1 <= _GEN_236;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_21) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_7_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_0_7_valid_1 <= _GEN_236;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_47) begin
          if (2'h1 == hitsVec_idx) begin
            sectored_entries_0_7_valid_1 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_21) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_7_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_0_7_valid_1 <= _GEN_236;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_21) begin
                if (invalidate_refill) begin
                  sectored_entries_0_7_valid_1 <= 1'h0;
                end else begin
                  sectored_entries_0_7_valid_1 <= _GEN_236;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_7_valid_1 <= _GEN_818;
      end
    end else begin
      sectored_entries_0_7_valid_1 <= _GEN_544;
    end
    if (metaReset) begin
      sectored_entries_0_7_valid_2 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_7_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_1032) begin
          if (sectored_entries_0_7_data_2[0]) begin
            sectored_entries_0_7_valid_2 <= 1'h0;
          end else if (_sector_hits_T_47) begin
            if (2'h2 == hitsVec_idx) begin
              sectored_entries_0_7_valid_2 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_21) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_7_valid_2 <= 1'h0;
                    end else begin
                      sectored_entries_0_7_valid_2 <= _GEN_237;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_21) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_7_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_0_7_valid_2 <= _GEN_237;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_47) begin
          if (2'h2 == hitsVec_idx) begin
            sectored_entries_0_7_valid_2 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_21) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_7_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_0_7_valid_2 <= _GEN_237;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_21) begin
                if (invalidate_refill) begin
                  sectored_entries_0_7_valid_2 <= 1'h0;
                end else begin
                  sectored_entries_0_7_valid_2 <= _GEN_237;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_7_valid_2 <= _GEN_819;
      end
    end else begin
      sectored_entries_0_7_valid_2 <= _GEN_545;
    end
    if (metaReset) begin
      sectored_entries_0_7_valid_3 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_7_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_1032) begin
          if (sectored_entries_0_7_data_3[0]) begin
            sectored_entries_0_7_valid_3 <= 1'h0;
          end else if (_sector_hits_T_47) begin
            if (2'h3 == hitsVec_idx) begin
              sectored_entries_0_7_valid_3 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_21) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_7_valid_3 <= 1'h0;
                    end else begin
                      sectored_entries_0_7_valid_3 <= _GEN_238;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_21) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_7_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_0_7_valid_3 <= _GEN_238;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_47) begin
          if (2'h3 == hitsVec_idx) begin
            sectored_entries_0_7_valid_3 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_21) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_7_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_0_7_valid_3 <= _GEN_238;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_21) begin
                if (invalidate_refill) begin
                  sectored_entries_0_7_valid_3 <= 1'h0;
                end else begin
                  sectored_entries_0_7_valid_3 <= _GEN_238;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_7_valid_3 <= _GEN_820;
      end
    end else begin
      sectored_entries_0_7_valid_3 <= _GEN_546;
    end
    if (metaReset) begin
      superpage_entries_0_level <= 2'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_2) begin
          if (_T_3) begin
            superpage_entries_0_level <= {{1'd0}, io_ptw_resp_bits_level[0]};
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_0_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_2) begin
          if (_T_3) begin
            superpage_entries_0_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_0_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_2) begin
          if (_T_3) begin
            superpage_entries_0_data_0 <= _special_entry_data_0_T;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_0_valid_0 <= 1'h0;
    end else if (_T_1326) begin
      superpage_entries_0_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (superpage_hits_0) begin
          superpage_entries_0_valid_0 <= 1'h0;
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (_T_2) begin
              if (_T_3) begin
                if (invalidate_refill) begin
                  superpage_entries_0_valid_0 <= 1'h0;
                end else begin
                  superpage_entries_0_valid_0 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        superpage_entries_0_valid_0 <= _GEN_827;
      end
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_2) begin
          if (_T_3) begin
            if (invalidate_refill) begin
              superpage_entries_0_valid_0 <= 1'h0;
            end else begin
              superpage_entries_0_valid_0 <= 1'h1;
            end
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_1_level <= 2'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_2) begin
          if (_T_4) begin
            superpage_entries_1_level <= {{1'd0}, io_ptw_resp_bits_level[0]};
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_1_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_2) begin
          if (_T_4) begin
            superpage_entries_1_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_1_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_2) begin
          if (_T_4) begin
            superpage_entries_1_data_0 <= _special_entry_data_0_T;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_1_valid_0 <= 1'h0;
    end else if (_T_1326) begin
      superpage_entries_1_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (superpage_hits_1) begin
          superpage_entries_1_valid_0 <= 1'h0;
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (_T_2) begin
              if (_T_4) begin
                if (invalidate_refill) begin
                  superpage_entries_1_valid_0 <= 1'h0;
                end else begin
                  superpage_entries_1_valid_0 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        superpage_entries_1_valid_0 <= _GEN_831;
      end
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_2) begin
          if (_T_4) begin
            if (invalidate_refill) begin
              superpage_entries_1_valid_0 <= 1'h0;
            end else begin
              superpage_entries_1_valid_0 <= 1'h1;
            end
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_2_level <= 2'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_2) begin
          if (_T_5) begin
            superpage_entries_2_level <= {{1'd0}, io_ptw_resp_bits_level[0]};
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_2_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_2) begin
          if (_T_5) begin
            superpage_entries_2_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_2_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_2) begin
          if (_T_5) begin
            superpage_entries_2_data_0 <= _special_entry_data_0_T;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_2_valid_0 <= 1'h0;
    end else if (_T_1326) begin
      superpage_entries_2_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (superpage_hits_2) begin
          superpage_entries_2_valid_0 <= 1'h0;
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (_T_2) begin
              if (_T_5) begin
                superpage_entries_2_valid_0 <= _GEN_32;
              end
            end
          end
        end
      end else begin
        superpage_entries_2_valid_0 <= _GEN_835;
      end
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_2) begin
          if (_T_5) begin
            superpage_entries_2_valid_0 <= _GEN_32;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_3_level <= 2'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_2) begin
          if (_T_6) begin
            superpage_entries_3_level <= {{1'd0}, io_ptw_resp_bits_level[0]};
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_3_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_2) begin
          if (_T_6) begin
            superpage_entries_3_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_3_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_2) begin
          if (_T_6) begin
            superpage_entries_3_data_0 <= _special_entry_data_0_T;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_3_valid_0 <= 1'h0;
    end else if (_T_1326) begin
      superpage_entries_3_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (superpage_hits_3) begin
          superpage_entries_3_valid_0 <= 1'h0;
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (_T_2) begin
              if (_T_6) begin
                superpage_entries_3_valid_0 <= _GEN_32;
              end
            end
          end
        end
      end else begin
        superpage_entries_3_valid_0 <= _GEN_839;
      end
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_2) begin
          if (_T_6) begin
            superpage_entries_3_valid_0 <= _GEN_32;
          end
        end
      end
    end
    if (metaReset) begin
      special_entry_level <= 2'h0;
    end else if (io_ptw_resp_valid) begin
      if (~io_ptw_resp_bits_homogeneous) begin
        special_entry_level <= io_ptw_resp_bits_level;
      end
    end
    if (metaReset) begin
      special_entry_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (~io_ptw_resp_bits_homogeneous) begin
        special_entry_tag <= r_refill_tag;
      end
    end
    if (metaReset) begin
      special_entry_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (~io_ptw_resp_bits_homogeneous) begin
        special_entry_data_0 <= _special_entry_data_0_T;
      end
    end
    if (metaReset) begin
      special_entry_valid_0 <= 1'h0;
    end else if (_T_1326) begin
      special_entry_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_hitsVec_T_106) begin
          special_entry_valid_0 <= 1'h0;
        end else if (io_ptw_resp_valid) begin
          if (~io_ptw_resp_bits_homogeneous) begin
            special_entry_valid_0 <= _GEN_32;
          end
        end
      end else begin
        special_entry_valid_0 <= _GEN_843;
      end
    end else if (io_ptw_resp_valid) begin
      if (~io_ptw_resp_bits_homogeneous) begin
        special_entry_valid_0 <= _GEN_32;
      end
    end
    if (metaReset) begin
      state <= 2'h0;
    end else if (reset) begin
      state <= 2'h0;
    end else if (io_ptw_resp_valid) begin
      state <= 2'h0;
    end else if (_T_45) begin
      state <= 2'h3;
    end else if (_invalidate_refill_T) begin
      if (io_ptw_req_ready) begin
        if (io_sfence_valid) begin
          state <= 2'h3;
        end else begin
          state <= 2'h2;
        end
      end else if (io_sfence_valid) begin
        state <= 2'h0;
      end else if (_T_42) begin
        state <= 2'h1;
      end
    end else if (_T_42) begin
      state <= 2'h1;
    end
    if (metaReset) begin
      r_refill_tag <= 27'h0;
    end else if (_T_42) begin
      r_refill_tag <= vpn;
    end
    if (metaReset) begin
      r_superpage_repl_addr <= 2'h0;
    end else if (_T_42) begin
      if (_r_superpage_repl_addr_T_3) begin
        r_superpage_repl_addr <= _r_superpage_repl_addr_T_2;
      end else if (_r_superpage_repl_addr_T_5) begin
        r_superpage_repl_addr <= 2'h0;
      end else if (_r_superpage_repl_addr_T_6) begin
        r_superpage_repl_addr <= 2'h1;
      end else if (_r_superpage_repl_addr_T_7) begin
        r_superpage_repl_addr <= 2'h2;
      end else begin
        r_superpage_repl_addr <= 2'h3;
      end
    end
    if (metaReset) begin
      r_sectored_repl_addr <= 3'h0;
    end else if (_T_42) begin
      if (_r_sectored_repl_addr_T_7) begin
        r_sectored_repl_addr <= _r_sectored_repl_addr_T_6;
      end else if (_r_sectored_repl_addr_T_9) begin
        r_sectored_repl_addr <= 3'h0;
      end else if (_r_sectored_repl_addr_T_10) begin
        r_sectored_repl_addr <= 3'h1;
      end else if (_r_sectored_repl_addr_T_11) begin
        r_sectored_repl_addr <= 3'h2;
      end else if (_r_sectored_repl_addr_T_12) begin
        r_sectored_repl_addr <= 3'h3;
      end else if (_r_sectored_repl_addr_T_13) begin
        r_sectored_repl_addr <= 3'h4;
      end else if (_r_sectored_repl_addr_T_14) begin
        r_sectored_repl_addr <= 3'h5;
      end else if (_r_sectored_repl_addr_T_15) begin
        r_sectored_repl_addr <= 3'h6;
      end else begin
        r_sectored_repl_addr <= 3'h7;
      end
    end
    if (metaReset) begin
      r_sectored_hit_addr <= 3'h0;
    end else if (_T_42) begin
      r_sectored_hit_addr <= state_vec_0_touch_way_sized;
    end
    if (metaReset) begin
      r_sectored_hit <= 1'h0;
    end else if (_T_42) begin
      r_sectored_hit <= _T_30;
    end
    if (metaReset) begin
      state_vec_0 <= 7'h0;
    end else if (reset) begin
      state_vec_0 <= 7'h0;
    end else if (_T_23) begin
      if (_T_30) begin
        state_vec_0 <= _state_vec_0_T_16;
      end
    end
    if (metaReset) begin
      state_reg_1 <= 3'h0;
    end else if (reset) begin
      state_reg_1 <= 3'h0;
    end else if (_T_23) begin
      if (_T_37) begin
        state_reg_1 <= _state_reg_T_6;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_sfence_valid & ~_T_51) begin
          $fwrite(32'h80000002,"Assertion failed\n    at TLB.scala:385 assert(!io.sfence.bits.rs1 || (io.sfence.bits.addr >> pgIdxBits) === vpn)\n"); // @[TLB.scala 385:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_sfence_valid & ~_T_51) begin
          $fatal; // @[TLB.scala 385:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    TLB_state <= TLB_xor0;
    if (!(TLB_cov_read_data)) begin
      TLB_covSum <= TLB_covSum + 1'h1;
    end
    if (metaReset) begin
      TLB_metaAssert <= 1'h0;
    end else begin
      TLB_metaAssert <= TLB_metaAssert | TLB_or0;
    end
  end
  always @(posedge clock) begin
    if(TLB_cov_write_en & TLB_cov_write_mask) begin
      TLB_cov[TLB_cov_write_addr] <= TLB_cov_write_data; // @[Coverage map for TLB]
    end
  end
endmodule
module MaxPeriodFibonacciLFSR(
  input         clock,
  input         reset,
  input         io_increment,
  output        io_out_0,
  output        io_out_1,
  output        io_out_2,
  output        io_out_3,
  output        io_out_4,
  output        io_out_5,
  output        io_out_6,
  output        io_out_7,
  output        io_out_8,
  output        io_out_9,
  output        io_out_10,
  output        io_out_11,
  output        io_out_12,
  output        io_out_13,
  output        io_out_14,
  output        io_out_15,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  reg  state_0; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_0;
  reg  state_1; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_1;
  reg  state_2; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_2;
  reg  state_3; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_3;
  reg  state_4; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_4;
  reg  state_5; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_5;
  reg  state_6; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_6;
  reg  state_7; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_7;
  reg  state_8; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_8;
  reg  state_9; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_9;
  reg  state_10; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_10;
  reg  state_11; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_11;
  reg  state_12; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_12;
  reg  state_13; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_13;
  reg  state_14; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_14;
  reg  state_15; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_15;
  wire  _T; // @[LFSR.scala 15:41]
  wire  _T_1; // @[LFSR.scala 15:41]
  wire  _T_2; // @[LFSR.scala 15:41]
  wire  _GEN_0; // @[PRNG.scala 61:23]
  wire [29:0] MaxPeriodFibonacciLFSR_covSum;
  assign _T = state_15 ^ state_13; // @[LFSR.scala 15:41]
  assign _T_1 = _T ^ state_12; // @[LFSR.scala 15:41]
  assign _T_2 = _T_1 ^ state_10; // @[LFSR.scala 15:41]
  assign _GEN_0 = io_increment ? _T_2 : state_0; // @[PRNG.scala 61:23]
  assign io_out_0 = state_0; // @[PRNG.scala 69:10]
  assign io_out_1 = state_1; // @[PRNG.scala 69:10]
  assign io_out_2 = state_2; // @[PRNG.scala 69:10]
  assign io_out_3 = state_3; // @[PRNG.scala 69:10]
  assign io_out_4 = state_4; // @[PRNG.scala 69:10]
  assign io_out_5 = state_5; // @[PRNG.scala 69:10]
  assign io_out_6 = state_6; // @[PRNG.scala 69:10]
  assign io_out_7 = state_7; // @[PRNG.scala 69:10]
  assign io_out_8 = state_8; // @[PRNG.scala 69:10]
  assign io_out_9 = state_9; // @[PRNG.scala 69:10]
  assign io_out_10 = state_10; // @[PRNG.scala 69:10]
  assign io_out_11 = state_11; // @[PRNG.scala 69:10]
  assign io_out_12 = state_12; // @[PRNG.scala 69:10]
  assign io_out_13 = state_13; // @[PRNG.scala 69:10]
  assign io_out_14 = state_14; // @[PRNG.scala 69:10]
  assign io_out_15 = state_15; // @[PRNG.scala 69:10]
  assign MaxPeriodFibonacciLFSR_covSum = 30'h0;
  assign io_covSum = MaxPeriodFibonacciLFSR_covSum;
  assign metaAssert = 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  state_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  state_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  state_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  state_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  state_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  state_6 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  state_7 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  state_8 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  state_9 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state_10 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state_11 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  state_12 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  state_13 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  state_14 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  state_15 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      state_0 <= 1'h0;
    end else begin
      state_0 <= reset | _GEN_0;
    end
    if (metaReset) begin
      state_1 <= 1'h0;
    end else if (reset) begin
      state_1 <= 1'h0;
    end else if (io_increment) begin
      state_1 <= state_0;
    end
    if (metaReset) begin
      state_2 <= 1'h0;
    end else if (reset) begin
      state_2 <= 1'h0;
    end else if (io_increment) begin
      state_2 <= state_1;
    end
    if (metaReset) begin
      state_3 <= 1'h0;
    end else if (reset) begin
      state_3 <= 1'h0;
    end else if (io_increment) begin
      state_3 <= state_2;
    end
    if (metaReset) begin
      state_4 <= 1'h0;
    end else if (reset) begin
      state_4 <= 1'h0;
    end else if (io_increment) begin
      state_4 <= state_3;
    end
    if (metaReset) begin
      state_5 <= 1'h0;
    end else if (reset) begin
      state_5 <= 1'h0;
    end else if (io_increment) begin
      state_5 <= state_4;
    end
    if (metaReset) begin
      state_6 <= 1'h0;
    end else if (reset) begin
      state_6 <= 1'h0;
    end else if (io_increment) begin
      state_6 <= state_5;
    end
    if (metaReset) begin
      state_7 <= 1'h0;
    end else if (reset) begin
      state_7 <= 1'h0;
    end else if (io_increment) begin
      state_7 <= state_6;
    end
    if (metaReset) begin
      state_8 <= 1'h0;
    end else if (reset) begin
      state_8 <= 1'h0;
    end else if (io_increment) begin
      state_8 <= state_7;
    end
    if (metaReset) begin
      state_9 <= 1'h0;
    end else if (reset) begin
      state_9 <= 1'h0;
    end else if (io_increment) begin
      state_9 <= state_8;
    end
    if (metaReset) begin
      state_10 <= 1'h0;
    end else if (reset) begin
      state_10 <= 1'h0;
    end else if (io_increment) begin
      state_10 <= state_9;
    end
    if (metaReset) begin
      state_11 <= 1'h0;
    end else if (reset) begin
      state_11 <= 1'h0;
    end else if (io_increment) begin
      state_11 <= state_10;
    end
    if (metaReset) begin
      state_12 <= 1'h0;
    end else if (reset) begin
      state_12 <= 1'h0;
    end else if (io_increment) begin
      state_12 <= state_11;
    end
    if (metaReset) begin
      state_13 <= 1'h0;
    end else if (reset) begin
      state_13 <= 1'h0;
    end else if (io_increment) begin
      state_13 <= state_12;
    end
    if (metaReset) begin
      state_14 <= 1'h0;
    end else if (reset) begin
      state_14 <= 1'h0;
    end else if (io_increment) begin
      state_14 <= state_13;
    end
    if (metaReset) begin
      state_15 <= 1'h0;
    end else if (reset) begin
      state_15 <= 1'h0;
    end else if (io_increment) begin
      state_15 <= state_14;
    end
  end
endmodule
module DCacheModuleImpl_Anon_1(
  input         io_in_0_valid,
  input  [39:0] io_in_0_bits_addr,
  input  [5:0]  io_in_0_bits_idx,
  input         io_in_1_valid,
  input  [39:0] io_in_1_bits_addr,
  input  [5:0]  io_in_1_bits_idx,
  input  [21:0] io_in_1_bits_data,
  input         io_in_2_valid,
  input  [39:0] io_in_2_bits_addr,
  input  [5:0]  io_in_2_bits_idx,
  input  [3:0]  io_in_2_bits_way_en,
  input  [21:0] io_in_2_bits_data,
  input         io_in_3_valid,
  input  [39:0] io_in_3_bits_addr,
  input  [5:0]  io_in_3_bits_idx,
  input  [3:0]  io_in_3_bits_way_en,
  input  [21:0] io_in_3_bits_data,
  output        io_in_4_ready,
  input         io_in_4_valid,
  input  [39:0] io_in_4_bits_addr,
  input  [5:0]  io_in_4_bits_idx,
  input  [3:0]  io_in_4_bits_way_en,
  input  [21:0] io_in_4_bits_data,
  output        io_in_5_ready,
  input         io_in_5_valid,
  input  [39:0] io_in_5_bits_addr,
  input  [5:0]  io_in_5_bits_idx,
  output        io_in_6_ready,
  input         io_in_6_valid,
  input  [39:0] io_in_6_bits_addr,
  input  [5:0]  io_in_6_bits_idx,
  input  [3:0]  io_in_6_bits_way_en,
  input  [21:0] io_in_6_bits_data,
  output        io_in_7_ready,
  input         io_in_7_valid,
  input  [39:0] io_in_7_bits_addr,
  input  [5:0]  io_in_7_bits_idx,
  input  [3:0]  io_in_7_bits_way_en,
  input  [21:0] io_in_7_bits_data,
  output        io_out_valid,
  output        io_out_bits_write,
  output [39:0] io_out_bits_addr,
  output [5:0]  io_out_bits_idx,
  output [3:0]  io_out_bits_way_en,
  output [21:0] io_out_bits_data,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire [21:0] _GEN_1; // @[Arbiter.scala 126:27]
  wire [3:0] _GEN_2; // @[Arbiter.scala 126:27]
  wire [5:0] _GEN_3; // @[Arbiter.scala 126:27]
  wire [39:0] _GEN_4; // @[Arbiter.scala 126:27]
  wire [21:0] _GEN_13; // @[Arbiter.scala 126:27]
  wire [3:0] _GEN_14; // @[Arbiter.scala 126:27]
  wire [5:0] _GEN_15; // @[Arbiter.scala 126:27]
  wire [39:0] _GEN_16; // @[Arbiter.scala 126:27]
  wire [21:0] _GEN_19; // @[Arbiter.scala 126:27]
  wire [3:0] _GEN_20; // @[Arbiter.scala 126:27]
  wire [5:0] _GEN_21; // @[Arbiter.scala 126:27]
  wire [39:0] _GEN_22; // @[Arbiter.scala 126:27]
  wire  _GEN_23; // @[Arbiter.scala 126:27]
  wire [21:0] _GEN_25; // @[Arbiter.scala 126:27]
  wire [3:0] _GEN_26; // @[Arbiter.scala 126:27]
  wire [5:0] _GEN_27; // @[Arbiter.scala 126:27]
  wire [39:0] _GEN_28; // @[Arbiter.scala 126:27]
  wire  _GEN_29; // @[Arbiter.scala 126:27]
  wire [21:0] _GEN_31; // @[Arbiter.scala 126:27]
  wire [3:0] _GEN_32; // @[Arbiter.scala 126:27]
  wire [5:0] _GEN_33; // @[Arbiter.scala 126:27]
  wire [39:0] _GEN_34; // @[Arbiter.scala 126:27]
  wire  _GEN_35; // @[Arbiter.scala 126:27]
  wire  _grant_T; // @[Arbiter.scala 31:68]
  wire  _grant_T_1; // @[Arbiter.scala 31:68]
  wire  _grant_T_2; // @[Arbiter.scala 31:68]
  wire  _grant_T_3; // @[Arbiter.scala 31:68]
  wire  _grant_T_5; // @[Arbiter.scala 31:68]
  wire  grant_7; // @[Arbiter.scala 31:78]
  wire [29:0] DCacheModuleImpl_Anon_1_covSum;
  assign _GEN_1 = io_in_6_valid ? io_in_6_bits_data : io_in_7_bits_data; // @[Arbiter.scala 126:27]
  assign _GEN_2 = io_in_6_valid ? io_in_6_bits_way_en : io_in_7_bits_way_en; // @[Arbiter.scala 126:27]
  assign _GEN_3 = io_in_6_valid ? io_in_6_bits_idx : io_in_7_bits_idx; // @[Arbiter.scala 126:27]
  assign _GEN_4 = io_in_6_valid ? io_in_6_bits_addr : io_in_7_bits_addr; // @[Arbiter.scala 126:27]
  assign _GEN_13 = io_in_4_valid ? io_in_4_bits_data : _GEN_1; // @[Arbiter.scala 126:27]
  assign _GEN_14 = io_in_4_valid ? io_in_4_bits_way_en : _GEN_2; // @[Arbiter.scala 126:27]
  assign _GEN_15 = io_in_4_valid ? io_in_4_bits_idx : _GEN_3; // @[Arbiter.scala 126:27]
  assign _GEN_16 = io_in_4_valid ? io_in_4_bits_addr : _GEN_4; // @[Arbiter.scala 126:27]
  assign _GEN_19 = io_in_3_valid ? io_in_3_bits_data : _GEN_13; // @[Arbiter.scala 126:27]
  assign _GEN_20 = io_in_3_valid ? io_in_3_bits_way_en : _GEN_14; // @[Arbiter.scala 126:27]
  assign _GEN_21 = io_in_3_valid ? io_in_3_bits_idx : _GEN_15; // @[Arbiter.scala 126:27]
  assign _GEN_22 = io_in_3_valid ? io_in_3_bits_addr : _GEN_16; // @[Arbiter.scala 126:27]
  assign _GEN_23 = io_in_3_valid | io_in_4_valid; // @[Arbiter.scala 126:27]
  assign _GEN_25 = io_in_2_valid ? io_in_2_bits_data : _GEN_19; // @[Arbiter.scala 126:27]
  assign _GEN_26 = io_in_2_valid ? io_in_2_bits_way_en : _GEN_20; // @[Arbiter.scala 126:27]
  assign _GEN_27 = io_in_2_valid ? io_in_2_bits_idx : _GEN_21; // @[Arbiter.scala 126:27]
  assign _GEN_28 = io_in_2_valid ? io_in_2_bits_addr : _GEN_22; // @[Arbiter.scala 126:27]
  assign _GEN_29 = io_in_2_valid | _GEN_23; // @[Arbiter.scala 126:27]
  assign _GEN_31 = io_in_1_valid ? io_in_1_bits_data : _GEN_25; // @[Arbiter.scala 126:27]
  assign _GEN_32 = io_in_1_valid ? 4'h0 : _GEN_26; // @[Arbiter.scala 126:27]
  assign _GEN_33 = io_in_1_valid ? io_in_1_bits_idx : _GEN_27; // @[Arbiter.scala 126:27]
  assign _GEN_34 = io_in_1_valid ? io_in_1_bits_addr : _GEN_28; // @[Arbiter.scala 126:27]
  assign _GEN_35 = io_in_1_valid | _GEN_29; // @[Arbiter.scala 126:27]
  assign _grant_T = io_in_0_valid | io_in_1_valid; // @[Arbiter.scala 31:68]
  assign _grant_T_1 = _grant_T | io_in_2_valid; // @[Arbiter.scala 31:68]
  assign _grant_T_2 = _grant_T_1 | io_in_3_valid; // @[Arbiter.scala 31:68]
  assign _grant_T_3 = _grant_T_2 | io_in_4_valid; // @[Arbiter.scala 31:68]
  assign _grant_T_5 = _grant_T_3 | io_in_6_valid; // @[Arbiter.scala 31:68]
  assign grant_7 = ~_grant_T_5; // @[Arbiter.scala 31:78]
  assign io_in_4_ready = ~_grant_T_2; // @[Arbiter.scala 134:14]
  assign io_in_5_ready = ~_grant_T_3; // @[Arbiter.scala 134:14]
  assign io_in_6_ready = ~_grant_T_3; // @[Arbiter.scala 134:14]
  assign io_in_7_ready = ~_grant_T_5; // @[Arbiter.scala 134:14]
  assign io_out_valid = ~grant_7 | io_in_7_valid; // @[Arbiter.scala 135:16]
  assign io_out_bits_write = io_in_0_valid | _GEN_35; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign io_out_bits_addr = io_in_0_valid ? io_in_0_bits_addr : _GEN_34; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign io_out_bits_idx = io_in_0_valid ? io_in_0_bits_idx : _GEN_33; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign io_out_bits_way_en = io_in_0_valid ? 4'hf : _GEN_32; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign io_out_bits_data = io_in_0_valid ? 22'h0 : _GEN_31; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign DCacheModuleImpl_Anon_1_covSum = 30'h0;
  assign io_covSum = DCacheModuleImpl_Anon_1_covSum;
  assign metaAssert = 1'h0;
endmodule
module DCacheDataArray(
  input         clock,
  input         io_req_valid,
  input  [11:0] io_req_bits_addr,
  input         io_req_bits_write,
  input  [63:0] io_req_bits_wdata,
  input  [7:0]  io_req_bits_eccMask,
  input  [3:0]  io_req_bits_way_en,
  output [63:0] io_resp_0,
  output [63:0] io_resp_1,
  output [63:0] io_resp_2,
  output [63:0] io_resp_3,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  reg [7:0] data_arrays_0_0 [0:511]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_0;
  wire [7:0] data_arrays_0_0_rdata_data_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_0_rdata_data_addr; // @[DescribedSRAM.scala 19:26]
  wire [7:0] data_arrays_0_0_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_0_rdata_MPORT_addr; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_0_rdata_MPORT_mask; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_0_rdata_MPORT_en; // @[DescribedSRAM.scala 19:26]
  reg  data_arrays_0_0_rdata_data_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [8:0] data_arrays_0_0_rdata_data_addr_pipe_0;
  reg [31:0] _RAND_2;
  reg [7:0] data_arrays_0_1 [0:511]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_3;
  wire [7:0] data_arrays_0_1_rdata_data_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_1_rdata_data_addr; // @[DescribedSRAM.scala 19:26]
  wire [7:0] data_arrays_0_1_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_1_rdata_MPORT_addr; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_1_rdata_MPORT_mask; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_1_rdata_MPORT_en; // @[DescribedSRAM.scala 19:26]
  reg  data_arrays_0_1_rdata_data_en_pipe_0;
  reg [31:0] _RAND_4;
  reg [8:0] data_arrays_0_1_rdata_data_addr_pipe_0;
  reg [31:0] _RAND_5;
  reg [7:0] data_arrays_0_2 [0:511]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_6;
  wire [7:0] data_arrays_0_2_rdata_data_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_2_rdata_data_addr; // @[DescribedSRAM.scala 19:26]
  wire [7:0] data_arrays_0_2_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_2_rdata_MPORT_addr; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_2_rdata_MPORT_mask; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_2_rdata_MPORT_en; // @[DescribedSRAM.scala 19:26]
  reg  data_arrays_0_2_rdata_data_en_pipe_0;
  reg [31:0] _RAND_7;
  reg [8:0] data_arrays_0_2_rdata_data_addr_pipe_0;
  reg [31:0] _RAND_8;
  reg [7:0] data_arrays_0_3 [0:511]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_9;
  wire [7:0] data_arrays_0_3_rdata_data_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_3_rdata_data_addr; // @[DescribedSRAM.scala 19:26]
  wire [7:0] data_arrays_0_3_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_3_rdata_MPORT_addr; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_3_rdata_MPORT_mask; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_3_rdata_MPORT_en; // @[DescribedSRAM.scala 19:26]
  reg  data_arrays_0_3_rdata_data_en_pipe_0;
  reg [31:0] _RAND_10;
  reg [8:0] data_arrays_0_3_rdata_data_addr_pipe_0;
  reg [31:0] _RAND_11;
  reg [7:0] data_arrays_0_4 [0:511]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_12;
  wire [7:0] data_arrays_0_4_rdata_data_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_4_rdata_data_addr; // @[DescribedSRAM.scala 19:26]
  wire [7:0] data_arrays_0_4_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_4_rdata_MPORT_addr; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_4_rdata_MPORT_mask; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_4_rdata_MPORT_en; // @[DescribedSRAM.scala 19:26]
  reg  data_arrays_0_4_rdata_data_en_pipe_0;
  reg [31:0] _RAND_13;
  reg [8:0] data_arrays_0_4_rdata_data_addr_pipe_0;
  reg [31:0] _RAND_14;
  reg [7:0] data_arrays_0_5 [0:511]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_15;
  wire [7:0] data_arrays_0_5_rdata_data_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_5_rdata_data_addr; // @[DescribedSRAM.scala 19:26]
  wire [7:0] data_arrays_0_5_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_5_rdata_MPORT_addr; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_5_rdata_MPORT_mask; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_5_rdata_MPORT_en; // @[DescribedSRAM.scala 19:26]
  reg  data_arrays_0_5_rdata_data_en_pipe_0;
  reg [31:0] _RAND_16;
  reg [8:0] data_arrays_0_5_rdata_data_addr_pipe_0;
  reg [31:0] _RAND_17;
  reg [7:0] data_arrays_0_6 [0:511]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_18;
  wire [7:0] data_arrays_0_6_rdata_data_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_6_rdata_data_addr; // @[DescribedSRAM.scala 19:26]
  wire [7:0] data_arrays_0_6_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_6_rdata_MPORT_addr; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_6_rdata_MPORT_mask; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_6_rdata_MPORT_en; // @[DescribedSRAM.scala 19:26]
  reg  data_arrays_0_6_rdata_data_en_pipe_0;
  reg [31:0] _RAND_19;
  reg [8:0] data_arrays_0_6_rdata_data_addr_pipe_0;
  reg [31:0] _RAND_20;
  reg [7:0] data_arrays_0_7 [0:511]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_21;
  wire [7:0] data_arrays_0_7_rdata_data_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_7_rdata_data_addr; // @[DescribedSRAM.scala 19:26]
  wire [7:0] data_arrays_0_7_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_7_rdata_MPORT_addr; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_7_rdata_MPORT_mask; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_7_rdata_MPORT_en; // @[DescribedSRAM.scala 19:26]
  reg  data_arrays_0_7_rdata_data_en_pipe_0;
  reg [31:0] _RAND_22;
  reg [8:0] data_arrays_0_7_rdata_data_addr_pipe_0;
  reg [31:0] _RAND_23;
  reg [7:0] data_arrays_0_8 [0:511]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_24;
  wire [7:0] data_arrays_0_8_rdata_data_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_8_rdata_data_addr; // @[DescribedSRAM.scala 19:26]
  wire [7:0] data_arrays_0_8_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_8_rdata_MPORT_addr; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_8_rdata_MPORT_mask; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_8_rdata_MPORT_en; // @[DescribedSRAM.scala 19:26]
  reg  data_arrays_0_8_rdata_data_en_pipe_0;
  reg [31:0] _RAND_25;
  reg [8:0] data_arrays_0_8_rdata_data_addr_pipe_0;
  reg [31:0] _RAND_26;
  reg [7:0] data_arrays_0_9 [0:511]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_27;
  wire [7:0] data_arrays_0_9_rdata_data_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_9_rdata_data_addr; // @[DescribedSRAM.scala 19:26]
  wire [7:0] data_arrays_0_9_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_9_rdata_MPORT_addr; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_9_rdata_MPORT_mask; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_9_rdata_MPORT_en; // @[DescribedSRAM.scala 19:26]
  reg  data_arrays_0_9_rdata_data_en_pipe_0;
  reg [31:0] _RAND_28;
  reg [8:0] data_arrays_0_9_rdata_data_addr_pipe_0;
  reg [31:0] _RAND_29;
  reg [7:0] data_arrays_0_10 [0:511]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_30;
  wire [7:0] data_arrays_0_10_rdata_data_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_10_rdata_data_addr; // @[DescribedSRAM.scala 19:26]
  wire [7:0] data_arrays_0_10_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_10_rdata_MPORT_addr; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_10_rdata_MPORT_mask; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_10_rdata_MPORT_en; // @[DescribedSRAM.scala 19:26]
  reg  data_arrays_0_10_rdata_data_en_pipe_0;
  reg [31:0] _RAND_31;
  reg [8:0] data_arrays_0_10_rdata_data_addr_pipe_0;
  reg [31:0] _RAND_32;
  reg [7:0] data_arrays_0_11 [0:511]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_33;
  wire [7:0] data_arrays_0_11_rdata_data_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_11_rdata_data_addr; // @[DescribedSRAM.scala 19:26]
  wire [7:0] data_arrays_0_11_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_11_rdata_MPORT_addr; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_11_rdata_MPORT_mask; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_11_rdata_MPORT_en; // @[DescribedSRAM.scala 19:26]
  reg  data_arrays_0_11_rdata_data_en_pipe_0;
  reg [31:0] _RAND_34;
  reg [8:0] data_arrays_0_11_rdata_data_addr_pipe_0;
  reg [31:0] _RAND_35;
  reg [7:0] data_arrays_0_12 [0:511]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_36;
  wire [7:0] data_arrays_0_12_rdata_data_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_12_rdata_data_addr; // @[DescribedSRAM.scala 19:26]
  wire [7:0] data_arrays_0_12_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_12_rdata_MPORT_addr; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_12_rdata_MPORT_mask; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_12_rdata_MPORT_en; // @[DescribedSRAM.scala 19:26]
  reg  data_arrays_0_12_rdata_data_en_pipe_0;
  reg [31:0] _RAND_37;
  reg [8:0] data_arrays_0_12_rdata_data_addr_pipe_0;
  reg [31:0] _RAND_38;
  reg [7:0] data_arrays_0_13 [0:511]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_39;
  wire [7:0] data_arrays_0_13_rdata_data_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_13_rdata_data_addr; // @[DescribedSRAM.scala 19:26]
  wire [7:0] data_arrays_0_13_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_13_rdata_MPORT_addr; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_13_rdata_MPORT_mask; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_13_rdata_MPORT_en; // @[DescribedSRAM.scala 19:26]
  reg  data_arrays_0_13_rdata_data_en_pipe_0;
  reg [31:0] _RAND_40;
  reg [8:0] data_arrays_0_13_rdata_data_addr_pipe_0;
  reg [31:0] _RAND_41;
  reg [7:0] data_arrays_0_14 [0:511]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_42;
  wire [7:0] data_arrays_0_14_rdata_data_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_14_rdata_data_addr; // @[DescribedSRAM.scala 19:26]
  wire [7:0] data_arrays_0_14_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_14_rdata_MPORT_addr; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_14_rdata_MPORT_mask; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_14_rdata_MPORT_en; // @[DescribedSRAM.scala 19:26]
  reg  data_arrays_0_14_rdata_data_en_pipe_0;
  reg [31:0] _RAND_43;
  reg [8:0] data_arrays_0_14_rdata_data_addr_pipe_0;
  reg [31:0] _RAND_44;
  reg [7:0] data_arrays_0_15 [0:511]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_45;
  wire [7:0] data_arrays_0_15_rdata_data_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_15_rdata_data_addr; // @[DescribedSRAM.scala 19:26]
  wire [7:0] data_arrays_0_15_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_15_rdata_MPORT_addr; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_15_rdata_MPORT_mask; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_15_rdata_MPORT_en; // @[DescribedSRAM.scala 19:26]
  reg  data_arrays_0_15_rdata_data_en_pipe_0;
  reg [31:0] _RAND_46;
  reg [8:0] data_arrays_0_15_rdata_data_addr_pipe_0;
  reg [31:0] _RAND_47;
  reg [7:0] data_arrays_0_16 [0:511]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_48;
  wire [7:0] data_arrays_0_16_rdata_data_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_16_rdata_data_addr; // @[DescribedSRAM.scala 19:26]
  wire [7:0] data_arrays_0_16_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_16_rdata_MPORT_addr; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_16_rdata_MPORT_mask; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_16_rdata_MPORT_en; // @[DescribedSRAM.scala 19:26]
  reg  data_arrays_0_16_rdata_data_en_pipe_0;
  reg [31:0] _RAND_49;
  reg [8:0] data_arrays_0_16_rdata_data_addr_pipe_0;
  reg [31:0] _RAND_50;
  reg [7:0] data_arrays_0_17 [0:511]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_51;
  wire [7:0] data_arrays_0_17_rdata_data_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_17_rdata_data_addr; // @[DescribedSRAM.scala 19:26]
  wire [7:0] data_arrays_0_17_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_17_rdata_MPORT_addr; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_17_rdata_MPORT_mask; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_17_rdata_MPORT_en; // @[DescribedSRAM.scala 19:26]
  reg  data_arrays_0_17_rdata_data_en_pipe_0;
  reg [31:0] _RAND_52;
  reg [8:0] data_arrays_0_17_rdata_data_addr_pipe_0;
  reg [31:0] _RAND_53;
  reg [7:0] data_arrays_0_18 [0:511]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_54;
  wire [7:0] data_arrays_0_18_rdata_data_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_18_rdata_data_addr; // @[DescribedSRAM.scala 19:26]
  wire [7:0] data_arrays_0_18_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_18_rdata_MPORT_addr; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_18_rdata_MPORT_mask; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_18_rdata_MPORT_en; // @[DescribedSRAM.scala 19:26]
  reg  data_arrays_0_18_rdata_data_en_pipe_0;
  reg [31:0] _RAND_55;
  reg [8:0] data_arrays_0_18_rdata_data_addr_pipe_0;
  reg [31:0] _RAND_56;
  reg [7:0] data_arrays_0_19 [0:511]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_57;
  wire [7:0] data_arrays_0_19_rdata_data_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_19_rdata_data_addr; // @[DescribedSRAM.scala 19:26]
  wire [7:0] data_arrays_0_19_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_19_rdata_MPORT_addr; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_19_rdata_MPORT_mask; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_19_rdata_MPORT_en; // @[DescribedSRAM.scala 19:26]
  reg  data_arrays_0_19_rdata_data_en_pipe_0;
  reg [31:0] _RAND_58;
  reg [8:0] data_arrays_0_19_rdata_data_addr_pipe_0;
  reg [31:0] _RAND_59;
  reg [7:0] data_arrays_0_20 [0:511]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_60;
  wire [7:0] data_arrays_0_20_rdata_data_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_20_rdata_data_addr; // @[DescribedSRAM.scala 19:26]
  wire [7:0] data_arrays_0_20_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_20_rdata_MPORT_addr; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_20_rdata_MPORT_mask; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_20_rdata_MPORT_en; // @[DescribedSRAM.scala 19:26]
  reg  data_arrays_0_20_rdata_data_en_pipe_0;
  reg [31:0] _RAND_61;
  reg [8:0] data_arrays_0_20_rdata_data_addr_pipe_0;
  reg [31:0] _RAND_62;
  reg [7:0] data_arrays_0_21 [0:511]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_63;
  wire [7:0] data_arrays_0_21_rdata_data_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_21_rdata_data_addr; // @[DescribedSRAM.scala 19:26]
  wire [7:0] data_arrays_0_21_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_21_rdata_MPORT_addr; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_21_rdata_MPORT_mask; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_21_rdata_MPORT_en; // @[DescribedSRAM.scala 19:26]
  reg  data_arrays_0_21_rdata_data_en_pipe_0;
  reg [31:0] _RAND_64;
  reg [8:0] data_arrays_0_21_rdata_data_addr_pipe_0;
  reg [31:0] _RAND_65;
  reg [7:0] data_arrays_0_22 [0:511]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_66;
  wire [7:0] data_arrays_0_22_rdata_data_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_22_rdata_data_addr; // @[DescribedSRAM.scala 19:26]
  wire [7:0] data_arrays_0_22_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_22_rdata_MPORT_addr; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_22_rdata_MPORT_mask; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_22_rdata_MPORT_en; // @[DescribedSRAM.scala 19:26]
  reg  data_arrays_0_22_rdata_data_en_pipe_0;
  reg [31:0] _RAND_67;
  reg [8:0] data_arrays_0_22_rdata_data_addr_pipe_0;
  reg [31:0] _RAND_68;
  reg [7:0] data_arrays_0_23 [0:511]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_69;
  wire [7:0] data_arrays_0_23_rdata_data_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_23_rdata_data_addr; // @[DescribedSRAM.scala 19:26]
  wire [7:0] data_arrays_0_23_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_23_rdata_MPORT_addr; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_23_rdata_MPORT_mask; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_23_rdata_MPORT_en; // @[DescribedSRAM.scala 19:26]
  reg  data_arrays_0_23_rdata_data_en_pipe_0;
  reg [31:0] _RAND_70;
  reg [8:0] data_arrays_0_23_rdata_data_addr_pipe_0;
  reg [31:0] _RAND_71;
  reg [7:0] data_arrays_0_24 [0:511]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_72;
  wire [7:0] data_arrays_0_24_rdata_data_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_24_rdata_data_addr; // @[DescribedSRAM.scala 19:26]
  wire [7:0] data_arrays_0_24_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_24_rdata_MPORT_addr; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_24_rdata_MPORT_mask; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_24_rdata_MPORT_en; // @[DescribedSRAM.scala 19:26]
  reg  data_arrays_0_24_rdata_data_en_pipe_0;
  reg [31:0] _RAND_73;
  reg [8:0] data_arrays_0_24_rdata_data_addr_pipe_0;
  reg [31:0] _RAND_74;
  reg [7:0] data_arrays_0_25 [0:511]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_75;
  wire [7:0] data_arrays_0_25_rdata_data_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_25_rdata_data_addr; // @[DescribedSRAM.scala 19:26]
  wire [7:0] data_arrays_0_25_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_25_rdata_MPORT_addr; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_25_rdata_MPORT_mask; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_25_rdata_MPORT_en; // @[DescribedSRAM.scala 19:26]
  reg  data_arrays_0_25_rdata_data_en_pipe_0;
  reg [31:0] _RAND_76;
  reg [8:0] data_arrays_0_25_rdata_data_addr_pipe_0;
  reg [31:0] _RAND_77;
  reg [7:0] data_arrays_0_26 [0:511]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_78;
  wire [7:0] data_arrays_0_26_rdata_data_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_26_rdata_data_addr; // @[DescribedSRAM.scala 19:26]
  wire [7:0] data_arrays_0_26_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_26_rdata_MPORT_addr; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_26_rdata_MPORT_mask; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_26_rdata_MPORT_en; // @[DescribedSRAM.scala 19:26]
  reg  data_arrays_0_26_rdata_data_en_pipe_0;
  reg [31:0] _RAND_79;
  reg [8:0] data_arrays_0_26_rdata_data_addr_pipe_0;
  reg [31:0] _RAND_80;
  reg [7:0] data_arrays_0_27 [0:511]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_81;
  wire [7:0] data_arrays_0_27_rdata_data_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_27_rdata_data_addr; // @[DescribedSRAM.scala 19:26]
  wire [7:0] data_arrays_0_27_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_27_rdata_MPORT_addr; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_27_rdata_MPORT_mask; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_27_rdata_MPORT_en; // @[DescribedSRAM.scala 19:26]
  reg  data_arrays_0_27_rdata_data_en_pipe_0;
  reg [31:0] _RAND_82;
  reg [8:0] data_arrays_0_27_rdata_data_addr_pipe_0;
  reg [31:0] _RAND_83;
  reg [7:0] data_arrays_0_28 [0:511]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_84;
  wire [7:0] data_arrays_0_28_rdata_data_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_28_rdata_data_addr; // @[DescribedSRAM.scala 19:26]
  wire [7:0] data_arrays_0_28_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_28_rdata_MPORT_addr; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_28_rdata_MPORT_mask; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_28_rdata_MPORT_en; // @[DescribedSRAM.scala 19:26]
  reg  data_arrays_0_28_rdata_data_en_pipe_0;
  reg [31:0] _RAND_85;
  reg [8:0] data_arrays_0_28_rdata_data_addr_pipe_0;
  reg [31:0] _RAND_86;
  reg [7:0] data_arrays_0_29 [0:511]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_87;
  wire [7:0] data_arrays_0_29_rdata_data_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_29_rdata_data_addr; // @[DescribedSRAM.scala 19:26]
  wire [7:0] data_arrays_0_29_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_29_rdata_MPORT_addr; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_29_rdata_MPORT_mask; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_29_rdata_MPORT_en; // @[DescribedSRAM.scala 19:26]
  reg  data_arrays_0_29_rdata_data_en_pipe_0;
  reg [31:0] _RAND_88;
  reg [8:0] data_arrays_0_29_rdata_data_addr_pipe_0;
  reg [31:0] _RAND_89;
  reg [7:0] data_arrays_0_30 [0:511]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_90;
  wire [7:0] data_arrays_0_30_rdata_data_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_30_rdata_data_addr; // @[DescribedSRAM.scala 19:26]
  wire [7:0] data_arrays_0_30_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_30_rdata_MPORT_addr; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_30_rdata_MPORT_mask; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_30_rdata_MPORT_en; // @[DescribedSRAM.scala 19:26]
  reg  data_arrays_0_30_rdata_data_en_pipe_0;
  reg [31:0] _RAND_91;
  reg [8:0] data_arrays_0_30_rdata_data_addr_pipe_0;
  reg [31:0] _RAND_92;
  reg [7:0] data_arrays_0_31 [0:511]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_93;
  wire [7:0] data_arrays_0_31_rdata_data_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_31_rdata_data_addr; // @[DescribedSRAM.scala 19:26]
  wire [7:0] data_arrays_0_31_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_31_rdata_MPORT_addr; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_31_rdata_MPORT_mask; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_31_rdata_MPORT_en; // @[DescribedSRAM.scala 19:26]
  reg  data_arrays_0_31_rdata_data_en_pipe_0;
  reg [31:0] _RAND_94;
  reg [8:0] data_arrays_0_31_rdata_data_addr_pipe_0;
  reg [31:0] _RAND_95;
  wire  eccMask_0; // @[DCache.scala 50:82]
  wire  eccMask_1; // @[DCache.scala 50:82]
  wire  eccMask_2; // @[DCache.scala 50:82]
  wire  eccMask_3; // @[DCache.scala 50:82]
  wire  eccMask_4; // @[DCache.scala 50:82]
  wire  eccMask_5; // @[DCache.scala 50:82]
  wire  eccMask_6; // @[DCache.scala 50:82]
  wire  eccMask_7; // @[DCache.scala 50:82]
  wire [31:0] rdata_lo; // @[Cat.scala 30:58]
  wire [31:0] rdata_hi; // @[Cat.scala 30:58]
  wire [31:0] lo; // @[Cat.scala 30:58]
  wire [31:0] hi; // @[Cat.scala 30:58]
  wire [31:0] lo_1; // @[Cat.scala 30:58]
  wire [31:0] hi_1; // @[Cat.scala 30:58]
  wire [31:0] lo_2; // @[Cat.scala 30:58]
  wire [31:0] hi_2; // @[Cat.scala 30:58]
  wire [29:0] DCacheDataArray_covSum;
  assign data_arrays_0_0_rdata_data_addr = data_arrays_0_0_rdata_data_addr_pipe_0;
  assign data_arrays_0_0_rdata_data_data = data_arrays_0_0[data_arrays_0_0_rdata_data_addr]; // @[DescribedSRAM.scala 19:26]
  assign data_arrays_0_0_rdata_MPORT_data = io_req_bits_wdata[7:0];
  assign data_arrays_0_0_rdata_MPORT_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_0_rdata_MPORT_mask = eccMask_0 & io_req_bits_way_en[0];
  assign data_arrays_0_0_rdata_MPORT_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_1_rdata_data_addr = data_arrays_0_1_rdata_data_addr_pipe_0;
  assign data_arrays_0_1_rdata_data_data = data_arrays_0_1[data_arrays_0_1_rdata_data_addr]; // @[DescribedSRAM.scala 19:26]
  assign data_arrays_0_1_rdata_MPORT_data = io_req_bits_wdata[15:8];
  assign data_arrays_0_1_rdata_MPORT_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_1_rdata_MPORT_mask = eccMask_1 & io_req_bits_way_en[0];
  assign data_arrays_0_1_rdata_MPORT_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_2_rdata_data_addr = data_arrays_0_2_rdata_data_addr_pipe_0;
  assign data_arrays_0_2_rdata_data_data = data_arrays_0_2[data_arrays_0_2_rdata_data_addr]; // @[DescribedSRAM.scala 19:26]
  assign data_arrays_0_2_rdata_MPORT_data = io_req_bits_wdata[23:16];
  assign data_arrays_0_2_rdata_MPORT_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_2_rdata_MPORT_mask = eccMask_2 & io_req_bits_way_en[0];
  assign data_arrays_0_2_rdata_MPORT_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_3_rdata_data_addr = data_arrays_0_3_rdata_data_addr_pipe_0;
  assign data_arrays_0_3_rdata_data_data = data_arrays_0_3[data_arrays_0_3_rdata_data_addr]; // @[DescribedSRAM.scala 19:26]
  assign data_arrays_0_3_rdata_MPORT_data = io_req_bits_wdata[31:24];
  assign data_arrays_0_3_rdata_MPORT_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_3_rdata_MPORT_mask = eccMask_3 & io_req_bits_way_en[0];
  assign data_arrays_0_3_rdata_MPORT_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_4_rdata_data_addr = data_arrays_0_4_rdata_data_addr_pipe_0;
  assign data_arrays_0_4_rdata_data_data = data_arrays_0_4[data_arrays_0_4_rdata_data_addr]; // @[DescribedSRAM.scala 19:26]
  assign data_arrays_0_4_rdata_MPORT_data = io_req_bits_wdata[39:32];
  assign data_arrays_0_4_rdata_MPORT_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_4_rdata_MPORT_mask = eccMask_4 & io_req_bits_way_en[0];
  assign data_arrays_0_4_rdata_MPORT_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_5_rdata_data_addr = data_arrays_0_5_rdata_data_addr_pipe_0;
  assign data_arrays_0_5_rdata_data_data = data_arrays_0_5[data_arrays_0_5_rdata_data_addr]; // @[DescribedSRAM.scala 19:26]
  assign data_arrays_0_5_rdata_MPORT_data = io_req_bits_wdata[47:40];
  assign data_arrays_0_5_rdata_MPORT_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_5_rdata_MPORT_mask = eccMask_5 & io_req_bits_way_en[0];
  assign data_arrays_0_5_rdata_MPORT_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_6_rdata_data_addr = data_arrays_0_6_rdata_data_addr_pipe_0;
  assign data_arrays_0_6_rdata_data_data = data_arrays_0_6[data_arrays_0_6_rdata_data_addr]; // @[DescribedSRAM.scala 19:26]
  assign data_arrays_0_6_rdata_MPORT_data = io_req_bits_wdata[55:48];
  assign data_arrays_0_6_rdata_MPORT_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_6_rdata_MPORT_mask = eccMask_6 & io_req_bits_way_en[0];
  assign data_arrays_0_6_rdata_MPORT_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_7_rdata_data_addr = data_arrays_0_7_rdata_data_addr_pipe_0;
  assign data_arrays_0_7_rdata_data_data = data_arrays_0_7[data_arrays_0_7_rdata_data_addr]; // @[DescribedSRAM.scala 19:26]
  assign data_arrays_0_7_rdata_MPORT_data = io_req_bits_wdata[63:56];
  assign data_arrays_0_7_rdata_MPORT_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_7_rdata_MPORT_mask = eccMask_7 & io_req_bits_way_en[0];
  assign data_arrays_0_7_rdata_MPORT_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_8_rdata_data_addr = data_arrays_0_8_rdata_data_addr_pipe_0;
  assign data_arrays_0_8_rdata_data_data = data_arrays_0_8[data_arrays_0_8_rdata_data_addr]; // @[DescribedSRAM.scala 19:26]
  assign data_arrays_0_8_rdata_MPORT_data = io_req_bits_wdata[7:0];
  assign data_arrays_0_8_rdata_MPORT_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_8_rdata_MPORT_mask = eccMask_0 & io_req_bits_way_en[1];
  assign data_arrays_0_8_rdata_MPORT_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_9_rdata_data_addr = data_arrays_0_9_rdata_data_addr_pipe_0;
  assign data_arrays_0_9_rdata_data_data = data_arrays_0_9[data_arrays_0_9_rdata_data_addr]; // @[DescribedSRAM.scala 19:26]
  assign data_arrays_0_9_rdata_MPORT_data = io_req_bits_wdata[15:8];
  assign data_arrays_0_9_rdata_MPORT_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_9_rdata_MPORT_mask = eccMask_1 & io_req_bits_way_en[1];
  assign data_arrays_0_9_rdata_MPORT_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_10_rdata_data_addr = data_arrays_0_10_rdata_data_addr_pipe_0;
  assign data_arrays_0_10_rdata_data_data = data_arrays_0_10[data_arrays_0_10_rdata_data_addr]; // @[DescribedSRAM.scala 19:26]
  assign data_arrays_0_10_rdata_MPORT_data = io_req_bits_wdata[23:16];
  assign data_arrays_0_10_rdata_MPORT_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_10_rdata_MPORT_mask = eccMask_2 & io_req_bits_way_en[1];
  assign data_arrays_0_10_rdata_MPORT_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_11_rdata_data_addr = data_arrays_0_11_rdata_data_addr_pipe_0;
  assign data_arrays_0_11_rdata_data_data = data_arrays_0_11[data_arrays_0_11_rdata_data_addr]; // @[DescribedSRAM.scala 19:26]
  assign data_arrays_0_11_rdata_MPORT_data = io_req_bits_wdata[31:24];
  assign data_arrays_0_11_rdata_MPORT_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_11_rdata_MPORT_mask = eccMask_3 & io_req_bits_way_en[1];
  assign data_arrays_0_11_rdata_MPORT_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_12_rdata_data_addr = data_arrays_0_12_rdata_data_addr_pipe_0;
  assign data_arrays_0_12_rdata_data_data = data_arrays_0_12[data_arrays_0_12_rdata_data_addr]; // @[DescribedSRAM.scala 19:26]
  assign data_arrays_0_12_rdata_MPORT_data = io_req_bits_wdata[39:32];
  assign data_arrays_0_12_rdata_MPORT_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_12_rdata_MPORT_mask = eccMask_4 & io_req_bits_way_en[1];
  assign data_arrays_0_12_rdata_MPORT_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_13_rdata_data_addr = data_arrays_0_13_rdata_data_addr_pipe_0;
  assign data_arrays_0_13_rdata_data_data = data_arrays_0_13[data_arrays_0_13_rdata_data_addr]; // @[DescribedSRAM.scala 19:26]
  assign data_arrays_0_13_rdata_MPORT_data = io_req_bits_wdata[47:40];
  assign data_arrays_0_13_rdata_MPORT_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_13_rdata_MPORT_mask = eccMask_5 & io_req_bits_way_en[1];
  assign data_arrays_0_13_rdata_MPORT_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_14_rdata_data_addr = data_arrays_0_14_rdata_data_addr_pipe_0;
  assign data_arrays_0_14_rdata_data_data = data_arrays_0_14[data_arrays_0_14_rdata_data_addr]; // @[DescribedSRAM.scala 19:26]
  assign data_arrays_0_14_rdata_MPORT_data = io_req_bits_wdata[55:48];
  assign data_arrays_0_14_rdata_MPORT_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_14_rdata_MPORT_mask = eccMask_6 & io_req_bits_way_en[1];
  assign data_arrays_0_14_rdata_MPORT_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_15_rdata_data_addr = data_arrays_0_15_rdata_data_addr_pipe_0;
  assign data_arrays_0_15_rdata_data_data = data_arrays_0_15[data_arrays_0_15_rdata_data_addr]; // @[DescribedSRAM.scala 19:26]
  assign data_arrays_0_15_rdata_MPORT_data = io_req_bits_wdata[63:56];
  assign data_arrays_0_15_rdata_MPORT_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_15_rdata_MPORT_mask = eccMask_7 & io_req_bits_way_en[1];
  assign data_arrays_0_15_rdata_MPORT_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_16_rdata_data_addr = data_arrays_0_16_rdata_data_addr_pipe_0;
  assign data_arrays_0_16_rdata_data_data = data_arrays_0_16[data_arrays_0_16_rdata_data_addr]; // @[DescribedSRAM.scala 19:26]
  assign data_arrays_0_16_rdata_MPORT_data = io_req_bits_wdata[7:0];
  assign data_arrays_0_16_rdata_MPORT_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_16_rdata_MPORT_mask = eccMask_0 & io_req_bits_way_en[2];
  assign data_arrays_0_16_rdata_MPORT_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_17_rdata_data_addr = data_arrays_0_17_rdata_data_addr_pipe_0;
  assign data_arrays_0_17_rdata_data_data = data_arrays_0_17[data_arrays_0_17_rdata_data_addr]; // @[DescribedSRAM.scala 19:26]
  assign data_arrays_0_17_rdata_MPORT_data = io_req_bits_wdata[15:8];
  assign data_arrays_0_17_rdata_MPORT_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_17_rdata_MPORT_mask = eccMask_1 & io_req_bits_way_en[2];
  assign data_arrays_0_17_rdata_MPORT_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_18_rdata_data_addr = data_arrays_0_18_rdata_data_addr_pipe_0;
  assign data_arrays_0_18_rdata_data_data = data_arrays_0_18[data_arrays_0_18_rdata_data_addr]; // @[DescribedSRAM.scala 19:26]
  assign data_arrays_0_18_rdata_MPORT_data = io_req_bits_wdata[23:16];
  assign data_arrays_0_18_rdata_MPORT_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_18_rdata_MPORT_mask = eccMask_2 & io_req_bits_way_en[2];
  assign data_arrays_0_18_rdata_MPORT_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_19_rdata_data_addr = data_arrays_0_19_rdata_data_addr_pipe_0;
  assign data_arrays_0_19_rdata_data_data = data_arrays_0_19[data_arrays_0_19_rdata_data_addr]; // @[DescribedSRAM.scala 19:26]
  assign data_arrays_0_19_rdata_MPORT_data = io_req_bits_wdata[31:24];
  assign data_arrays_0_19_rdata_MPORT_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_19_rdata_MPORT_mask = eccMask_3 & io_req_bits_way_en[2];
  assign data_arrays_0_19_rdata_MPORT_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_20_rdata_data_addr = data_arrays_0_20_rdata_data_addr_pipe_0;
  assign data_arrays_0_20_rdata_data_data = data_arrays_0_20[data_arrays_0_20_rdata_data_addr]; // @[DescribedSRAM.scala 19:26]
  assign data_arrays_0_20_rdata_MPORT_data = io_req_bits_wdata[39:32];
  assign data_arrays_0_20_rdata_MPORT_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_20_rdata_MPORT_mask = eccMask_4 & io_req_bits_way_en[2];
  assign data_arrays_0_20_rdata_MPORT_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_21_rdata_data_addr = data_arrays_0_21_rdata_data_addr_pipe_0;
  assign data_arrays_0_21_rdata_data_data = data_arrays_0_21[data_arrays_0_21_rdata_data_addr]; // @[DescribedSRAM.scala 19:26]
  assign data_arrays_0_21_rdata_MPORT_data = io_req_bits_wdata[47:40];
  assign data_arrays_0_21_rdata_MPORT_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_21_rdata_MPORT_mask = eccMask_5 & io_req_bits_way_en[2];
  assign data_arrays_0_21_rdata_MPORT_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_22_rdata_data_addr = data_arrays_0_22_rdata_data_addr_pipe_0;
  assign data_arrays_0_22_rdata_data_data = data_arrays_0_22[data_arrays_0_22_rdata_data_addr]; // @[DescribedSRAM.scala 19:26]
  assign data_arrays_0_22_rdata_MPORT_data = io_req_bits_wdata[55:48];
  assign data_arrays_0_22_rdata_MPORT_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_22_rdata_MPORT_mask = eccMask_6 & io_req_bits_way_en[2];
  assign data_arrays_0_22_rdata_MPORT_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_23_rdata_data_addr = data_arrays_0_23_rdata_data_addr_pipe_0;
  assign data_arrays_0_23_rdata_data_data = data_arrays_0_23[data_arrays_0_23_rdata_data_addr]; // @[DescribedSRAM.scala 19:26]
  assign data_arrays_0_23_rdata_MPORT_data = io_req_bits_wdata[63:56];
  assign data_arrays_0_23_rdata_MPORT_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_23_rdata_MPORT_mask = eccMask_7 & io_req_bits_way_en[2];
  assign data_arrays_0_23_rdata_MPORT_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_24_rdata_data_addr = data_arrays_0_24_rdata_data_addr_pipe_0;
  assign data_arrays_0_24_rdata_data_data = data_arrays_0_24[data_arrays_0_24_rdata_data_addr]; // @[DescribedSRAM.scala 19:26]
  assign data_arrays_0_24_rdata_MPORT_data = io_req_bits_wdata[7:0];
  assign data_arrays_0_24_rdata_MPORT_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_24_rdata_MPORT_mask = eccMask_0 & io_req_bits_way_en[3];
  assign data_arrays_0_24_rdata_MPORT_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_25_rdata_data_addr = data_arrays_0_25_rdata_data_addr_pipe_0;
  assign data_arrays_0_25_rdata_data_data = data_arrays_0_25[data_arrays_0_25_rdata_data_addr]; // @[DescribedSRAM.scala 19:26]
  assign data_arrays_0_25_rdata_MPORT_data = io_req_bits_wdata[15:8];
  assign data_arrays_0_25_rdata_MPORT_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_25_rdata_MPORT_mask = eccMask_1 & io_req_bits_way_en[3];
  assign data_arrays_0_25_rdata_MPORT_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_26_rdata_data_addr = data_arrays_0_26_rdata_data_addr_pipe_0;
  assign data_arrays_0_26_rdata_data_data = data_arrays_0_26[data_arrays_0_26_rdata_data_addr]; // @[DescribedSRAM.scala 19:26]
  assign data_arrays_0_26_rdata_MPORT_data = io_req_bits_wdata[23:16];
  assign data_arrays_0_26_rdata_MPORT_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_26_rdata_MPORT_mask = eccMask_2 & io_req_bits_way_en[3];
  assign data_arrays_0_26_rdata_MPORT_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_27_rdata_data_addr = data_arrays_0_27_rdata_data_addr_pipe_0;
  assign data_arrays_0_27_rdata_data_data = data_arrays_0_27[data_arrays_0_27_rdata_data_addr]; // @[DescribedSRAM.scala 19:26]
  assign data_arrays_0_27_rdata_MPORT_data = io_req_bits_wdata[31:24];
  assign data_arrays_0_27_rdata_MPORT_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_27_rdata_MPORT_mask = eccMask_3 & io_req_bits_way_en[3];
  assign data_arrays_0_27_rdata_MPORT_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_28_rdata_data_addr = data_arrays_0_28_rdata_data_addr_pipe_0;
  assign data_arrays_0_28_rdata_data_data = data_arrays_0_28[data_arrays_0_28_rdata_data_addr]; // @[DescribedSRAM.scala 19:26]
  assign data_arrays_0_28_rdata_MPORT_data = io_req_bits_wdata[39:32];
  assign data_arrays_0_28_rdata_MPORT_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_28_rdata_MPORT_mask = eccMask_4 & io_req_bits_way_en[3];
  assign data_arrays_0_28_rdata_MPORT_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_29_rdata_data_addr = data_arrays_0_29_rdata_data_addr_pipe_0;
  assign data_arrays_0_29_rdata_data_data = data_arrays_0_29[data_arrays_0_29_rdata_data_addr]; // @[DescribedSRAM.scala 19:26]
  assign data_arrays_0_29_rdata_MPORT_data = io_req_bits_wdata[47:40];
  assign data_arrays_0_29_rdata_MPORT_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_29_rdata_MPORT_mask = eccMask_5 & io_req_bits_way_en[3];
  assign data_arrays_0_29_rdata_MPORT_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_30_rdata_data_addr = data_arrays_0_30_rdata_data_addr_pipe_0;
  assign data_arrays_0_30_rdata_data_data = data_arrays_0_30[data_arrays_0_30_rdata_data_addr]; // @[DescribedSRAM.scala 19:26]
  assign data_arrays_0_30_rdata_MPORT_data = io_req_bits_wdata[55:48];
  assign data_arrays_0_30_rdata_MPORT_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_30_rdata_MPORT_mask = eccMask_6 & io_req_bits_way_en[3];
  assign data_arrays_0_30_rdata_MPORT_en = io_req_valid & io_req_bits_write;
  assign data_arrays_0_31_rdata_data_addr = data_arrays_0_31_rdata_data_addr_pipe_0;
  assign data_arrays_0_31_rdata_data_data = data_arrays_0_31[data_arrays_0_31_rdata_data_addr]; // @[DescribedSRAM.scala 19:26]
  assign data_arrays_0_31_rdata_MPORT_data = io_req_bits_wdata[63:56];
  assign data_arrays_0_31_rdata_MPORT_addr = io_req_bits_addr[11:3];
  assign data_arrays_0_31_rdata_MPORT_mask = eccMask_7 & io_req_bits_way_en[3];
  assign data_arrays_0_31_rdata_MPORT_en = io_req_valid & io_req_bits_write;
  assign eccMask_0 = io_req_bits_eccMask[0]; // @[DCache.scala 50:82]
  assign eccMask_1 = io_req_bits_eccMask[1]; // @[DCache.scala 50:82]
  assign eccMask_2 = io_req_bits_eccMask[2]; // @[DCache.scala 50:82]
  assign eccMask_3 = io_req_bits_eccMask[3]; // @[DCache.scala 50:82]
  assign eccMask_4 = io_req_bits_eccMask[4]; // @[DCache.scala 50:82]
  assign eccMask_5 = io_req_bits_eccMask[5]; // @[DCache.scala 50:82]
  assign eccMask_6 = io_req_bits_eccMask[6]; // @[DCache.scala 50:82]
  assign eccMask_7 = io_req_bits_eccMask[7]; // @[DCache.scala 50:82]
  assign rdata_lo = {data_arrays_0_3_rdata_data_data,data_arrays_0_2_rdata_data_data,data_arrays_0_1_rdata_data_data,data_arrays_0_0_rdata_data_data}; // @[Cat.scala 30:58]
  assign rdata_hi = {data_arrays_0_7_rdata_data_data,data_arrays_0_6_rdata_data_data,data_arrays_0_5_rdata_data_data,data_arrays_0_4_rdata_data_data}; // @[Cat.scala 30:58]
  assign lo = {data_arrays_0_11_rdata_data_data,data_arrays_0_10_rdata_data_data,data_arrays_0_9_rdata_data_data,data_arrays_0_8_rdata_data_data}; // @[Cat.scala 30:58]
  assign hi = {data_arrays_0_15_rdata_data_data,data_arrays_0_14_rdata_data_data,data_arrays_0_13_rdata_data_data,data_arrays_0_12_rdata_data_data}; // @[Cat.scala 30:58]
  assign lo_1 = {data_arrays_0_19_rdata_data_data,data_arrays_0_18_rdata_data_data,data_arrays_0_17_rdata_data_data,data_arrays_0_16_rdata_data_data}; // @[Cat.scala 30:58]
  assign hi_1 = {data_arrays_0_23_rdata_data_data,data_arrays_0_22_rdata_data_data,data_arrays_0_21_rdata_data_data,data_arrays_0_20_rdata_data_data}; // @[Cat.scala 30:58]
  assign lo_2 = {data_arrays_0_27_rdata_data_data,data_arrays_0_26_rdata_data_data,data_arrays_0_25_rdata_data_data,data_arrays_0_24_rdata_data_data}; // @[Cat.scala 30:58]
  assign hi_2 = {data_arrays_0_31_rdata_data_data,data_arrays_0_30_rdata_data_data,data_arrays_0_29_rdata_data_data,data_arrays_0_28_rdata_data_data}; // @[Cat.scala 30:58]
  assign io_resp_0 = {rdata_hi,rdata_lo}; // @[DCache.scala 74:69]
  assign io_resp_1 = {hi,lo}; // @[DCache.scala 74:69]
  assign io_resp_2 = {hi_1,lo_1}; // @[DCache.scala 74:69]
  assign io_resp_3 = {hi_2,lo_2}; // @[DCache.scala 74:69]
  assign DCacheDataArray_covSum = 30'h0;
  assign io_covSum = DCacheDataArray_covSum;
  assign metaAssert = 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_0[initvar] = _RAND_0[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  data_arrays_0_0_rdata_data_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  data_arrays_0_0_rdata_data_addr_pipe_0 = _RAND_2[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_1[initvar] = _RAND_3[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  data_arrays_0_1_rdata_data_en_pipe_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  data_arrays_0_1_rdata_data_addr_pipe_0 = _RAND_5[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_2[initvar] = _RAND_6[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  data_arrays_0_2_rdata_data_en_pipe_0 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  data_arrays_0_2_rdata_data_addr_pipe_0 = _RAND_8[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_3[initvar] = _RAND_9[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  data_arrays_0_3_rdata_data_en_pipe_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  data_arrays_0_3_rdata_data_addr_pipe_0 = _RAND_11[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_4[initvar] = _RAND_12[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  data_arrays_0_4_rdata_data_en_pipe_0 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  data_arrays_0_4_rdata_data_addr_pipe_0 = _RAND_14[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_5[initvar] = _RAND_15[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  data_arrays_0_5_rdata_data_en_pipe_0 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  data_arrays_0_5_rdata_data_addr_pipe_0 = _RAND_17[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_6[initvar] = _RAND_18[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  data_arrays_0_6_rdata_data_en_pipe_0 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  data_arrays_0_6_rdata_data_addr_pipe_0 = _RAND_20[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_7[initvar] = _RAND_21[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  data_arrays_0_7_rdata_data_en_pipe_0 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  data_arrays_0_7_rdata_data_addr_pipe_0 = _RAND_23[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_8[initvar] = _RAND_24[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  data_arrays_0_8_rdata_data_en_pipe_0 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  data_arrays_0_8_rdata_data_addr_pipe_0 = _RAND_26[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_9[initvar] = _RAND_27[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  data_arrays_0_9_rdata_data_en_pipe_0 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  data_arrays_0_9_rdata_data_addr_pipe_0 = _RAND_29[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_10[initvar] = _RAND_30[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  data_arrays_0_10_rdata_data_en_pipe_0 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  data_arrays_0_10_rdata_data_addr_pipe_0 = _RAND_32[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_11[initvar] = _RAND_33[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  data_arrays_0_11_rdata_data_en_pipe_0 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  data_arrays_0_11_rdata_data_addr_pipe_0 = _RAND_35[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_12[initvar] = _RAND_36[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  data_arrays_0_12_rdata_data_en_pipe_0 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  data_arrays_0_12_rdata_data_addr_pipe_0 = _RAND_38[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_13[initvar] = _RAND_39[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  data_arrays_0_13_rdata_data_en_pipe_0 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  data_arrays_0_13_rdata_data_addr_pipe_0 = _RAND_41[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_14[initvar] = _RAND_42[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  data_arrays_0_14_rdata_data_en_pipe_0 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  data_arrays_0_14_rdata_data_addr_pipe_0 = _RAND_44[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_15[initvar] = _RAND_45[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  data_arrays_0_15_rdata_data_en_pipe_0 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  data_arrays_0_15_rdata_data_addr_pipe_0 = _RAND_47[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_16[initvar] = _RAND_48[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  data_arrays_0_16_rdata_data_en_pipe_0 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  data_arrays_0_16_rdata_data_addr_pipe_0 = _RAND_50[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_17[initvar] = _RAND_51[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  data_arrays_0_17_rdata_data_en_pipe_0 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  data_arrays_0_17_rdata_data_addr_pipe_0 = _RAND_53[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_18[initvar] = _RAND_54[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  data_arrays_0_18_rdata_data_en_pipe_0 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  data_arrays_0_18_rdata_data_addr_pipe_0 = _RAND_56[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_19[initvar] = _RAND_57[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  data_arrays_0_19_rdata_data_en_pipe_0 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  data_arrays_0_19_rdata_data_addr_pipe_0 = _RAND_59[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_20[initvar] = _RAND_60[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  data_arrays_0_20_rdata_data_en_pipe_0 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  data_arrays_0_20_rdata_data_addr_pipe_0 = _RAND_62[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_21[initvar] = _RAND_63[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  data_arrays_0_21_rdata_data_en_pipe_0 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  data_arrays_0_21_rdata_data_addr_pipe_0 = _RAND_65[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_22[initvar] = _RAND_66[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  data_arrays_0_22_rdata_data_en_pipe_0 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  data_arrays_0_22_rdata_data_addr_pipe_0 = _RAND_68[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_23[initvar] = _RAND_69[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  data_arrays_0_23_rdata_data_en_pipe_0 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  data_arrays_0_23_rdata_data_addr_pipe_0 = _RAND_71[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_24[initvar] = _RAND_72[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  data_arrays_0_24_rdata_data_en_pipe_0 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  data_arrays_0_24_rdata_data_addr_pipe_0 = _RAND_74[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_25[initvar] = _RAND_75[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  data_arrays_0_25_rdata_data_en_pipe_0 = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  data_arrays_0_25_rdata_data_addr_pipe_0 = _RAND_77[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_26[initvar] = _RAND_78[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  data_arrays_0_26_rdata_data_en_pipe_0 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  data_arrays_0_26_rdata_data_addr_pipe_0 = _RAND_80[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_27[initvar] = _RAND_81[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  data_arrays_0_27_rdata_data_en_pipe_0 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  data_arrays_0_27_rdata_data_addr_pipe_0 = _RAND_83[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_28[initvar] = _RAND_84[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  data_arrays_0_28_rdata_data_en_pipe_0 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  data_arrays_0_28_rdata_data_addr_pipe_0 = _RAND_86[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_29[initvar] = _RAND_87[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  data_arrays_0_29_rdata_data_en_pipe_0 = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  data_arrays_0_29_rdata_data_addr_pipe_0 = _RAND_89[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_30[initvar] = _RAND_90[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  data_arrays_0_30_rdata_data_en_pipe_0 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  data_arrays_0_30_rdata_data_addr_pipe_0 = _RAND_92[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_31[initvar] = _RAND_93[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  data_arrays_0_31_rdata_data_en_pipe_0 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  data_arrays_0_31_rdata_data_addr_pipe_0 = _RAND_95[8:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(data_arrays_0_0_rdata_MPORT_en & data_arrays_0_0_rdata_MPORT_mask) begin
      data_arrays_0_0[data_arrays_0_0_rdata_MPORT_addr] <= data_arrays_0_0_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      data_arrays_0_0_rdata_data_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_0_rdata_data_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_0_rdata_data_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_0_rdata_data_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_1_rdata_MPORT_en & data_arrays_0_1_rdata_MPORT_mask) begin
      data_arrays_0_1[data_arrays_0_1_rdata_MPORT_addr] <= data_arrays_0_1_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      data_arrays_0_1_rdata_data_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_1_rdata_data_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_1_rdata_data_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_1_rdata_data_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_2_rdata_MPORT_en & data_arrays_0_2_rdata_MPORT_mask) begin
      data_arrays_0_2[data_arrays_0_2_rdata_MPORT_addr] <= data_arrays_0_2_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      data_arrays_0_2_rdata_data_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_2_rdata_data_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_2_rdata_data_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_2_rdata_data_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_3_rdata_MPORT_en & data_arrays_0_3_rdata_MPORT_mask) begin
      data_arrays_0_3[data_arrays_0_3_rdata_MPORT_addr] <= data_arrays_0_3_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      data_arrays_0_3_rdata_data_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_3_rdata_data_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_3_rdata_data_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_3_rdata_data_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_4_rdata_MPORT_en & data_arrays_0_4_rdata_MPORT_mask) begin
      data_arrays_0_4[data_arrays_0_4_rdata_MPORT_addr] <= data_arrays_0_4_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      data_arrays_0_4_rdata_data_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_4_rdata_data_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_4_rdata_data_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_4_rdata_data_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_5_rdata_MPORT_en & data_arrays_0_5_rdata_MPORT_mask) begin
      data_arrays_0_5[data_arrays_0_5_rdata_MPORT_addr] <= data_arrays_0_5_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      data_arrays_0_5_rdata_data_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_5_rdata_data_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_5_rdata_data_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_5_rdata_data_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_6_rdata_MPORT_en & data_arrays_0_6_rdata_MPORT_mask) begin
      data_arrays_0_6[data_arrays_0_6_rdata_MPORT_addr] <= data_arrays_0_6_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      data_arrays_0_6_rdata_data_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_6_rdata_data_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_6_rdata_data_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_6_rdata_data_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_7_rdata_MPORT_en & data_arrays_0_7_rdata_MPORT_mask) begin
      data_arrays_0_7[data_arrays_0_7_rdata_MPORT_addr] <= data_arrays_0_7_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      data_arrays_0_7_rdata_data_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_7_rdata_data_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_7_rdata_data_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_7_rdata_data_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_8_rdata_MPORT_en & data_arrays_0_8_rdata_MPORT_mask) begin
      data_arrays_0_8[data_arrays_0_8_rdata_MPORT_addr] <= data_arrays_0_8_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      data_arrays_0_8_rdata_data_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_8_rdata_data_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_8_rdata_data_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_8_rdata_data_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_9_rdata_MPORT_en & data_arrays_0_9_rdata_MPORT_mask) begin
      data_arrays_0_9[data_arrays_0_9_rdata_MPORT_addr] <= data_arrays_0_9_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      data_arrays_0_9_rdata_data_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_9_rdata_data_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_9_rdata_data_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_9_rdata_data_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_10_rdata_MPORT_en & data_arrays_0_10_rdata_MPORT_mask) begin
      data_arrays_0_10[data_arrays_0_10_rdata_MPORT_addr] <= data_arrays_0_10_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      data_arrays_0_10_rdata_data_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_10_rdata_data_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_10_rdata_data_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_10_rdata_data_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_11_rdata_MPORT_en & data_arrays_0_11_rdata_MPORT_mask) begin
      data_arrays_0_11[data_arrays_0_11_rdata_MPORT_addr] <= data_arrays_0_11_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      data_arrays_0_11_rdata_data_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_11_rdata_data_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_11_rdata_data_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_11_rdata_data_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_12_rdata_MPORT_en & data_arrays_0_12_rdata_MPORT_mask) begin
      data_arrays_0_12[data_arrays_0_12_rdata_MPORT_addr] <= data_arrays_0_12_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      data_arrays_0_12_rdata_data_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_12_rdata_data_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_12_rdata_data_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_12_rdata_data_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_13_rdata_MPORT_en & data_arrays_0_13_rdata_MPORT_mask) begin
      data_arrays_0_13[data_arrays_0_13_rdata_MPORT_addr] <= data_arrays_0_13_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      data_arrays_0_13_rdata_data_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_13_rdata_data_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_13_rdata_data_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_13_rdata_data_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_14_rdata_MPORT_en & data_arrays_0_14_rdata_MPORT_mask) begin
      data_arrays_0_14[data_arrays_0_14_rdata_MPORT_addr] <= data_arrays_0_14_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      data_arrays_0_14_rdata_data_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_14_rdata_data_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_14_rdata_data_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_14_rdata_data_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_15_rdata_MPORT_en & data_arrays_0_15_rdata_MPORT_mask) begin
      data_arrays_0_15[data_arrays_0_15_rdata_MPORT_addr] <= data_arrays_0_15_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      data_arrays_0_15_rdata_data_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_15_rdata_data_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_15_rdata_data_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_15_rdata_data_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_16_rdata_MPORT_en & data_arrays_0_16_rdata_MPORT_mask) begin
      data_arrays_0_16[data_arrays_0_16_rdata_MPORT_addr] <= data_arrays_0_16_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      data_arrays_0_16_rdata_data_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_16_rdata_data_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_16_rdata_data_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_16_rdata_data_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_17_rdata_MPORT_en & data_arrays_0_17_rdata_MPORT_mask) begin
      data_arrays_0_17[data_arrays_0_17_rdata_MPORT_addr] <= data_arrays_0_17_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      data_arrays_0_17_rdata_data_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_17_rdata_data_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_17_rdata_data_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_17_rdata_data_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_18_rdata_MPORT_en & data_arrays_0_18_rdata_MPORT_mask) begin
      data_arrays_0_18[data_arrays_0_18_rdata_MPORT_addr] <= data_arrays_0_18_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      data_arrays_0_18_rdata_data_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_18_rdata_data_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_18_rdata_data_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_18_rdata_data_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_19_rdata_MPORT_en & data_arrays_0_19_rdata_MPORT_mask) begin
      data_arrays_0_19[data_arrays_0_19_rdata_MPORT_addr] <= data_arrays_0_19_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      data_arrays_0_19_rdata_data_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_19_rdata_data_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_19_rdata_data_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_19_rdata_data_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_20_rdata_MPORT_en & data_arrays_0_20_rdata_MPORT_mask) begin
      data_arrays_0_20[data_arrays_0_20_rdata_MPORT_addr] <= data_arrays_0_20_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      data_arrays_0_20_rdata_data_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_20_rdata_data_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_20_rdata_data_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_20_rdata_data_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_21_rdata_MPORT_en & data_arrays_0_21_rdata_MPORT_mask) begin
      data_arrays_0_21[data_arrays_0_21_rdata_MPORT_addr] <= data_arrays_0_21_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      data_arrays_0_21_rdata_data_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_21_rdata_data_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_21_rdata_data_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_21_rdata_data_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_22_rdata_MPORT_en & data_arrays_0_22_rdata_MPORT_mask) begin
      data_arrays_0_22[data_arrays_0_22_rdata_MPORT_addr] <= data_arrays_0_22_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      data_arrays_0_22_rdata_data_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_22_rdata_data_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_22_rdata_data_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_22_rdata_data_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_23_rdata_MPORT_en & data_arrays_0_23_rdata_MPORT_mask) begin
      data_arrays_0_23[data_arrays_0_23_rdata_MPORT_addr] <= data_arrays_0_23_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      data_arrays_0_23_rdata_data_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_23_rdata_data_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_23_rdata_data_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_23_rdata_data_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_24_rdata_MPORT_en & data_arrays_0_24_rdata_MPORT_mask) begin
      data_arrays_0_24[data_arrays_0_24_rdata_MPORT_addr] <= data_arrays_0_24_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      data_arrays_0_24_rdata_data_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_24_rdata_data_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_24_rdata_data_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_24_rdata_data_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_25_rdata_MPORT_en & data_arrays_0_25_rdata_MPORT_mask) begin
      data_arrays_0_25[data_arrays_0_25_rdata_MPORT_addr] <= data_arrays_0_25_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      data_arrays_0_25_rdata_data_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_25_rdata_data_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_25_rdata_data_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_25_rdata_data_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_26_rdata_MPORT_en & data_arrays_0_26_rdata_MPORT_mask) begin
      data_arrays_0_26[data_arrays_0_26_rdata_MPORT_addr] <= data_arrays_0_26_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      data_arrays_0_26_rdata_data_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_26_rdata_data_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_26_rdata_data_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_26_rdata_data_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_27_rdata_MPORT_en & data_arrays_0_27_rdata_MPORT_mask) begin
      data_arrays_0_27[data_arrays_0_27_rdata_MPORT_addr] <= data_arrays_0_27_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      data_arrays_0_27_rdata_data_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_27_rdata_data_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_27_rdata_data_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_27_rdata_data_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_28_rdata_MPORT_en & data_arrays_0_28_rdata_MPORT_mask) begin
      data_arrays_0_28[data_arrays_0_28_rdata_MPORT_addr] <= data_arrays_0_28_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      data_arrays_0_28_rdata_data_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_28_rdata_data_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_28_rdata_data_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_28_rdata_data_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_29_rdata_MPORT_en & data_arrays_0_29_rdata_MPORT_mask) begin
      data_arrays_0_29[data_arrays_0_29_rdata_MPORT_addr] <= data_arrays_0_29_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      data_arrays_0_29_rdata_data_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_29_rdata_data_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_29_rdata_data_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_29_rdata_data_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_30_rdata_MPORT_en & data_arrays_0_30_rdata_MPORT_mask) begin
      data_arrays_0_30[data_arrays_0_30_rdata_MPORT_addr] <= data_arrays_0_30_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      data_arrays_0_30_rdata_data_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_30_rdata_data_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_30_rdata_data_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_30_rdata_data_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
    if(data_arrays_0_31_rdata_MPORT_en & data_arrays_0_31_rdata_MPORT_mask) begin
      data_arrays_0_31[data_arrays_0_31_rdata_MPORT_addr] <= data_arrays_0_31_rdata_MPORT_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      data_arrays_0_31_rdata_data_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_31_rdata_data_en_pipe_0 <= io_req_valid & ~io_req_bits_write;
    end
    if (metaReset) begin
      data_arrays_0_31_rdata_data_addr_pipe_0 <= 9'h0;
    end else if (io_req_valid & ~io_req_bits_write) begin
      data_arrays_0_31_rdata_data_addr_pipe_0 <= io_req_bits_addr[11:3];
    end
  end
endmodule
module DCacheModuleImpl_Anon_2(
  input         io_in_0_valid,
  input  [11:0] io_in_0_bits_addr,
  input         io_in_0_bits_write,
  input  [63:0] io_in_0_bits_wdata,
  input  [7:0]  io_in_0_bits_eccMask,
  input  [3:0]  io_in_0_bits_way_en,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [11:0] io_in_1_bits_addr,
  input         io_in_1_bits_write,
  input  [63:0] io_in_1_bits_wdata,
  input  [3:0]  io_in_1_bits_way_en,
  output        io_in_2_ready,
  input         io_in_2_valid,
  input  [11:0] io_in_2_bits_addr,
  input  [63:0] io_in_2_bits_wdata,
  output        io_in_3_ready,
  input         io_in_3_valid,
  input  [11:0] io_in_3_bits_addr,
  input  [63:0] io_in_3_bits_wdata,
  input         io_in_3_bits_wordMask,
  output        io_out_valid,
  output [11:0] io_out_bits_addr,
  output        io_out_bits_write,
  output [63:0] io_out_bits_wdata,
  output [7:0]  io_out_bits_eccMask,
  output [3:0]  io_out_bits_way_en,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire [63:0] _GEN_4; // @[Arbiter.scala 126:27]
  wire [11:0] _GEN_6; // @[Arbiter.scala 126:27]
  wire [3:0] _GEN_8; // @[Arbiter.scala 126:27]
  wire [63:0] _GEN_11; // @[Arbiter.scala 126:27]
  wire  _GEN_12; // @[Arbiter.scala 126:27]
  wire [11:0] _GEN_13; // @[Arbiter.scala 126:27]
  wire  _grant_T; // @[Arbiter.scala 31:68]
  wire  _grant_T_1; // @[Arbiter.scala 31:68]
  wire  grant_3; // @[Arbiter.scala 31:78]
  wire [29:0] DCacheModuleImpl_Anon_2_covSum;
  assign _GEN_4 = io_in_2_valid ? io_in_2_bits_wdata : io_in_3_bits_wdata; // @[Arbiter.scala 126:27]
  assign _GEN_6 = io_in_2_valid ? io_in_2_bits_addr : io_in_3_bits_addr; // @[Arbiter.scala 126:27]
  assign _GEN_8 = io_in_1_valid ? io_in_1_bits_way_en : 4'hf; // @[Arbiter.scala 126:27]
  assign _GEN_11 = io_in_1_valid ? io_in_1_bits_wdata : _GEN_4; // @[Arbiter.scala 126:27]
  assign _GEN_12 = io_in_1_valid & io_in_1_bits_write; // @[Arbiter.scala 126:27]
  assign _GEN_13 = io_in_1_valid ? io_in_1_bits_addr : _GEN_6; // @[Arbiter.scala 126:27]
  assign _grant_T = io_in_0_valid | io_in_1_valid; // @[Arbiter.scala 31:68]
  assign _grant_T_1 = _grant_T | io_in_2_valid; // @[Arbiter.scala 31:68]
  assign grant_3 = ~_grant_T_1; // @[Arbiter.scala 31:78]
  assign io_in_1_ready = ~io_in_0_valid; // @[Arbiter.scala 134:14]
  assign io_in_2_ready = ~_grant_T; // @[Arbiter.scala 134:14]
  assign io_in_3_ready = ~_grant_T_1; // @[Arbiter.scala 134:14]
  assign io_out_valid = ~grant_3 | io_in_3_valid; // @[Arbiter.scala 135:16]
  assign io_out_bits_addr = io_in_0_valid ? io_in_0_bits_addr : _GEN_13; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign io_out_bits_write = io_in_0_valid ? io_in_0_bits_write : _GEN_12; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign io_out_bits_wdata = io_in_0_valid ? io_in_0_bits_wdata : _GEN_11; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign io_out_bits_eccMask = io_in_0_valid ? io_in_0_bits_eccMask : 8'hff; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign io_out_bits_way_en = io_in_0_valid ? io_in_0_bits_way_en : _GEN_8; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign DCacheModuleImpl_Anon_2_covSum = 30'h0;
  assign io_covSum = DCacheModuleImpl_Anon_2_covSum;
  assign metaAssert = 1'h0;
endmodule
module AMOALU(
  input  [7:0]  io_mask,
  input  [4:0]  io_cmd,
  input  [63:0] io_lhs,
  input  [63:0] io_rhs,
  output [63:0] io_out,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  _max_T; // @[AMOALU.scala 64:20]
  wire  _max_T_1; // @[AMOALU.scala 64:43]
  wire  max; // @[AMOALU.scala 64:33]
  wire  _min_T; // @[AMOALU.scala 65:20]
  wire  _min_T_1; // @[AMOALU.scala 65:43]
  wire  min; // @[AMOALU.scala 65:33]
  wire  add; // @[AMOALU.scala 66:20]
  wire  _logic_and_T; // @[AMOALU.scala 67:26]
  wire  _logic_and_T_1; // @[AMOALU.scala 67:48]
  wire  logic_and; // @[AMOALU.scala 67:38]
  wire  _logic_xor_T; // @[AMOALU.scala 68:26]
  wire  logic_xor; // @[AMOALU.scala 68:39]
  wire [31:0] _adder_out_mask_T_2; // @[AMOALU.scala 72:79]
  wire [63:0] _adder_out_mask_T_3; // @[AMOALU.scala 72:98]
  wire [63:0] adder_out_mask; // @[AMOALU.scala 72:16]
  wire [63:0] _adder_out_T; // @[AMOALU.scala 73:13]
  wire [63:0] _adder_out_T_1; // @[AMOALU.scala 73:31]
  wire [63:0] adder_out; // @[AMOALU.scala 73:21]
  wire [4:0] _less_signed_T; // @[AMOALU.scala 86:17]
  wire  less_signed; // @[AMOALU.scala 86:25]
  wire  _less_T_3; // @[AMOALU.scala 88:18]
  wire  _less_T_6; // @[AMOALU.scala 80:24]
  wire  _less_T_9; // @[AMOALU.scala 80:53]
  wire  _less_T_12; // @[AMOALU.scala 79:35]
  wire  _less_T_13; // @[AMOALU.scala 80:69]
  wire  _less_T_14; // @[AMOALU.scala 80:38]
  wire  _less_T_17; // @[AMOALU.scala 88:58]
  wire  _less_T_18; // @[AMOALU.scala 88:10]
  wire  _less_T_22; // @[AMOALU.scala 88:18]
  wire  _less_T_28; // @[AMOALU.scala 88:58]
  wire  _less_T_29; // @[AMOALU.scala 88:10]
  wire  less; // @[Mux.scala 47:69]
  wire  _minmax_T; // @[AMOALU.scala 94:23]
  wire [63:0] minmax; // @[AMOALU.scala 94:19]
  wire [63:0] _logic_T; // @[AMOALU.scala 96:27]
  wire [63:0] _logic_T_1; // @[AMOALU.scala 96:8]
  wire [63:0] _logic_T_2; // @[AMOALU.scala 97:27]
  wire [63:0] _logic_T_3; // @[AMOALU.scala 97:8]
  wire [63:0] logic_; // @[AMOALU.scala 96:42]
  wire  _out_T; // @[AMOALU.scala 100:19]
  wire [63:0] _out_T_1; // @[AMOALU.scala 100:8]
  wire [63:0] out; // @[AMOALU.scala 99:8]
  wire [7:0] wmask_lo_lo_lo; // @[Bitwise.scala 72:12]
  wire [7:0] wmask_lo_lo_hi; // @[Bitwise.scala 72:12]
  wire [7:0] wmask_lo_hi_lo; // @[Bitwise.scala 72:12]
  wire [7:0] wmask_lo_hi_hi; // @[Bitwise.scala 72:12]
  wire [7:0] wmask_hi_lo_lo; // @[Bitwise.scala 72:12]
  wire [7:0] wmask_hi_lo_hi; // @[Bitwise.scala 72:12]
  wire [7:0] wmask_hi_hi_lo; // @[Bitwise.scala 72:12]
  wire [7:0] wmask_hi_hi_hi; // @[Bitwise.scala 72:12]
  wire [63:0] wmask; // @[Cat.scala 30:58]
  wire [63:0] _io_out_T; // @[AMOALU.scala 104:19]
  wire [63:0] _io_out_T_2; // @[AMOALU.scala 104:34]
  wire [29:0] AMOALU_covSum;
  assign _max_T = io_cmd == 5'hd; // @[AMOALU.scala 64:20]
  assign _max_T_1 = io_cmd == 5'hf; // @[AMOALU.scala 64:43]
  assign max = _max_T | _max_T_1; // @[AMOALU.scala 64:33]
  assign _min_T = io_cmd == 5'hc; // @[AMOALU.scala 65:20]
  assign _min_T_1 = io_cmd == 5'he; // @[AMOALU.scala 65:43]
  assign min = _min_T | _min_T_1; // @[AMOALU.scala 65:33]
  assign add = io_cmd == 5'h8; // @[AMOALU.scala 66:20]
  assign _logic_and_T = io_cmd == 5'ha; // @[AMOALU.scala 67:26]
  assign _logic_and_T_1 = io_cmd == 5'hb; // @[AMOALU.scala 67:48]
  assign logic_and = _logic_and_T | _logic_and_T_1; // @[AMOALU.scala 67:38]
  assign _logic_xor_T = io_cmd == 5'h9; // @[AMOALU.scala 68:26]
  assign logic_xor = _logic_xor_T | _logic_and_T; // @[AMOALU.scala 68:39]
  assign _adder_out_mask_T_2 = {~io_mask[3], 31'h0}; // @[AMOALU.scala 72:79]
  assign _adder_out_mask_T_3 = {{32'd0}, _adder_out_mask_T_2}; // @[AMOALU.scala 72:98]
  assign adder_out_mask = ~_adder_out_mask_T_3; // @[AMOALU.scala 72:16]
  assign _adder_out_T = io_lhs & adder_out_mask; // @[AMOALU.scala 73:13]
  assign _adder_out_T_1 = io_rhs & adder_out_mask; // @[AMOALU.scala 73:31]
  assign adder_out = _adder_out_T + _adder_out_T_1; // @[AMOALU.scala 73:21]
  assign _less_signed_T = io_cmd & 5'h2; // @[AMOALU.scala 86:17]
  assign less_signed = _less_signed_T == 5'h0; // @[AMOALU.scala 86:25]
  assign _less_T_3 = io_lhs[63] == io_rhs[63]; // @[AMOALU.scala 88:18]
  assign _less_T_6 = io_lhs[63:32] < io_rhs[63:32]; // @[AMOALU.scala 80:24]
  assign _less_T_9 = io_lhs[63:32] == io_rhs[63:32]; // @[AMOALU.scala 80:53]
  assign _less_T_12 = io_lhs[31:0] < io_rhs[31:0]; // @[AMOALU.scala 79:35]
  assign _less_T_13 = _less_T_9 & _less_T_12; // @[AMOALU.scala 80:69]
  assign _less_T_14 = _less_T_6 | _less_T_13; // @[AMOALU.scala 80:38]
  assign _less_T_17 = less_signed ? io_lhs[63] : io_rhs[63]; // @[AMOALU.scala 88:58]
  assign _less_T_18 = _less_T_3 ? _less_T_14 : _less_T_17; // @[AMOALU.scala 88:10]
  assign _less_T_22 = io_lhs[31] == io_rhs[31]; // @[AMOALU.scala 88:18]
  assign _less_T_28 = less_signed ? io_lhs[31] : io_rhs[31]; // @[AMOALU.scala 88:58]
  assign _less_T_29 = _less_T_22 ? _less_T_12 : _less_T_28; // @[AMOALU.scala 88:10]
  assign less = io_mask[4] ? _less_T_18 : _less_T_29; // @[Mux.scala 47:69]
  assign _minmax_T = less ? min : max; // @[AMOALU.scala 94:23]
  assign minmax = _minmax_T ? io_lhs : io_rhs; // @[AMOALU.scala 94:19]
  assign _logic_T = io_lhs & io_rhs; // @[AMOALU.scala 96:27]
  assign _logic_T_1 = logic_and ? _logic_T : 64'h0; // @[AMOALU.scala 96:8]
  assign _logic_T_2 = io_lhs ^ io_rhs; // @[AMOALU.scala 97:27]
  assign _logic_T_3 = logic_xor ? _logic_T_2 : 64'h0; // @[AMOALU.scala 97:8]
  assign logic_ = _logic_T_1 | _logic_T_3; // @[AMOALU.scala 96:42]
  assign _out_T = logic_and | logic_xor; // @[AMOALU.scala 100:19]
  assign _out_T_1 = _out_T ? logic_ : minmax; // @[AMOALU.scala 100:8]
  assign out = add ? adder_out : _out_T_1; // @[AMOALU.scala 99:8]
  assign wmask_lo_lo_lo = io_mask[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign wmask_lo_lo_hi = io_mask[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign wmask_lo_hi_lo = io_mask[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign wmask_lo_hi_hi = io_mask[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign wmask_hi_lo_lo = io_mask[4] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign wmask_hi_lo_hi = io_mask[5] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign wmask_hi_hi_lo = io_mask[6] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign wmask_hi_hi_hi = io_mask[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign wmask = {wmask_hi_hi_hi,wmask_hi_hi_lo,wmask_hi_lo_hi,wmask_hi_lo_lo,wmask_lo_hi_hi,wmask_lo_hi_lo,wmask_lo_lo_hi,wmask_lo_lo_lo}; // @[Cat.scala 30:58]
  assign _io_out_T = wmask & out; // @[AMOALU.scala 104:19]
  assign _io_out_T_2 = ~wmask & io_lhs; // @[AMOALU.scala 104:34]
  assign io_out = _io_out_T | _io_out_T_2; // @[AMOALU.scala 104:10]
  assign AMOALU_covSum = 30'h0;
  assign io_covSum = AMOALU_covSum;
  assign metaAssert = 1'h0;
endmodule
module ICache(
  input         clock,
  input         reset,
  input         auto_master_out_a_ready,
  output        auto_master_out_a_valid,
  output [31:0] auto_master_out_a_bits_address,
  input         auto_master_out_d_valid,
  input  [2:0]  auto_master_out_d_bits_opcode,
  input  [3:0]  auto_master_out_d_bits_size,
  input  [63:0] auto_master_out_d_bits_data,
  input         auto_master_out_d_bits_corrupt,
  output        io_req_ready,
  input         io_req_valid,
  input  [38:0] io_req_bits_addr,
  input  [31:0] io_s1_paddr,
  input         io_s1_kill,
  input         io_s2_kill,
  output        io_resp_valid,
  output [31:0] io_resp_bits_data,
  output        io_resp_bits_replay,
  output        io_resp_bits_ae,
  input         io_invalidate,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset,
  input         repl_way_v0_prng_halt
);
  wire  repl_way_v0_prng_clock; // @[PRNG.scala 82:22]
  wire  repl_way_v0_prng_reset; // @[PRNG.scala 82:22]
  wire  repl_way_v0_prng_io_increment; // @[PRNG.scala 82:22]
  wire  repl_way_v0_prng_io_out_0; // @[PRNG.scala 82:22]
  wire  repl_way_v0_prng_io_out_1; // @[PRNG.scala 82:22]
  wire  repl_way_v0_prng_io_out_2; // @[PRNG.scala 82:22]
  wire  repl_way_v0_prng_io_out_3; // @[PRNG.scala 82:22]
  wire  repl_way_v0_prng_io_out_4; // @[PRNG.scala 82:22]
  wire  repl_way_v0_prng_io_out_5; // @[PRNG.scala 82:22]
  wire  repl_way_v0_prng_io_out_6; // @[PRNG.scala 82:22]
  wire  repl_way_v0_prng_io_out_7; // @[PRNG.scala 82:22]
  wire  repl_way_v0_prng_io_out_8; // @[PRNG.scala 82:22]
  wire  repl_way_v0_prng_io_out_9; // @[PRNG.scala 82:22]
  wire  repl_way_v0_prng_io_out_10; // @[PRNG.scala 82:22]
  wire  repl_way_v0_prng_io_out_11; // @[PRNG.scala 82:22]
  wire  repl_way_v0_prng_io_out_12; // @[PRNG.scala 82:22]
  wire  repl_way_v0_prng_io_out_13; // @[PRNG.scala 82:22]
  wire  repl_way_v0_prng_io_out_14; // @[PRNG.scala 82:22]
  wire  repl_way_v0_prng_io_out_15; // @[PRNG.scala 82:22]
  wire [29:0] repl_way_v0_prng_io_covSum; // @[PRNG.scala 82:22]
  wire  repl_way_v0_prng_metaAssert; // @[PRNG.scala 82:22]
  wire  repl_way_v0_prng_metaReset; // @[PRNG.scala 82:22]
  reg [20:0] tag_array_0 [0:63]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_0;
  wire [20:0] tag_array_0_tag_rdata_data; // @[DescribedSRAM.scala 19:26]
  wire [5:0] tag_array_0_tag_rdata_addr; // @[DescribedSRAM.scala 19:26]
  wire [20:0] tag_array_0_MPORT_data; // @[DescribedSRAM.scala 19:26]
  wire [5:0] tag_array_0_MPORT_addr; // @[DescribedSRAM.scala 19:26]
  wire  tag_array_0_MPORT_mask; // @[DescribedSRAM.scala 19:26]
  wire  tag_array_0_MPORT_en; // @[DescribedSRAM.scala 19:26]
  reg  tag_array_0_tag_rdata_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [5:0] tag_array_0_tag_rdata_addr_pipe_0;
  reg [31:0] _RAND_2;
  reg [20:0] tag_array_1 [0:63]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_3;
  wire [20:0] tag_array_1_tag_rdata_data; // @[DescribedSRAM.scala 19:26]
  wire [5:0] tag_array_1_tag_rdata_addr; // @[DescribedSRAM.scala 19:26]
  wire [20:0] tag_array_1_MPORT_data; // @[DescribedSRAM.scala 19:26]
  wire [5:0] tag_array_1_MPORT_addr; // @[DescribedSRAM.scala 19:26]
  wire  tag_array_1_MPORT_mask; // @[DescribedSRAM.scala 19:26]
  wire  tag_array_1_MPORT_en; // @[DescribedSRAM.scala 19:26]
  reg  tag_array_1_tag_rdata_en_pipe_0;
  reg [31:0] _RAND_4;
  reg [5:0] tag_array_1_tag_rdata_addr_pipe_0;
  reg [31:0] _RAND_5;
  reg [20:0] tag_array_2 [0:63]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_6;
  wire [20:0] tag_array_2_tag_rdata_data; // @[DescribedSRAM.scala 19:26]
  wire [5:0] tag_array_2_tag_rdata_addr; // @[DescribedSRAM.scala 19:26]
  wire [20:0] tag_array_2_MPORT_data; // @[DescribedSRAM.scala 19:26]
  wire [5:0] tag_array_2_MPORT_addr; // @[DescribedSRAM.scala 19:26]
  wire  tag_array_2_MPORT_mask; // @[DescribedSRAM.scala 19:26]
  wire  tag_array_2_MPORT_en; // @[DescribedSRAM.scala 19:26]
  reg  tag_array_2_tag_rdata_en_pipe_0;
  reg [31:0] _RAND_7;
  reg [5:0] tag_array_2_tag_rdata_addr_pipe_0;
  reg [31:0] _RAND_8;
  reg [20:0] tag_array_3 [0:63]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_9;
  wire [20:0] tag_array_3_tag_rdata_data; // @[DescribedSRAM.scala 19:26]
  wire [5:0] tag_array_3_tag_rdata_addr; // @[DescribedSRAM.scala 19:26]
  wire [20:0] tag_array_3_MPORT_data; // @[DescribedSRAM.scala 19:26]
  wire [5:0] tag_array_3_MPORT_addr; // @[DescribedSRAM.scala 19:26]
  wire  tag_array_3_MPORT_mask; // @[DescribedSRAM.scala 19:26]
  wire  tag_array_3_MPORT_en; // @[DescribedSRAM.scala 19:26]
  reg  tag_array_3_tag_rdata_en_pipe_0;
  reg [31:0] _RAND_10;
  reg [5:0] tag_array_3_tag_rdata_addr_pipe_0;
  reg [31:0] _RAND_11;
  reg [31:0] data_arrays_0_0 [0:511]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_12;
  wire [31:0] data_arrays_0_0_dout_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_0_dout_addr; // @[DescribedSRAM.scala 19:26]
  wire [31:0] data_arrays_0_0_MPORT_1_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_0_MPORT_1_addr; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_0_MPORT_1_mask; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_0_MPORT_1_en; // @[DescribedSRAM.scala 19:26]
  reg  data_arrays_0_0_dout_en_pipe_0;
  reg [31:0] _RAND_13;
  reg [8:0] data_arrays_0_0_dout_addr_pipe_0;
  reg [31:0] _RAND_14;
  reg [31:0] data_arrays_0_1 [0:511]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_15;
  wire [31:0] data_arrays_0_1_dout_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_1_dout_addr; // @[DescribedSRAM.scala 19:26]
  wire [31:0] data_arrays_0_1_MPORT_1_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_1_MPORT_1_addr; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_1_MPORT_1_mask; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_1_MPORT_1_en; // @[DescribedSRAM.scala 19:26]
  reg  data_arrays_0_1_dout_en_pipe_0;
  reg [31:0] _RAND_16;
  reg [8:0] data_arrays_0_1_dout_addr_pipe_0;
  reg [31:0] _RAND_17;
  reg [31:0] data_arrays_0_2 [0:511]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_18;
  wire [31:0] data_arrays_0_2_dout_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_2_dout_addr; // @[DescribedSRAM.scala 19:26]
  wire [31:0] data_arrays_0_2_MPORT_1_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_2_MPORT_1_addr; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_2_MPORT_1_mask; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_2_MPORT_1_en; // @[DescribedSRAM.scala 19:26]
  reg  data_arrays_0_2_dout_en_pipe_0;
  reg [31:0] _RAND_19;
  reg [8:0] data_arrays_0_2_dout_addr_pipe_0;
  reg [31:0] _RAND_20;
  reg [31:0] data_arrays_0_3 [0:511]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_21;
  wire [31:0] data_arrays_0_3_dout_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_3_dout_addr; // @[DescribedSRAM.scala 19:26]
  wire [31:0] data_arrays_0_3_MPORT_1_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_0_3_MPORT_1_addr; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_3_MPORT_1_mask; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_0_3_MPORT_1_en; // @[DescribedSRAM.scala 19:26]
  reg  data_arrays_0_3_dout_en_pipe_0;
  reg [31:0] _RAND_22;
  reg [8:0] data_arrays_0_3_dout_addr_pipe_0;
  reg [31:0] _RAND_23;
  reg [31:0] data_arrays_1_0 [0:511]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_24;
  wire [31:0] data_arrays_1_0_dout_1_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_1_0_dout_1_addr; // @[DescribedSRAM.scala 19:26]
  wire [31:0] data_arrays_1_0_MPORT_2_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_1_0_MPORT_2_addr; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_1_0_MPORT_2_mask; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_1_0_MPORT_2_en; // @[DescribedSRAM.scala 19:26]
  reg  data_arrays_1_0_dout_1_en_pipe_0;
  reg [31:0] _RAND_25;
  reg [8:0] data_arrays_1_0_dout_1_addr_pipe_0;
  reg [31:0] _RAND_26;
  reg [31:0] data_arrays_1_1 [0:511]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_27;
  wire [31:0] data_arrays_1_1_dout_1_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_1_1_dout_1_addr; // @[DescribedSRAM.scala 19:26]
  wire [31:0] data_arrays_1_1_MPORT_2_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_1_1_MPORT_2_addr; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_1_1_MPORT_2_mask; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_1_1_MPORT_2_en; // @[DescribedSRAM.scala 19:26]
  reg  data_arrays_1_1_dout_1_en_pipe_0;
  reg [31:0] _RAND_28;
  reg [8:0] data_arrays_1_1_dout_1_addr_pipe_0;
  reg [31:0] _RAND_29;
  reg [31:0] data_arrays_1_2 [0:511]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_30;
  wire [31:0] data_arrays_1_2_dout_1_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_1_2_dout_1_addr; // @[DescribedSRAM.scala 19:26]
  wire [31:0] data_arrays_1_2_MPORT_2_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_1_2_MPORT_2_addr; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_1_2_MPORT_2_mask; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_1_2_MPORT_2_en; // @[DescribedSRAM.scala 19:26]
  reg  data_arrays_1_2_dout_1_en_pipe_0;
  reg [31:0] _RAND_31;
  reg [8:0] data_arrays_1_2_dout_1_addr_pipe_0;
  reg [31:0] _RAND_32;
  reg [31:0] data_arrays_1_3 [0:511]; // @[DescribedSRAM.scala 19:26]
  reg [31:0] _RAND_33;
  wire [31:0] data_arrays_1_3_dout_1_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_1_3_dout_1_addr; // @[DescribedSRAM.scala 19:26]
  wire [31:0] data_arrays_1_3_MPORT_2_data; // @[DescribedSRAM.scala 19:26]
  wire [8:0] data_arrays_1_3_MPORT_2_addr; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_1_3_MPORT_2_mask; // @[DescribedSRAM.scala 19:26]
  wire  data_arrays_1_3_MPORT_2_en; // @[DescribedSRAM.scala 19:26]
  reg  data_arrays_1_3_dout_1_en_pipe_0;
  reg [31:0] _RAND_34;
  reg [8:0] data_arrays_1_3_dout_1_addr_pipe_0;
  reg [31:0] _RAND_35;
  wire  s0_valid; // @[Decoupled.scala 40:37]
  reg  s1_valid; // @[ICache.scala 169:21]
  reg [31:0] _RAND_36;
  reg [255:0] vb_array; // @[ICache.scala 231:21]
  reg [255:0] _RAND_37;
  wire [5:0] s1_vb_lo; // @[ICache.scala 486:21]
  wire [6:0] _s1_vb_T; // @[Cat.scala 30:58]
  wire [255:0] _s1_vb_T_1; // @[ICache.scala 259:25]
  wire  s1_vb; // @[ICache.scala 259:25]
  wire [19:0] tag; // @[package.scala 154:13]
  wire [19:0] s1_tag; // @[ICache.scala 254:30]
  wire  _tagMatch_T; // @[ICache.scala 262:33]
  wire  tagMatch; // @[ICache.scala 262:26]
  wire [6:0] _s1_vb_T_4; // @[Cat.scala 30:58]
  wire [255:0] _s1_vb_T_5; // @[ICache.scala 259:25]
  wire  s1_vb_1; // @[ICache.scala 259:25]
  wire [19:0] tag_1; // @[package.scala 154:13]
  wire  _tagMatch_T_1; // @[ICache.scala 262:33]
  wire  tagMatch_1; // @[ICache.scala 262:26]
  wire  _s1_hit_T; // @[ICache.scala 172:35]
  wire [7:0] _s1_vb_T_8; // @[Cat.scala 30:58]
  wire [255:0] _s1_vb_T_9; // @[ICache.scala 259:25]
  wire  s1_vb_2; // @[ICache.scala 259:25]
  wire [19:0] tag_2; // @[package.scala 154:13]
  wire  _tagMatch_T_2; // @[ICache.scala 262:33]
  wire  tagMatch_2; // @[ICache.scala 262:26]
  wire  _s1_hit_T_1; // @[ICache.scala 172:35]
  wire [7:0] _s1_vb_T_12; // @[Cat.scala 30:58]
  wire [255:0] _s1_vb_T_13; // @[ICache.scala 259:25]
  wire  s1_vb_3; // @[ICache.scala 259:25]
  wire [19:0] tag_3; // @[package.scala 154:13]
  wire  _tagMatch_T_3; // @[ICache.scala 262:33]
  wire  tagMatch_3; // @[ICache.scala 262:26]
  wire  _s2_valid_T_1; // @[ICache.scala 174:35]
  reg  s2_valid; // @[ICache.scala 174:25]
  reg [31:0] _RAND_38;
  reg  s2_hit; // @[ICache.scala 175:23]
  reg [31:0] _RAND_39;
  reg  invalidated; // @[ICache.scala 177:24]
  reg [31:0] _RAND_40;
  reg  refill_valid; // @[ICache.scala 178:29]
  reg [31:0] _RAND_41;
  wire  _s2_miss_T_1; // @[ICache.scala 182:26]
  wire  s2_miss; // @[ICache.scala 182:37]
  reg  s2_request_refill_REG; // @[ICache.scala 184:45]
  reg [31:0] _RAND_42;
  wire  s2_request_refill; // @[ICache.scala 184:35]
  wire  refill_fire; // @[Decoupled.scala 40:37]
  wire  _s1_can_request_refill_T; // @[ICache.scala 183:41]
  wire  s1_can_request_refill; // @[ICache.scala 183:31]
  wire  _refill_paddr_T; // @[ICache.scala 185:54]
  reg [31:0] refill_paddr; // @[Reg.scala 15:16]
  reg [31:0] _RAND_43;
  wire [19:0] refill_tag; // @[ICache.scala 187:33]
  wire [5:0] refill_idx; // @[ICache.scala 486:21]
  wire  refill_one_beat_opdata; // @[Edges.scala 105:36]
  wire  refill_one_beat; // @[ICache.scala 189:41]
  wire [26:0] _beats1_decode_T_1; // @[package.scala 234:77]
  wire [8:0] beats1_decode; // @[Edges.scala 219:59]
  wire [8:0] beats1; // @[Edges.scala 220:14]
  reg [8:0] counter; // @[Edges.scala 228:27]
  reg [31:0] _RAND_44;
  wire [8:0] counter1; // @[Edges.scala 229:28]
  wire  first; // @[Edges.scala 230:25]
  wire  _last_T; // @[Edges.scala 231:25]
  wire  _last_T_1; // @[Edges.scala 231:47]
  wire  last; // @[Edges.scala 231:37]
  wire  d_done; // @[Edges.scala 232:22]
  wire [8:0] refill_cnt; // @[Edges.scala 233:25]
  wire  refill_done; // @[ICache.scala 195:37]
  wire [7:0] repl_way_v0_lo; // @[PRNG.scala 86:17]
  wire [15:0] _repl_way_v0_T; // @[PRNG.scala 86:17]
  wire [1:0] repl_way_v0; // @[ICache.scala 201:35]
  wire [7:0] _repl_way_T; // @[Cat.scala 30:58]
  reg  accruedRefillError; // @[ICache.scala 219:31]
  reg [31:0] _RAND_45;
  wire  _refillError_T; // @[ICache.scala 220:58]
  wire  _refillError_T_1; // @[ICache.scala 220:62]
  wire  refillError; // @[ICache.scala 220:43]
  wire  _vb_array_T_2; // @[ICache.scala 235:72]
  wire [255:0] _vb_array_T_3; // @[ICache.scala 235:32]
  wire [255:0] _vb_array_T_4; // @[ICache.scala 235:32]
  wire [255:0] _vb_array_T_6; // @[ICache.scala 235:32]
  wire  s2_tag_disparity; // @[ICache.scala 312:72]
  wire  _T_40; // @[ICache.scala 334:22]
  wire  invalidate; // @[ICache.scala 334:39]
  wire  _GEN_30; // @[ICache.scala 238:21]
  wire  tl_error; // @[package.scala 154:13]
  wire  s1_tl_error_0; // @[ICache.scala 264:32]
  wire  tl_error_1; // @[package.scala 154:13]
  wire  s1_tl_error_1; // @[ICache.scala 264:32]
  wire  tl_error_2; // @[package.scala 154:13]
  wire  s1_tl_error_2; // @[ICache.scala 264:32]
  wire  tl_error_3; // @[package.scala 154:13]
  wire  s1_tl_error_3; // @[ICache.scala 264:32]
  wire [1:0] _T_15; // @[Bitwise.scala 47:55]
  wire [1:0] _T_17; // @[Bitwise.scala 47:55]
  wire [2:0] _T_19; // @[Bitwise.scala 47:55]
  wire  _T_21; // @[ICache.scala 267:115]
  wire  _T_22; // @[ICache.scala 267:39]
  wire  _T_24; // @[ICache.scala 267:9]
  wire  s0_ren; // @[ICache.scala 284:28]
  wire  wen; // @[ICache.scala 285:32]
  wire [8:0] _mem_idx_T; // @[ICache.scala 286:52]
  wire [8:0] _mem_idx_T_1; // @[ICache.scala 286:79]
  wire [31:0] _GEN_54; // @[ICache.scala 296:71]
  wire [31:0] _GEN_55; // @[ICache.scala 296:71]
  wire [31:0] _GEN_56; // @[ICache.scala 296:71]
  wire [31:0] _GEN_57; // @[ICache.scala 296:71]
  wire  s0_ren_1; // @[ICache.scala 284:28]
  reg  s2_tag_hit_0; // @[Reg.scala 15:16]
  reg [31:0] _RAND_46;
  reg  s2_tag_hit_1; // @[Reg.scala 15:16]
  reg [31:0] _RAND_47;
  reg  s2_tag_hit_2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_48;
  reg  s2_tag_hit_3; // @[Reg.scala 15:16]
  reg [31:0] _RAND_49;
  reg [31:0] s2_dout_0; // @[Reg.scala 15:16]
  reg [31:0] _RAND_50;
  reg [31:0] s2_dout_1; // @[Reg.scala 15:16]
  reg [31:0] _RAND_51;
  reg [31:0] s2_dout_2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_52;
  reg [31:0] s2_dout_3; // @[Reg.scala 15:16]
  reg [31:0] _RAND_53;
  wire [31:0] _s2_way_mux_T; // @[Mux.scala 27:72]
  wire [31:0] _s2_way_mux_T_1; // @[Mux.scala 27:72]
  wire [31:0] _s2_way_mux_T_2; // @[Mux.scala 27:72]
  wire [31:0] _s2_way_mux_T_3; // @[Mux.scala 27:72]
  wire [31:0] _s2_way_mux_T_4; // @[Mux.scala 27:72]
  wire [31:0] _s2_way_mux_T_5; // @[Mux.scala 27:72]
  wire [3:0] _s2_tl_error_T; // @[ICache.scala 313:43]
  wire  _s2_tl_error_T_1; // @[ICache.scala 313:50]
  reg  s2_tl_error; // @[Reg.scala 15:16]
  reg [31:0] _RAND_54;
  wire  _GEN_101; // @[ICache.scala 477:22]
  reg [5:0] ICache_state; // @[Register tracking ICache state]
  reg [31:0] _RAND_55;
  reg  ICache_cov [0:63]; // @[Coverage map for ICache]
  reg [31:0] _RAND_56;
  wire  ICache_cov_read_data; // @[Coverage map for ICache]
  wire [5:0] ICache_cov_read_addr; // @[Coverage map for ICache]
  wire  ICache_cov_write_data; // @[Coverage map for ICache]
  wire [5:0] ICache_cov_write_addr; // @[Coverage map for ICache]
  wire  ICache_cov_write_mask; // @[Coverage map for ICache]
  wire  ICache_cov_write_en; // @[Coverage map for ICache]
  reg [29:0] ICache_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_57;
  wire  s2_valid_shl;
  wire [5:0] s2_valid_pad;
  wire [1:0] s1_valid_shl;
  wire [5:0] s1_valid_pad;
  wire [2:0] refill_valid_shl;
  wire [5:0] refill_valid_pad;
  wire [3:0] invalidated_shl;
  wire [5:0] invalidated_pad;
  wire [4:0] s2_hit_shl;
  wire [5:0] s2_hit_pad;
  wire [5:0] s2_tag_hit_0_shl;
  wire [5:0] s2_tag_hit_0_pad;
  wire [5:0] s2_tag_hit_1_shl;
  wire [5:0] s2_tag_hit_1_pad;
  wire [5:0] s2_tag_hit_2_shl;
  wire [5:0] s2_tag_hit_2_pad;
  wire [5:0] s2_tag_hit_3_shl;
  wire [5:0] s2_tag_hit_3_pad;
  wire [5:0] ICache_xor3;
  wire [5:0] ICache_xor4;
  wire [5:0] ICache_xor1;
  wire [5:0] ICache_xor5;
  wire [5:0] ICache_xor14;
  wire [5:0] ICache_xor6;
  wire [5:0] ICache_xor2;
  wire [5:0] ICache_xor0;
  wire [29:0] repl_way_v0_prng_sum;
  wire  stopEn0;
  wire  repl_way_v0_prng_metaAssert_wire;
  wire  ICache_or0;
  reg  ICache_metaAssert;
  reg [31:0] _RAND_58;
  MaxPeriodFibonacciLFSR repl_way_v0_prng ( // @[PRNG.scala 82:22]
    .clock(repl_way_v0_prng_clock),
    .reset(repl_way_v0_prng_reset),
    .io_increment(repl_way_v0_prng_io_increment),
    .io_out_0(repl_way_v0_prng_io_out_0),
    .io_out_1(repl_way_v0_prng_io_out_1),
    .io_out_2(repl_way_v0_prng_io_out_2),
    .io_out_3(repl_way_v0_prng_io_out_3),
    .io_out_4(repl_way_v0_prng_io_out_4),
    .io_out_5(repl_way_v0_prng_io_out_5),
    .io_out_6(repl_way_v0_prng_io_out_6),
    .io_out_7(repl_way_v0_prng_io_out_7),
    .io_out_8(repl_way_v0_prng_io_out_8),
    .io_out_9(repl_way_v0_prng_io_out_9),
    .io_out_10(repl_way_v0_prng_io_out_10),
    .io_out_11(repl_way_v0_prng_io_out_11),
    .io_out_12(repl_way_v0_prng_io_out_12),
    .io_out_13(repl_way_v0_prng_io_out_13),
    .io_out_14(repl_way_v0_prng_io_out_14),
    .io_out_15(repl_way_v0_prng_io_out_15),
    .io_covSum(repl_way_v0_prng_io_covSum),
    .metaAssert(repl_way_v0_prng_metaAssert),
    .metaReset(repl_way_v0_prng_metaReset)
  );
  assign tag_array_0_tag_rdata_addr = tag_array_0_tag_rdata_addr_pipe_0;
  assign tag_array_0_tag_rdata_data = tag_array_0[tag_array_0_tag_rdata_addr]; // @[DescribedSRAM.scala 19:26]
  assign tag_array_0_MPORT_data = {refillError,refill_tag};
  assign tag_array_0_MPORT_addr = refill_paddr[11:6];
  assign tag_array_0_MPORT_mask = repl_way_v0 == 2'h0;
  assign tag_array_0_MPORT_en = refill_one_beat & d_done;
  assign tag_array_1_tag_rdata_addr = tag_array_1_tag_rdata_addr_pipe_0;
  assign tag_array_1_tag_rdata_data = tag_array_1[tag_array_1_tag_rdata_addr]; // @[DescribedSRAM.scala 19:26]
  assign tag_array_1_MPORT_data = {refillError,refill_tag};
  assign tag_array_1_MPORT_addr = refill_paddr[11:6];
  assign tag_array_1_MPORT_mask = repl_way_v0 == 2'h1;
  assign tag_array_1_MPORT_en = refill_one_beat & d_done;
  assign tag_array_2_tag_rdata_addr = tag_array_2_tag_rdata_addr_pipe_0;
  assign tag_array_2_tag_rdata_data = tag_array_2[tag_array_2_tag_rdata_addr]; // @[DescribedSRAM.scala 19:26]
  assign tag_array_2_MPORT_data = {refillError,refill_tag};
  assign tag_array_2_MPORT_addr = refill_paddr[11:6];
  assign tag_array_2_MPORT_mask = repl_way_v0 == 2'h2;
  assign tag_array_2_MPORT_en = refill_one_beat & d_done;
  assign tag_array_3_tag_rdata_addr = tag_array_3_tag_rdata_addr_pipe_0;
  assign tag_array_3_tag_rdata_data = tag_array_3[tag_array_3_tag_rdata_addr]; // @[DescribedSRAM.scala 19:26]
  assign tag_array_3_MPORT_data = {refillError,refill_tag};
  assign tag_array_3_MPORT_addr = refill_paddr[11:6];
  assign tag_array_3_MPORT_mask = repl_way_v0 == 2'h3;
  assign tag_array_3_MPORT_en = refill_one_beat & d_done;
  assign data_arrays_0_0_dout_addr = data_arrays_0_0_dout_addr_pipe_0;
  assign data_arrays_0_0_dout_data = data_arrays_0_0[data_arrays_0_0_dout_addr]; // @[DescribedSRAM.scala 19:26]
  assign data_arrays_0_0_MPORT_1_data = auto_master_out_d_bits_data[31:0];
  assign data_arrays_0_0_MPORT_1_addr = refill_one_beat ? _mem_idx_T_1 : io_req_bits_addr[11:3];
  assign data_arrays_0_0_MPORT_1_mask = repl_way_v0 == 2'h0;
  assign data_arrays_0_0_MPORT_1_en = refill_one_beat & ~invalidated;
  assign data_arrays_0_1_dout_addr = data_arrays_0_1_dout_addr_pipe_0;
  assign data_arrays_0_1_dout_data = data_arrays_0_1[data_arrays_0_1_dout_addr]; // @[DescribedSRAM.scala 19:26]
  assign data_arrays_0_1_MPORT_1_data = auto_master_out_d_bits_data[31:0];
  assign data_arrays_0_1_MPORT_1_addr = refill_one_beat ? _mem_idx_T_1 : io_req_bits_addr[11:3];
  assign data_arrays_0_1_MPORT_1_mask = repl_way_v0 == 2'h1;
  assign data_arrays_0_1_MPORT_1_en = refill_one_beat & ~invalidated;
  assign data_arrays_0_2_dout_addr = data_arrays_0_2_dout_addr_pipe_0;
  assign data_arrays_0_2_dout_data = data_arrays_0_2[data_arrays_0_2_dout_addr]; // @[DescribedSRAM.scala 19:26]
  assign data_arrays_0_2_MPORT_1_data = auto_master_out_d_bits_data[31:0];
  assign data_arrays_0_2_MPORT_1_addr = refill_one_beat ? _mem_idx_T_1 : io_req_bits_addr[11:3];
  assign data_arrays_0_2_MPORT_1_mask = repl_way_v0 == 2'h2;
  assign data_arrays_0_2_MPORT_1_en = refill_one_beat & ~invalidated;
  assign data_arrays_0_3_dout_addr = data_arrays_0_3_dout_addr_pipe_0;
  assign data_arrays_0_3_dout_data = data_arrays_0_3[data_arrays_0_3_dout_addr]; // @[DescribedSRAM.scala 19:26]
  assign data_arrays_0_3_MPORT_1_data = auto_master_out_d_bits_data[31:0];
  assign data_arrays_0_3_MPORT_1_addr = refill_one_beat ? _mem_idx_T_1 : io_req_bits_addr[11:3];
  assign data_arrays_0_3_MPORT_1_mask = repl_way_v0 == 2'h3;
  assign data_arrays_0_3_MPORT_1_en = refill_one_beat & ~invalidated;
  assign data_arrays_1_0_dout_1_addr = data_arrays_1_0_dout_1_addr_pipe_0;
  assign data_arrays_1_0_dout_1_data = data_arrays_1_0[data_arrays_1_0_dout_1_addr]; // @[DescribedSRAM.scala 19:26]
  assign data_arrays_1_0_MPORT_2_data = auto_master_out_d_bits_data[63:32];
  assign data_arrays_1_0_MPORT_2_addr = refill_one_beat ? _mem_idx_T_1 : io_req_bits_addr[11:3];
  assign data_arrays_1_0_MPORT_2_mask = repl_way_v0 == 2'h0;
  assign data_arrays_1_0_MPORT_2_en = refill_one_beat & ~invalidated;
  assign data_arrays_1_1_dout_1_addr = data_arrays_1_1_dout_1_addr_pipe_0;
  assign data_arrays_1_1_dout_1_data = data_arrays_1_1[data_arrays_1_1_dout_1_addr]; // @[DescribedSRAM.scala 19:26]
  assign data_arrays_1_1_MPORT_2_data = auto_master_out_d_bits_data[63:32];
  assign data_arrays_1_1_MPORT_2_addr = refill_one_beat ? _mem_idx_T_1 : io_req_bits_addr[11:3];
  assign data_arrays_1_1_MPORT_2_mask = repl_way_v0 == 2'h1;
  assign data_arrays_1_1_MPORT_2_en = refill_one_beat & ~invalidated;
  assign data_arrays_1_2_dout_1_addr = data_arrays_1_2_dout_1_addr_pipe_0;
  assign data_arrays_1_2_dout_1_data = data_arrays_1_2[data_arrays_1_2_dout_1_addr]; // @[DescribedSRAM.scala 19:26]
  assign data_arrays_1_2_MPORT_2_data = auto_master_out_d_bits_data[63:32];
  assign data_arrays_1_2_MPORT_2_addr = refill_one_beat ? _mem_idx_T_1 : io_req_bits_addr[11:3];
  assign data_arrays_1_2_MPORT_2_mask = repl_way_v0 == 2'h2;
  assign data_arrays_1_2_MPORT_2_en = refill_one_beat & ~invalidated;
  assign data_arrays_1_3_dout_1_addr = data_arrays_1_3_dout_1_addr_pipe_0;
  assign data_arrays_1_3_dout_1_data = data_arrays_1_3[data_arrays_1_3_dout_1_addr]; // @[DescribedSRAM.scala 19:26]
  assign data_arrays_1_3_MPORT_2_data = auto_master_out_d_bits_data[63:32];
  assign data_arrays_1_3_MPORT_2_addr = refill_one_beat ? _mem_idx_T_1 : io_req_bits_addr[11:3];
  assign data_arrays_1_3_MPORT_2_mask = repl_way_v0 == 2'h3;
  assign data_arrays_1_3_MPORT_2_en = refill_one_beat & ~invalidated;
  assign s0_valid = io_req_ready & io_req_valid; // @[Decoupled.scala 40:37]
  assign s1_vb_lo = io_s1_paddr[11:6]; // @[ICache.scala 486:21]
  assign _s1_vb_T = {1'h0,s1_vb_lo}; // @[Cat.scala 30:58]
  assign _s1_vb_T_1 = vb_array >> _s1_vb_T; // @[ICache.scala 259:25]
  assign s1_vb = _s1_vb_T_1[0]; // @[ICache.scala 259:25]
  assign tag = tag_array_0_tag_rdata_data[19:0]; // @[package.scala 154:13]
  assign s1_tag = io_s1_paddr[31:12]; // @[ICache.scala 254:30]
  assign _tagMatch_T = tag == s1_tag; // @[ICache.scala 262:33]
  assign tagMatch = s1_vb & _tagMatch_T; // @[ICache.scala 262:26]
  assign _s1_vb_T_4 = {1'h1,s1_vb_lo}; // @[Cat.scala 30:58]
  assign _s1_vb_T_5 = vb_array >> _s1_vb_T_4; // @[ICache.scala 259:25]
  assign s1_vb_1 = _s1_vb_T_5[0]; // @[ICache.scala 259:25]
  assign tag_1 = tag_array_1_tag_rdata_data[19:0]; // @[package.scala 154:13]
  assign _tagMatch_T_1 = tag_1 == s1_tag; // @[ICache.scala 262:33]
  assign tagMatch_1 = s1_vb_1 & _tagMatch_T_1; // @[ICache.scala 262:26]
  assign _s1_hit_T = tagMatch | tagMatch_1; // @[ICache.scala 172:35]
  assign _s1_vb_T_8 = {2'h2,s1_vb_lo}; // @[Cat.scala 30:58]
  assign _s1_vb_T_9 = vb_array >> _s1_vb_T_8; // @[ICache.scala 259:25]
  assign s1_vb_2 = _s1_vb_T_9[0]; // @[ICache.scala 259:25]
  assign tag_2 = tag_array_2_tag_rdata_data[19:0]; // @[package.scala 154:13]
  assign _tagMatch_T_2 = tag_2 == s1_tag; // @[ICache.scala 262:33]
  assign tagMatch_2 = s1_vb_2 & _tagMatch_T_2; // @[ICache.scala 262:26]
  assign _s1_hit_T_1 = _s1_hit_T | tagMatch_2; // @[ICache.scala 172:35]
  assign _s1_vb_T_12 = {2'h3,s1_vb_lo}; // @[Cat.scala 30:58]
  assign _s1_vb_T_13 = vb_array >> _s1_vb_T_12; // @[ICache.scala 259:25]
  assign s1_vb_3 = _s1_vb_T_13[0]; // @[ICache.scala 259:25]
  assign tag_3 = tag_array_3_tag_rdata_data[19:0]; // @[package.scala 154:13]
  assign _tagMatch_T_3 = tag_3 == s1_tag; // @[ICache.scala 262:33]
  assign tagMatch_3 = s1_vb_3 & _tagMatch_T_3; // @[ICache.scala 262:26]
  assign _s2_valid_T_1 = s1_valid & ~io_s1_kill; // @[ICache.scala 174:35]
  assign _s2_miss_T_1 = s2_valid & ~s2_hit; // @[ICache.scala 182:26]
  assign s2_miss = _s2_miss_T_1 & ~io_s2_kill; // @[ICache.scala 182:37]
  assign s2_request_refill = s2_miss & s2_request_refill_REG; // @[ICache.scala 184:35]
  assign refill_fire = auto_master_out_a_ready & s2_request_refill; // @[Decoupled.scala 40:37]
  assign _s1_can_request_refill_T = s2_miss | refill_valid; // @[ICache.scala 183:41]
  assign s1_can_request_refill = ~_s1_can_request_refill_T; // @[ICache.scala 183:31]
  assign _refill_paddr_T = s1_valid & s1_can_request_refill; // @[ICache.scala 185:54]
  assign refill_tag = refill_paddr[31:12]; // @[ICache.scala 187:33]
  assign refill_idx = refill_paddr[11:6]; // @[ICache.scala 486:21]
  assign refill_one_beat_opdata = auto_master_out_d_bits_opcode[0]; // @[Edges.scala 105:36]
  assign refill_one_beat = auto_master_out_d_valid & refill_one_beat_opdata; // @[ICache.scala 189:41]
  assign _beats1_decode_T_1 = 27'hfff << auto_master_out_d_bits_size; // @[package.scala 234:77]
  assign beats1_decode = ~_beats1_decode_T_1[11:3]; // @[Edges.scala 219:59]
  assign beats1 = refill_one_beat_opdata ? beats1_decode : 9'h0; // @[Edges.scala 220:14]
  assign counter1 = counter - 9'h1; // @[Edges.scala 229:28]
  assign first = counter == 9'h0; // @[Edges.scala 230:25]
  assign _last_T = counter == 9'h1; // @[Edges.scala 231:25]
  assign _last_T_1 = beats1 == 9'h0; // @[Edges.scala 231:47]
  assign last = _last_T | _last_T_1; // @[Edges.scala 231:37]
  assign d_done = last & auto_master_out_d_valid; // @[Edges.scala 232:22]
  assign refill_cnt = beats1 & ~counter1; // @[Edges.scala 233:25]
  assign refill_done = refill_one_beat & d_done; // @[ICache.scala 195:37]
  assign repl_way_v0_lo = {repl_way_v0_prng_io_out_7,repl_way_v0_prng_io_out_6,repl_way_v0_prng_io_out_5,repl_way_v0_prng_io_out_4,repl_way_v0_prng_io_out_3,repl_way_v0_prng_io_out_2,repl_way_v0_prng_io_out_1,repl_way_v0_prng_io_out_0}; // @[PRNG.scala 86:17]
  assign _repl_way_v0_T = {repl_way_v0_prng_io_out_15,repl_way_v0_prng_io_out_14,repl_way_v0_prng_io_out_13,repl_way_v0_prng_io_out_12,repl_way_v0_prng_io_out_11,repl_way_v0_prng_io_out_10,repl_way_v0_prng_io_out_9,repl_way_v0_prng_io_out_8,repl_way_v0_lo}; // @[PRNG.scala 86:17]
  assign repl_way_v0 = _repl_way_v0_T[1:0]; // @[ICache.scala 201:35]
  assign _repl_way_T = {repl_way_v0,refill_idx}; // @[Cat.scala 30:58]
  assign _refillError_T = refill_cnt > 9'h0; // @[ICache.scala 220:58]
  assign _refillError_T_1 = _refillError_T & accruedRefillError; // @[ICache.scala 220:62]
  assign refillError = auto_master_out_d_bits_corrupt | _refillError_T_1; // @[ICache.scala 220:43]
  assign _vb_array_T_2 = refill_done & ~invalidated; // @[ICache.scala 235:72]
  assign _vb_array_T_3 = 256'h1 << _repl_way_T; // @[ICache.scala 235:32]
  assign _vb_array_T_4 = vb_array | _vb_array_T_3; // @[ICache.scala 235:32]
  assign _vb_array_T_6 = ~vb_array | _vb_array_T_3; // @[ICache.scala 235:32]
  assign s2_tag_disparity = |4'h0; // @[ICache.scala 312:72]
  assign _T_40 = s2_valid & s2_tag_disparity; // @[ICache.scala 334:22]
  assign invalidate = _T_40 | io_invalidate; // @[ICache.scala 334:39]
  assign _GEN_30 = invalidate | invalidated; // @[ICache.scala 238:21]
  assign tl_error = tag_array_0_tag_rdata_data[20]; // @[package.scala 154:13]
  assign s1_tl_error_0 = tagMatch & tl_error; // @[ICache.scala 264:32]
  assign tl_error_1 = tag_array_1_tag_rdata_data[20]; // @[package.scala 154:13]
  assign s1_tl_error_1 = tagMatch_1 & tl_error_1; // @[ICache.scala 264:32]
  assign tl_error_2 = tag_array_2_tag_rdata_data[20]; // @[package.scala 154:13]
  assign s1_tl_error_2 = tagMatch_2 & tl_error_2; // @[ICache.scala 264:32]
  assign tl_error_3 = tag_array_3_tag_rdata_data[20]; // @[package.scala 154:13]
  assign s1_tl_error_3 = tagMatch_3 & tl_error_3; // @[ICache.scala 264:32]
  assign _T_15 = tagMatch + tagMatch_1; // @[Bitwise.scala 47:55]
  assign _T_17 = tagMatch_2 + tagMatch_3; // @[Bitwise.scala 47:55]
  assign _T_19 = _T_15 + _T_17; // @[Bitwise.scala 47:55]
  assign _T_21 = _T_19 <= 3'h1; // @[ICache.scala 267:115]
  assign _T_22 = ~s1_valid | _T_21; // @[ICache.scala 267:39]
  assign _T_24 = _T_22 | reset; // @[ICache.scala 267:9]
  assign s0_ren = s0_valid & ~io_req_bits_addr[2]; // @[ICache.scala 284:28]
  assign wen = refill_one_beat & ~invalidated; // @[ICache.scala 285:32]
  assign _mem_idx_T = {refill_idx, 3'h0}; // @[ICache.scala 286:52]
  assign _mem_idx_T_1 = _mem_idx_T | refill_cnt; // @[ICache.scala 286:79]
  assign _GEN_54 = data_arrays_0_0_dout_data; // @[ICache.scala 296:71]
  assign _GEN_55 = data_arrays_0_1_dout_data; // @[ICache.scala 296:71]
  assign _GEN_56 = data_arrays_0_2_dout_data; // @[ICache.scala 296:71]
  assign _GEN_57 = data_arrays_0_3_dout_data; // @[ICache.scala 296:71]
  assign s0_ren_1 = s0_valid & io_req_bits_addr[2]; // @[ICache.scala 284:28]
  assign _s2_way_mux_T = s2_tag_hit_0 ? s2_dout_0 : 32'h0; // @[Mux.scala 27:72]
  assign _s2_way_mux_T_1 = s2_tag_hit_1 ? s2_dout_1 : 32'h0; // @[Mux.scala 27:72]
  assign _s2_way_mux_T_2 = s2_tag_hit_2 ? s2_dout_2 : 32'h0; // @[Mux.scala 27:72]
  assign _s2_way_mux_T_3 = s2_tag_hit_3 ? s2_dout_3 : 32'h0; // @[Mux.scala 27:72]
  assign _s2_way_mux_T_4 = _s2_way_mux_T | _s2_way_mux_T_1; // @[Mux.scala 27:72]
  assign _s2_way_mux_T_5 = _s2_way_mux_T_4 | _s2_way_mux_T_2; // @[Mux.scala 27:72]
  assign _s2_tl_error_T = {s1_tl_error_3,s1_tl_error_2,s1_tl_error_1,s1_tl_error_0}; // @[ICache.scala 313:43]
  assign _s2_tl_error_T_1 = |_s2_tl_error_T; // @[ICache.scala 313:50]
  assign _GEN_101 = refill_fire | refill_valid; // @[ICache.scala 477:22]
  assign auto_master_out_a_valid = s2_miss & s2_request_refill_REG; // @[LazyModule.scala 311:12]
  assign auto_master_out_a_bits_address = {refill_paddr[31:6], 6'h0}; // @[LazyModule.scala 311:12]
  assign io_req_ready = ~refill_one_beat; // @[ICache.scala 191:16]
  assign io_resp_valid = s2_valid & s2_hit; // @[ICache.scala 339:21]
  assign io_resp_bits_data = _s2_way_mux_T_5 | _s2_way_mux_T_3; // @[ICache.scala 336:25]
  assign io_resp_bits_replay = |4'h0; // @[ICache.scala 338:27]
  assign io_resp_bits_ae = s2_tl_error; // @[ICache.scala 337:23]
  assign repl_way_v0_prng_clock = clock;
  assign repl_way_v0_prng_reset = reset;
  assign repl_way_v0_prng_io_increment = auto_master_out_a_ready & s2_request_refill; // @[PRNG.scala 85:23]
  assign ICache_cov_read_addr = ICache_state;
  assign ICache_cov_read_data = ICache_cov[ICache_cov_read_addr]; // @[Coverage map for ICache]
  assign ICache_cov_write_data = 1'h1;
  assign ICache_cov_write_addr = ICache_state;
  assign ICache_cov_write_mask = 1'h1;
  assign ICache_cov_write_en = 1'h1;
  assign s2_valid_shl = s2_valid;
  assign s2_valid_pad = {5'h0,s2_valid_shl};
  assign s1_valid_shl = {s1_valid, 1'h0};
  assign s1_valid_pad = {4'h0,s1_valid_shl};
  assign refill_valid_shl = {refill_valid, 2'h0};
  assign refill_valid_pad = {3'h0,refill_valid_shl};
  assign invalidated_shl = {invalidated, 3'h0};
  assign invalidated_pad = {2'h0,invalidated_shl};
  assign s2_hit_shl = {s2_hit, 4'h0};
  assign s2_hit_pad = {1'h0,s2_hit_shl};
  assign s2_tag_hit_0_shl = {s2_tag_hit_0, 5'h0};
  assign s2_tag_hit_0_pad = s2_tag_hit_0_shl;
  assign s2_tag_hit_1_shl = {s2_tag_hit_1, 5'h0};
  assign s2_tag_hit_1_pad = s2_tag_hit_1_shl;
  assign s2_tag_hit_2_shl = {s2_tag_hit_2, 5'h0};
  assign s2_tag_hit_2_pad = s2_tag_hit_2_shl;
  assign s2_tag_hit_3_shl = {s2_tag_hit_3, 5'h0};
  assign s2_tag_hit_3_pad = s2_tag_hit_3_shl;
  assign ICache_xor3 = s2_valid_pad ^ s1_valid_pad;
  assign ICache_xor4 = refill_valid_pad ^ invalidated_pad;
  assign ICache_xor1 = ICache_xor3 ^ ICache_xor4;
  assign ICache_xor5 = s2_hit_pad ^ s2_tag_hit_0_pad;
  assign ICache_xor14 = s2_tag_hit_2_pad ^ s2_tag_hit_3_pad;
  assign ICache_xor6 = s2_tag_hit_1_pad ^ ICache_xor14;
  assign ICache_xor2 = ICache_xor5 ^ ICache_xor6;
  assign ICache_xor0 = ICache_xor1 ^ ICache_xor2;
  assign repl_way_v0_prng_sum = ICache_covSum + repl_way_v0_prng_io_covSum;
  assign io_covSum = repl_way_v0_prng_sum;
  assign stopEn0 = ~_T_24;
  assign repl_way_v0_prng_metaAssert_wire = repl_way_v0_prng_metaAssert;
  assign ICache_or0 = stopEn0 | repl_way_v0_prng_metaAssert_wire;
  assign metaAssert = ICache_metaAssert;
  assign repl_way_v0_prng_metaReset = metaReset | repl_way_v0_prng_halt;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tag_array_0[initvar] = _RAND_0[20:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  tag_array_0_tag_rdata_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  tag_array_0_tag_rdata_addr_pipe_0 = _RAND_2[5:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tag_array_1[initvar] = _RAND_3[20:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  tag_array_1_tag_rdata_en_pipe_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  tag_array_1_tag_rdata_addr_pipe_0 = _RAND_5[5:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tag_array_2[initvar] = _RAND_6[20:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  tag_array_2_tag_rdata_en_pipe_0 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  tag_array_2_tag_rdata_addr_pipe_0 = _RAND_8[5:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tag_array_3[initvar] = _RAND_9[20:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  tag_array_3_tag_rdata_en_pipe_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  tag_array_3_tag_rdata_addr_pipe_0 = _RAND_11[5:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_0[initvar] = _RAND_12[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  data_arrays_0_0_dout_en_pipe_0 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  data_arrays_0_0_dout_addr_pipe_0 = _RAND_14[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_1[initvar] = _RAND_15[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  data_arrays_0_1_dout_en_pipe_0 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  data_arrays_0_1_dout_addr_pipe_0 = _RAND_17[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_2[initvar] = _RAND_18[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  data_arrays_0_2_dout_en_pipe_0 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  data_arrays_0_2_dout_addr_pipe_0 = _RAND_20[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_0_3[initvar] = _RAND_21[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  data_arrays_0_3_dout_en_pipe_0 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  data_arrays_0_3_dout_addr_pipe_0 = _RAND_23[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_1_0[initvar] = _RAND_24[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  data_arrays_1_0_dout_1_en_pipe_0 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  data_arrays_1_0_dout_1_addr_pipe_0 = _RAND_26[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_1_1[initvar] = _RAND_27[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  data_arrays_1_1_dout_1_en_pipe_0 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  data_arrays_1_1_dout_1_addr_pipe_0 = _RAND_29[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_1_2[initvar] = _RAND_30[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  data_arrays_1_2_dout_1_en_pipe_0 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  data_arrays_1_2_dout_1_addr_pipe_0 = _RAND_32[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    data_arrays_1_3[initvar] = _RAND_33[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  data_arrays_1_3_dout_1_en_pipe_0 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  data_arrays_1_3_dout_1_addr_pipe_0 = _RAND_35[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  s1_valid = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {8{`RANDOM}};
  vb_array = _RAND_37[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  s2_valid = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  s2_hit = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  invalidated = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  refill_valid = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  s2_request_refill_REG = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  refill_paddr = _RAND_43[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  counter = _RAND_44[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  accruedRefillError = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  s2_tag_hit_0 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  s2_tag_hit_1 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  s2_tag_hit_2 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  s2_tag_hit_3 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  s2_dout_0 = _RAND_50[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  s2_dout_1 = _RAND_51[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  s2_dout_2 = _RAND_52[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  s2_dout_3 = _RAND_53[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  s2_tl_error = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  ICache_state = _RAND_55[5:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    ICache_cov[initvar] = _RAND_56[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  ICache_covSum = _RAND_57[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  ICache_metaAssert = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(tag_array_0_MPORT_en & tag_array_0_MPORT_mask) begin
      tag_array_0[tag_array_0_MPORT_addr] <= tag_array_0_MPORT_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      tag_array_0_tag_rdata_en_pipe_0 <= 1'h0;
    end else begin
      tag_array_0_tag_rdata_en_pipe_0 <= ~refill_done & s0_valid;
    end
    if (metaReset) begin
      tag_array_0_tag_rdata_addr_pipe_0 <= 6'h0;
    end else if (~refill_done & s0_valid) begin
      tag_array_0_tag_rdata_addr_pipe_0 <= io_req_bits_addr[11:6];
    end
    if(tag_array_1_MPORT_en & tag_array_1_MPORT_mask) begin
      tag_array_1[tag_array_1_MPORT_addr] <= tag_array_1_MPORT_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      tag_array_1_tag_rdata_en_pipe_0 <= 1'h0;
    end else begin
      tag_array_1_tag_rdata_en_pipe_0 <= ~refill_done & s0_valid;
    end
    if (metaReset) begin
      tag_array_1_tag_rdata_addr_pipe_0 <= 6'h0;
    end else if (~refill_done & s0_valid) begin
      tag_array_1_tag_rdata_addr_pipe_0 <= io_req_bits_addr[11:6];
    end
    if(tag_array_2_MPORT_en & tag_array_2_MPORT_mask) begin
      tag_array_2[tag_array_2_MPORT_addr] <= tag_array_2_MPORT_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      tag_array_2_tag_rdata_en_pipe_0 <= 1'h0;
    end else begin
      tag_array_2_tag_rdata_en_pipe_0 <= ~refill_done & s0_valid;
    end
    if (metaReset) begin
      tag_array_2_tag_rdata_addr_pipe_0 <= 6'h0;
    end else if (~refill_done & s0_valid) begin
      tag_array_2_tag_rdata_addr_pipe_0 <= io_req_bits_addr[11:6];
    end
    if(tag_array_3_MPORT_en & tag_array_3_MPORT_mask) begin
      tag_array_3[tag_array_3_MPORT_addr] <= tag_array_3_MPORT_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      tag_array_3_tag_rdata_en_pipe_0 <= 1'h0;
    end else begin
      tag_array_3_tag_rdata_en_pipe_0 <= ~refill_done & s0_valid;
    end
    if (metaReset) begin
      tag_array_3_tag_rdata_addr_pipe_0 <= 6'h0;
    end else if (~refill_done & s0_valid) begin
      tag_array_3_tag_rdata_addr_pipe_0 <= io_req_bits_addr[11:6];
    end
    if(data_arrays_0_0_MPORT_1_en & data_arrays_0_0_MPORT_1_mask) begin
      data_arrays_0_0[data_arrays_0_0_MPORT_1_addr] <= data_arrays_0_0_MPORT_1_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      data_arrays_0_0_dout_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_0_dout_en_pipe_0 <= ~wen & s0_ren;
    end
    if (metaReset) begin
      data_arrays_0_0_dout_addr_pipe_0 <= 9'h0;
    end else if (~wen & s0_ren) begin
      if (refill_one_beat) begin
        data_arrays_0_0_dout_addr_pipe_0 <= _mem_idx_T_1;
      end else begin
        data_arrays_0_0_dout_addr_pipe_0 <= io_req_bits_addr[11:3];
      end
    end
    if(data_arrays_0_1_MPORT_1_en & data_arrays_0_1_MPORT_1_mask) begin
      data_arrays_0_1[data_arrays_0_1_MPORT_1_addr] <= data_arrays_0_1_MPORT_1_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      data_arrays_0_1_dout_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_1_dout_en_pipe_0 <= ~wen & s0_ren;
    end
    if (metaReset) begin
      data_arrays_0_1_dout_addr_pipe_0 <= 9'h0;
    end else if (~wen & s0_ren) begin
      if (refill_one_beat) begin
        data_arrays_0_1_dout_addr_pipe_0 <= _mem_idx_T_1;
      end else begin
        data_arrays_0_1_dout_addr_pipe_0 <= io_req_bits_addr[11:3];
      end
    end
    if(data_arrays_0_2_MPORT_1_en & data_arrays_0_2_MPORT_1_mask) begin
      data_arrays_0_2[data_arrays_0_2_MPORT_1_addr] <= data_arrays_0_2_MPORT_1_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      data_arrays_0_2_dout_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_2_dout_en_pipe_0 <= ~wen & s0_ren;
    end
    if (metaReset) begin
      data_arrays_0_2_dout_addr_pipe_0 <= 9'h0;
    end else if (~wen & s0_ren) begin
      if (refill_one_beat) begin
        data_arrays_0_2_dout_addr_pipe_0 <= _mem_idx_T_1;
      end else begin
        data_arrays_0_2_dout_addr_pipe_0 <= io_req_bits_addr[11:3];
      end
    end
    if(data_arrays_0_3_MPORT_1_en & data_arrays_0_3_MPORT_1_mask) begin
      data_arrays_0_3[data_arrays_0_3_MPORT_1_addr] <= data_arrays_0_3_MPORT_1_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      data_arrays_0_3_dout_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_0_3_dout_en_pipe_0 <= ~wen & s0_ren;
    end
    if (metaReset) begin
      data_arrays_0_3_dout_addr_pipe_0 <= 9'h0;
    end else if (~wen & s0_ren) begin
      if (refill_one_beat) begin
        data_arrays_0_3_dout_addr_pipe_0 <= _mem_idx_T_1;
      end else begin
        data_arrays_0_3_dout_addr_pipe_0 <= io_req_bits_addr[11:3];
      end
    end
    if(data_arrays_1_0_MPORT_2_en & data_arrays_1_0_MPORT_2_mask) begin
      data_arrays_1_0[data_arrays_1_0_MPORT_2_addr] <= data_arrays_1_0_MPORT_2_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      data_arrays_1_0_dout_1_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_1_0_dout_1_en_pipe_0 <= ~wen & s0_ren_1;
    end
    if (metaReset) begin
      data_arrays_1_0_dout_1_addr_pipe_0 <= 9'h0;
    end else if (~wen & s0_ren_1) begin
      if (refill_one_beat) begin
        data_arrays_1_0_dout_1_addr_pipe_0 <= _mem_idx_T_1;
      end else begin
        data_arrays_1_0_dout_1_addr_pipe_0 <= io_req_bits_addr[11:3];
      end
    end
    if(data_arrays_1_1_MPORT_2_en & data_arrays_1_1_MPORT_2_mask) begin
      data_arrays_1_1[data_arrays_1_1_MPORT_2_addr] <= data_arrays_1_1_MPORT_2_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      data_arrays_1_1_dout_1_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_1_1_dout_1_en_pipe_0 <= ~wen & s0_ren_1;
    end
    if (metaReset) begin
      data_arrays_1_1_dout_1_addr_pipe_0 <= 9'h0;
    end else if (~wen & s0_ren_1) begin
      if (refill_one_beat) begin
        data_arrays_1_1_dout_1_addr_pipe_0 <= _mem_idx_T_1;
      end else begin
        data_arrays_1_1_dout_1_addr_pipe_0 <= io_req_bits_addr[11:3];
      end
    end
    if(data_arrays_1_2_MPORT_2_en & data_arrays_1_2_MPORT_2_mask) begin
      data_arrays_1_2[data_arrays_1_2_MPORT_2_addr] <= data_arrays_1_2_MPORT_2_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      data_arrays_1_2_dout_1_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_1_2_dout_1_en_pipe_0 <= ~wen & s0_ren_1;
    end
    if (metaReset) begin
      data_arrays_1_2_dout_1_addr_pipe_0 <= 9'h0;
    end else if (~wen & s0_ren_1) begin
      if (refill_one_beat) begin
        data_arrays_1_2_dout_1_addr_pipe_0 <= _mem_idx_T_1;
      end else begin
        data_arrays_1_2_dout_1_addr_pipe_0 <= io_req_bits_addr[11:3];
      end
    end
    if(data_arrays_1_3_MPORT_2_en & data_arrays_1_3_MPORT_2_mask) begin
      data_arrays_1_3[data_arrays_1_3_MPORT_2_addr] <= data_arrays_1_3_MPORT_2_data; // @[DescribedSRAM.scala 19:26]
    end
    if (metaReset) begin
      data_arrays_1_3_dout_1_en_pipe_0 <= 1'h0;
    end else begin
      data_arrays_1_3_dout_1_en_pipe_0 <= ~wen & s0_ren_1;
    end
    if (metaReset) begin
      data_arrays_1_3_dout_1_addr_pipe_0 <= 9'h0;
    end else if (~wen & s0_ren_1) begin
      if (refill_one_beat) begin
        data_arrays_1_3_dout_1_addr_pipe_0 <= _mem_idx_T_1;
      end else begin
        data_arrays_1_3_dout_1_addr_pipe_0 <= io_req_bits_addr[11:3];
      end
    end
    if (metaReset) begin
      s1_valid <= 1'h0;
    end else if (reset) begin
      s1_valid <= 1'h0;
    end else begin
      s1_valid <= s0_valid;
    end
    if (metaReset) begin
      vb_array <= 256'h0;
    end else if (reset) begin
      vb_array <= 256'h0;
    end else if (invalidate) begin
      vb_array <= 256'h0;
    end else if (refill_one_beat) begin
      if (_vb_array_T_2) begin
        vb_array <= _vb_array_T_4;
      end else begin
        vb_array <= ~_vb_array_T_6;
      end
    end
    if (metaReset) begin
      s2_valid <= 1'h0;
    end else if (reset) begin
      s2_valid <= 1'h0;
    end else begin
      s2_valid <= _s2_valid_T_1;
    end
    if (metaReset) begin
      s2_hit <= 1'h0;
    end else begin
      s2_hit <= _s1_hit_T_1 | tagMatch_3;
    end
    if (metaReset) begin
      invalidated <= 1'h0;
    end else if (~refill_valid) begin
      invalidated <= 1'h0;
    end else begin
      invalidated <= _GEN_30;
    end
    if (metaReset) begin
      refill_valid <= 1'h0;
    end else if (reset) begin
      refill_valid <= 1'h0;
    end else if (refill_done) begin
      refill_valid <= 1'h0;
    end else begin
      refill_valid <= _GEN_101;
    end
    if (metaReset) begin
      s2_request_refill_REG <= 1'h0;
    end else begin
      s2_request_refill_REG <= ~_s1_can_request_refill_T;
    end
    if (metaReset) begin
      refill_paddr <= 32'h0;
    end else if (_refill_paddr_T) begin
      refill_paddr <= io_s1_paddr;
    end
    if (metaReset) begin
      counter <= 9'h0;
    end else if (reset) begin
      counter <= 9'h0;
    end else if (auto_master_out_d_valid) begin
      if (first) begin
        if (refill_one_beat_opdata) begin
          counter <= beats1_decode;
        end else begin
          counter <= 9'h0;
        end
      end else begin
        counter <= counter1;
      end
    end
    if (metaReset) begin
      accruedRefillError <= 1'h0;
    end else if (refill_one_beat) begin
      accruedRefillError <= refillError;
    end
    if (metaReset) begin
      s2_tag_hit_0 <= 1'h0;
    end else if (s1_valid) begin
      s2_tag_hit_0 <= tagMatch;
    end
    if (metaReset) begin
      s2_tag_hit_1 <= 1'h0;
    end else if (s1_valid) begin
      s2_tag_hit_1 <= tagMatch_1;
    end
    if (metaReset) begin
      s2_tag_hit_2 <= 1'h0;
    end else if (s1_valid) begin
      s2_tag_hit_2 <= tagMatch_2;
    end
    if (metaReset) begin
      s2_tag_hit_3 <= 1'h0;
    end else if (s1_valid) begin
      s2_tag_hit_3 <= tagMatch_3;
    end
    if (metaReset) begin
      s2_dout_0 <= 32'h0;
    end else if (s1_valid) begin
      if (io_s1_paddr[2]) begin
        s2_dout_0 <= data_arrays_1_0_dout_1_data;
      end else begin
        s2_dout_0 <= _GEN_54;
      end
    end
    if (metaReset) begin
      s2_dout_1 <= 32'h0;
    end else if (s1_valid) begin
      if (io_s1_paddr[2]) begin
        s2_dout_1 <= data_arrays_1_1_dout_1_data;
      end else begin
        s2_dout_1 <= _GEN_55;
      end
    end
    if (metaReset) begin
      s2_dout_2 <= 32'h0;
    end else if (s1_valid) begin
      if (io_s1_paddr[2]) begin
        s2_dout_2 <= data_arrays_1_2_dout_1_data;
      end else begin
        s2_dout_2 <= _GEN_56;
      end
    end
    if (metaReset) begin
      s2_dout_3 <= 32'h0;
    end else if (s1_valid) begin
      if (io_s1_paddr[2]) begin
        s2_dout_3 <= data_arrays_1_3_dout_1_data;
      end else begin
        s2_dout_3 <= _GEN_57;
      end
    end
    if (metaReset) begin
      s2_tl_error <= 1'h0;
    end else if (s1_valid) begin
      s2_tl_error <= _s2_tl_error_T_1;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_24) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ICache.scala:267 assert(!(s1_valid || s1_slaveValid) || PopCount(s1_tag_hit zip s1_tag_disparity map { case (h, d) => h && !d }) <= 1)\n"); // @[ICache.scala 267:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_24) begin
          $fatal; // @[ICache.scala 267:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    ICache_state <= ICache_xor0;
    if (!(ICache_cov_read_data)) begin
      ICache_covSum <= ICache_covSum + 1'h1;
    end
    if (metaReset) begin
      ICache_metaAssert <= 1'h0;
    end else begin
      ICache_metaAssert <= ICache_metaAssert | ICache_or0;
    end
  end
  always @(posedge clock) begin
    if(ICache_cov_write_en & ICache_cov_write_mask) begin
      ICache_cov[ICache_cov_write_addr] <= ICache_cov_write_data; // @[Coverage map for ICache]
    end
  end
endmodule
module ShiftQueue(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_btb_taken,
  input         io_enq_bits_btb_bridx,
  input  [4:0]  io_enq_bits_btb_entry,
  input  [7:0]  io_enq_bits_btb_bht_history,
  input  [39:0] io_enq_bits_pc,
  input  [31:0] io_enq_bits_data,
  input  [1:0]  io_enq_bits_mask,
  input         io_enq_bits_xcpt_pf_inst,
  input         io_enq_bits_xcpt_ae_inst,
  input         io_enq_bits_replay,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_btb_taken,
  output        io_deq_bits_btb_bridx,
  output [4:0]  io_deq_bits_btb_entry,
  output [7:0]  io_deq_bits_btb_bht_history,
  output [39:0] io_deq_bits_pc,
  output [31:0] io_deq_bits_data,
  output        io_deq_bits_xcpt_pf_inst,
  output        io_deq_bits_xcpt_ae_inst,
  output        io_deq_bits_replay,
  output [4:0]  io_mask,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  reg  valid_0; // @[ShiftQueue.scala 21:30]
  reg [31:0] _RAND_0;
  reg  valid_1; // @[ShiftQueue.scala 21:30]
  reg [31:0] _RAND_1;
  reg  valid_2; // @[ShiftQueue.scala 21:30]
  reg [31:0] _RAND_2;
  reg  valid_3; // @[ShiftQueue.scala 21:30]
  reg [31:0] _RAND_3;
  reg  valid_4; // @[ShiftQueue.scala 21:30]
  reg [31:0] _RAND_4;
  reg  elts_0_btb_taken; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_5;
  reg  elts_0_btb_bridx; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_6;
  reg [4:0] elts_0_btb_entry; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_7;
  reg [7:0] elts_0_btb_bht_history; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_8;
  reg [39:0] elts_0_pc; // @[ShiftQueue.scala 22:25]
  reg [63:0] _RAND_9;
  reg [31:0] elts_0_data; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_10;
  reg  elts_0_xcpt_pf_inst; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_11;
  reg  elts_0_xcpt_ae_inst; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_12;
  reg  elts_0_replay; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_13;
  reg  elts_1_btb_taken; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_14;
  reg  elts_1_btb_bridx; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_15;
  reg [4:0] elts_1_btb_entry; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_16;
  reg [7:0] elts_1_btb_bht_history; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_17;
  reg [39:0] elts_1_pc; // @[ShiftQueue.scala 22:25]
  reg [63:0] _RAND_18;
  reg [31:0] elts_1_data; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_19;
  reg  elts_1_xcpt_pf_inst; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_20;
  reg  elts_1_xcpt_ae_inst; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_21;
  reg  elts_1_replay; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_22;
  reg  elts_2_btb_taken; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_23;
  reg  elts_2_btb_bridx; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_24;
  reg [4:0] elts_2_btb_entry; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_25;
  reg [7:0] elts_2_btb_bht_history; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_26;
  reg [39:0] elts_2_pc; // @[ShiftQueue.scala 22:25]
  reg [63:0] _RAND_27;
  reg [31:0] elts_2_data; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_28;
  reg  elts_2_xcpt_pf_inst; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_29;
  reg  elts_2_xcpt_ae_inst; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_30;
  reg  elts_2_replay; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_31;
  reg  elts_3_btb_taken; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_32;
  reg  elts_3_btb_bridx; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_33;
  reg [4:0] elts_3_btb_entry; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_34;
  reg [7:0] elts_3_btb_bht_history; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_35;
  reg [39:0] elts_3_pc; // @[ShiftQueue.scala 22:25]
  reg [63:0] _RAND_36;
  reg [31:0] elts_3_data; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_37;
  reg  elts_3_xcpt_pf_inst; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_38;
  reg  elts_3_xcpt_ae_inst; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_39;
  reg  elts_3_replay; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_40;
  reg  elts_4_btb_taken; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_41;
  reg  elts_4_btb_bridx; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_42;
  reg [4:0] elts_4_btb_entry; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_43;
  reg [7:0] elts_4_btb_bht_history; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_44;
  reg [39:0] elts_4_pc; // @[ShiftQueue.scala 22:25]
  reg [63:0] _RAND_45;
  reg [31:0] elts_4_data; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_46;
  reg  elts_4_xcpt_pf_inst; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_47;
  reg  elts_4_xcpt_ae_inst; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_48;
  reg  elts_4_replay; // @[ShiftQueue.scala 22:25]
  reg [31:0] _RAND_49;
  wire  _wen_T; // @[Decoupled.scala 40:37]
  wire  _wen_T_2; // @[ShiftQueue.scala 30:45]
  wire  _wen_T_3; // @[ShiftQueue.scala 30:28]
  wire  _wen_T_7; // @[ShiftQueue.scala 31:45]
  wire  wen; // @[ShiftQueue.scala 29:10]
  wire  _valid_0_T_6; // @[ShiftQueue.scala 37:45]
  wire  _wen_T_10; // @[ShiftQueue.scala 30:45]
  wire  _wen_T_11; // @[ShiftQueue.scala 30:28]
  wire  _wen_T_15; // @[ShiftQueue.scala 31:45]
  wire  wen_1; // @[ShiftQueue.scala 29:10]
  wire  _valid_1_T_6; // @[ShiftQueue.scala 37:45]
  wire  _wen_T_18; // @[ShiftQueue.scala 30:45]
  wire  _wen_T_19; // @[ShiftQueue.scala 30:28]
  wire  _wen_T_23; // @[ShiftQueue.scala 31:45]
  wire  wen_2; // @[ShiftQueue.scala 29:10]
  wire  _valid_2_T_6; // @[ShiftQueue.scala 37:45]
  wire  _wen_T_26; // @[ShiftQueue.scala 30:45]
  wire  _wen_T_27; // @[ShiftQueue.scala 30:28]
  wire  _wen_T_31; // @[ShiftQueue.scala 31:45]
  wire  wen_3; // @[ShiftQueue.scala 29:10]
  wire  _valid_3_T_6; // @[ShiftQueue.scala 37:45]
  wire  _wen_T_34; // @[ShiftQueue.scala 30:45]
  wire  _wen_T_39; // @[ShiftQueue.scala 31:45]
  wire  wen_4; // @[ShiftQueue.scala 29:10]
  wire  _valid_4_T_6; // @[ShiftQueue.scala 37:45]
  wire [1:0] io_mask_lo; // @[ShiftQueue.scala 53:20]
  wire [2:0] io_mask_hi; // @[ShiftQueue.scala 53:20]
  reg  ShiftQueue_state; // @[Register tracking ShiftQueue state]
  reg [31:0] _RAND_50;
  reg  ShiftQueue_cov [0:1]; // @[Coverage map for ShiftQueue]
  reg [31:0] _RAND_51;
  wire  ShiftQueue_cov_read_data; // @[Coverage map for ShiftQueue]
  wire  ShiftQueue_cov_read_addr; // @[Coverage map for ShiftQueue]
  wire  ShiftQueue_cov_write_data; // @[Coverage map for ShiftQueue]
  wire  ShiftQueue_cov_write_addr; // @[Coverage map for ShiftQueue]
  wire  ShiftQueue_cov_write_mask; // @[Coverage map for ShiftQueue]
  wire  ShiftQueue_cov_write_en; // @[Coverage map for ShiftQueue]
  reg [29:0] ShiftQueue_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_52;
  wire  valid_1_shl;
  wire  valid_1_pad;
  wire  valid_0_shl;
  wire  valid_0_pad;
  wire  valid_2_shl;
  wire  valid_2_pad;
  wire  valid_4_shl;
  wire  valid_4_pad;
  wire  valid_3_shl;
  wire  valid_3_pad;
  wire  ShiftQueue_xor1;
  wire  ShiftQueue_xor6;
  wire  ShiftQueue_xor2;
  wire  ShiftQueue_xor0;
  assign _wen_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _wen_T_2 = _wen_T & valid_0; // @[ShiftQueue.scala 30:45]
  assign _wen_T_3 = valid_1 | _wen_T_2; // @[ShiftQueue.scala 30:28]
  assign _wen_T_7 = _wen_T & ~valid_0; // @[ShiftQueue.scala 31:45]
  assign wen = io_deq_ready ? _wen_T_3 : _wen_T_7; // @[ShiftQueue.scala 29:10]
  assign _valid_0_T_6 = _wen_T | valid_0; // @[ShiftQueue.scala 37:45]
  assign _wen_T_10 = _wen_T & valid_1; // @[ShiftQueue.scala 30:45]
  assign _wen_T_11 = valid_2 | _wen_T_10; // @[ShiftQueue.scala 30:28]
  assign _wen_T_15 = _wen_T_2 & ~valid_1; // @[ShiftQueue.scala 31:45]
  assign wen_1 = io_deq_ready ? _wen_T_11 : _wen_T_15; // @[ShiftQueue.scala 29:10]
  assign _valid_1_T_6 = _wen_T_2 | valid_1; // @[ShiftQueue.scala 37:45]
  assign _wen_T_18 = _wen_T & valid_2; // @[ShiftQueue.scala 30:45]
  assign _wen_T_19 = valid_3 | _wen_T_18; // @[ShiftQueue.scala 30:28]
  assign _wen_T_23 = _wen_T_10 & ~valid_2; // @[ShiftQueue.scala 31:45]
  assign wen_2 = io_deq_ready ? _wen_T_19 : _wen_T_23; // @[ShiftQueue.scala 29:10]
  assign _valid_2_T_6 = _wen_T_10 | valid_2; // @[ShiftQueue.scala 37:45]
  assign _wen_T_26 = _wen_T & valid_3; // @[ShiftQueue.scala 30:45]
  assign _wen_T_27 = valid_4 | _wen_T_26; // @[ShiftQueue.scala 30:28]
  assign _wen_T_31 = _wen_T_18 & ~valid_3; // @[ShiftQueue.scala 31:45]
  assign wen_3 = io_deq_ready ? _wen_T_27 : _wen_T_31; // @[ShiftQueue.scala 29:10]
  assign _valid_3_T_6 = _wen_T_18 | valid_3; // @[ShiftQueue.scala 37:45]
  assign _wen_T_34 = _wen_T & valid_4; // @[ShiftQueue.scala 30:45]
  assign _wen_T_39 = _wen_T_26 & ~valid_4; // @[ShiftQueue.scala 31:45]
  assign wen_4 = io_deq_ready ? _wen_T_34 : _wen_T_39; // @[ShiftQueue.scala 29:10]
  assign _valid_4_T_6 = _wen_T_26 | valid_4; // @[ShiftQueue.scala 37:45]
  assign io_mask_lo = {valid_1,valid_0}; // @[ShiftQueue.scala 53:20]
  assign io_mask_hi = {valid_4,valid_3,valid_2}; // @[ShiftQueue.scala 53:20]
  assign io_enq_ready = ~valid_4; // @[ShiftQueue.scala 40:16]
  assign io_deq_valid = io_enq_valid | valid_0; // @[ShiftQueue.scala 41:16 ShiftQueue.scala 45:40]
  assign io_deq_bits_btb_taken = valid_0 ? elts_0_btb_taken : io_enq_bits_btb_taken; // @[ShiftQueue.scala 42:15 ShiftQueue.scala 46:36]
  assign io_deq_bits_btb_bridx = valid_0 ? elts_0_btb_bridx : io_enq_bits_btb_bridx; // @[ShiftQueue.scala 42:15 ShiftQueue.scala 46:36]
  assign io_deq_bits_btb_entry = valid_0 ? elts_0_btb_entry : io_enq_bits_btb_entry; // @[ShiftQueue.scala 42:15 ShiftQueue.scala 46:36]
  assign io_deq_bits_btb_bht_history = valid_0 ? elts_0_btb_bht_history : io_enq_bits_btb_bht_history; // @[ShiftQueue.scala 42:15 ShiftQueue.scala 46:36]
  assign io_deq_bits_pc = valid_0 ? elts_0_pc : io_enq_bits_pc; // @[ShiftQueue.scala 42:15 ShiftQueue.scala 46:36]
  assign io_deq_bits_data = valid_0 ? elts_0_data : io_enq_bits_data; // @[ShiftQueue.scala 42:15 ShiftQueue.scala 46:36]
  assign io_deq_bits_xcpt_pf_inst = valid_0 ? elts_0_xcpt_pf_inst : io_enq_bits_xcpt_pf_inst; // @[ShiftQueue.scala 42:15 ShiftQueue.scala 46:36]
  assign io_deq_bits_xcpt_ae_inst = valid_0 ? elts_0_xcpt_ae_inst : io_enq_bits_xcpt_ae_inst; // @[ShiftQueue.scala 42:15 ShiftQueue.scala 46:36]
  assign io_deq_bits_replay = valid_0 ? elts_0_replay : io_enq_bits_replay; // @[ShiftQueue.scala 42:15 ShiftQueue.scala 46:36]
  assign io_mask = {io_mask_hi,io_mask_lo}; // @[ShiftQueue.scala 53:11]
  assign ShiftQueue_cov_read_addr = ShiftQueue_state;
  assign ShiftQueue_cov_read_data = ShiftQueue_cov[ShiftQueue_cov_read_addr]; // @[Coverage map for ShiftQueue]
  assign ShiftQueue_cov_write_data = 1'h1;
  assign ShiftQueue_cov_write_addr = ShiftQueue_state;
  assign ShiftQueue_cov_write_mask = 1'h1;
  assign ShiftQueue_cov_write_en = 1'h1;
  assign valid_1_shl = valid_1;
  assign valid_1_pad = valid_1_shl;
  assign valid_0_shl = valid_0;
  assign valid_0_pad = valid_0_shl;
  assign valid_2_shl = valid_2;
  assign valid_2_pad = valid_2_shl;
  assign valid_4_shl = valid_4;
  assign valid_4_pad = valid_4_shl;
  assign valid_3_shl = valid_3;
  assign valid_3_pad = valid_3_shl;
  assign ShiftQueue_xor1 = valid_1_pad ^ valid_0_pad;
  assign ShiftQueue_xor6 = valid_4_pad ^ valid_3_pad;
  assign ShiftQueue_xor2 = valid_2_pad ^ ShiftQueue_xor6;
  assign ShiftQueue_xor0 = ShiftQueue_xor1 ^ ShiftQueue_xor2;
  assign io_covSum = ShiftQueue_covSum;
  assign metaAssert = 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  valid_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  valid_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  valid_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  valid_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  valid_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  elts_0_btb_taken = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  elts_0_btb_bridx = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  elts_0_btb_entry = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  elts_0_btb_bht_history = _RAND_8[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {2{`RANDOM}};
  elts_0_pc = _RAND_9[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  elts_0_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  elts_0_xcpt_pf_inst = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  elts_0_xcpt_ae_inst = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  elts_0_replay = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  elts_1_btb_taken = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  elts_1_btb_bridx = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  elts_1_btb_entry = _RAND_16[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  elts_1_btb_bht_history = _RAND_17[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {2{`RANDOM}};
  elts_1_pc = _RAND_18[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  elts_1_data = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  elts_1_xcpt_pf_inst = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  elts_1_xcpt_ae_inst = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  elts_1_replay = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  elts_2_btb_taken = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  elts_2_btb_bridx = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  elts_2_btb_entry = _RAND_25[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  elts_2_btb_bht_history = _RAND_26[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {2{`RANDOM}};
  elts_2_pc = _RAND_27[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  elts_2_data = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  elts_2_xcpt_pf_inst = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  elts_2_xcpt_ae_inst = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  elts_2_replay = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  elts_3_btb_taken = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  elts_3_btb_bridx = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  elts_3_btb_entry = _RAND_34[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  elts_3_btb_bht_history = _RAND_35[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {2{`RANDOM}};
  elts_3_pc = _RAND_36[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  elts_3_data = _RAND_37[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  elts_3_xcpt_pf_inst = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  elts_3_xcpt_ae_inst = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  elts_3_replay = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  elts_4_btb_taken = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  elts_4_btb_bridx = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  elts_4_btb_entry = _RAND_43[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  elts_4_btb_bht_history = _RAND_44[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {2{`RANDOM}};
  elts_4_pc = _RAND_45[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  elts_4_data = _RAND_46[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  elts_4_xcpt_pf_inst = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  elts_4_xcpt_ae_inst = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  elts_4_replay = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  ShiftQueue_state = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ShiftQueue_cov[initvar] = _RAND_51[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  ShiftQueue_covSum = _RAND_52[29:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      valid_0 <= 1'h0;
    end else if (reset) begin
      valid_0 <= 1'h0;
    end else if (io_deq_ready) begin
      valid_0 <= _wen_T_3;
    end else begin
      valid_0 <= _valid_0_T_6;
    end
    if (metaReset) begin
      valid_1 <= 1'h0;
    end else if (reset) begin
      valid_1 <= 1'h0;
    end else if (io_deq_ready) begin
      valid_1 <= _wen_T_11;
    end else begin
      valid_1 <= _valid_1_T_6;
    end
    if (metaReset) begin
      valid_2 <= 1'h0;
    end else if (reset) begin
      valid_2 <= 1'h0;
    end else if (io_deq_ready) begin
      valid_2 <= _wen_T_19;
    end else begin
      valid_2 <= _valid_2_T_6;
    end
    if (metaReset) begin
      valid_3 <= 1'h0;
    end else if (reset) begin
      valid_3 <= 1'h0;
    end else if (io_deq_ready) begin
      valid_3 <= _wen_T_27;
    end else begin
      valid_3 <= _valid_3_T_6;
    end
    if (metaReset) begin
      valid_4 <= 1'h0;
    end else if (reset) begin
      valid_4 <= 1'h0;
    end else if (io_deq_ready) begin
      valid_4 <= _wen_T_34;
    end else begin
      valid_4 <= _valid_4_T_6;
    end
    if (metaReset) begin
      elts_0_btb_taken <= 1'h0;
    end else if (wen) begin
      if (valid_1) begin
        elts_0_btb_taken <= elts_1_btb_taken;
      end else begin
        elts_0_btb_taken <= io_enq_bits_btb_taken;
      end
    end
    if (metaReset) begin
      elts_0_btb_bridx <= 1'h0;
    end else if (wen) begin
      if (valid_1) begin
        elts_0_btb_bridx <= elts_1_btb_bridx;
      end else begin
        elts_0_btb_bridx <= io_enq_bits_btb_bridx;
      end
    end
    if (metaReset) begin
      elts_0_btb_entry <= 5'h0;
    end else if (wen) begin
      if (valid_1) begin
        elts_0_btb_entry <= elts_1_btb_entry;
      end else begin
        elts_0_btb_entry <= io_enq_bits_btb_entry;
      end
    end
    if (metaReset) begin
      elts_0_btb_bht_history <= 8'h0;
    end else if (wen) begin
      if (valid_1) begin
        elts_0_btb_bht_history <= elts_1_btb_bht_history;
      end else begin
        elts_0_btb_bht_history <= io_enq_bits_btb_bht_history;
      end
    end
    if (metaReset) begin
      elts_0_pc <= 40'h0;
    end else if (wen) begin
      if (valid_1) begin
        elts_0_pc <= elts_1_pc;
      end else begin
        elts_0_pc <= io_enq_bits_pc;
      end
    end
    if (metaReset) begin
      elts_0_data <= 32'h0;
    end else if (wen) begin
      if (valid_1) begin
        elts_0_data <= elts_1_data;
      end else begin
        elts_0_data <= io_enq_bits_data;
      end
    end
    if (metaReset) begin
      elts_0_xcpt_pf_inst <= 1'h0;
    end else if (wen) begin
      if (valid_1) begin
        elts_0_xcpt_pf_inst <= elts_1_xcpt_pf_inst;
      end else begin
        elts_0_xcpt_pf_inst <= io_enq_bits_xcpt_pf_inst;
      end
    end
    if (metaReset) begin
      elts_0_xcpt_ae_inst <= 1'h0;
    end else if (wen) begin
      if (valid_1) begin
        elts_0_xcpt_ae_inst <= elts_1_xcpt_ae_inst;
      end else begin
        elts_0_xcpt_ae_inst <= io_enq_bits_xcpt_ae_inst;
      end
    end
    if (metaReset) begin
      elts_0_replay <= 1'h0;
    end else if (wen) begin
      if (valid_1) begin
        elts_0_replay <= elts_1_replay;
      end else begin
        elts_0_replay <= io_enq_bits_replay;
      end
    end
    if (metaReset) begin
      elts_1_btb_taken <= 1'h0;
    end else if (wen_1) begin
      if (valid_2) begin
        elts_1_btb_taken <= elts_2_btb_taken;
      end else begin
        elts_1_btb_taken <= io_enq_bits_btb_taken;
      end
    end
    if (metaReset) begin
      elts_1_btb_bridx <= 1'h0;
    end else if (wen_1) begin
      if (valid_2) begin
        elts_1_btb_bridx <= elts_2_btb_bridx;
      end else begin
        elts_1_btb_bridx <= io_enq_bits_btb_bridx;
      end
    end
    if (metaReset) begin
      elts_1_btb_entry <= 5'h0;
    end else if (wen_1) begin
      if (valid_2) begin
        elts_1_btb_entry <= elts_2_btb_entry;
      end else begin
        elts_1_btb_entry <= io_enq_bits_btb_entry;
      end
    end
    if (metaReset) begin
      elts_1_btb_bht_history <= 8'h0;
    end else if (wen_1) begin
      if (valid_2) begin
        elts_1_btb_bht_history <= elts_2_btb_bht_history;
      end else begin
        elts_1_btb_bht_history <= io_enq_bits_btb_bht_history;
      end
    end
    if (metaReset) begin
      elts_1_pc <= 40'h0;
    end else if (wen_1) begin
      if (valid_2) begin
        elts_1_pc <= elts_2_pc;
      end else begin
        elts_1_pc <= io_enq_bits_pc;
      end
    end
    if (metaReset) begin
      elts_1_data <= 32'h0;
    end else if (wen_1) begin
      if (valid_2) begin
        elts_1_data <= elts_2_data;
      end else begin
        elts_1_data <= io_enq_bits_data;
      end
    end
    if (metaReset) begin
      elts_1_xcpt_pf_inst <= 1'h0;
    end else if (wen_1) begin
      if (valid_2) begin
        elts_1_xcpt_pf_inst <= elts_2_xcpt_pf_inst;
      end else begin
        elts_1_xcpt_pf_inst <= io_enq_bits_xcpt_pf_inst;
      end
    end
    if (metaReset) begin
      elts_1_xcpt_ae_inst <= 1'h0;
    end else if (wen_1) begin
      if (valid_2) begin
        elts_1_xcpt_ae_inst <= elts_2_xcpt_ae_inst;
      end else begin
        elts_1_xcpt_ae_inst <= io_enq_bits_xcpt_ae_inst;
      end
    end
    if (metaReset) begin
      elts_1_replay <= 1'h0;
    end else if (wen_1) begin
      if (valid_2) begin
        elts_1_replay <= elts_2_replay;
      end else begin
        elts_1_replay <= io_enq_bits_replay;
      end
    end
    if (metaReset) begin
      elts_2_btb_taken <= 1'h0;
    end else if (wen_2) begin
      if (valid_3) begin
        elts_2_btb_taken <= elts_3_btb_taken;
      end else begin
        elts_2_btb_taken <= io_enq_bits_btb_taken;
      end
    end
    if (metaReset) begin
      elts_2_btb_bridx <= 1'h0;
    end else if (wen_2) begin
      if (valid_3) begin
        elts_2_btb_bridx <= elts_3_btb_bridx;
      end else begin
        elts_2_btb_bridx <= io_enq_bits_btb_bridx;
      end
    end
    if (metaReset) begin
      elts_2_btb_entry <= 5'h0;
    end else if (wen_2) begin
      if (valid_3) begin
        elts_2_btb_entry <= elts_3_btb_entry;
      end else begin
        elts_2_btb_entry <= io_enq_bits_btb_entry;
      end
    end
    if (metaReset) begin
      elts_2_btb_bht_history <= 8'h0;
    end else if (wen_2) begin
      if (valid_3) begin
        elts_2_btb_bht_history <= elts_3_btb_bht_history;
      end else begin
        elts_2_btb_bht_history <= io_enq_bits_btb_bht_history;
      end
    end
    if (metaReset) begin
      elts_2_pc <= 40'h0;
    end else if (wen_2) begin
      if (valid_3) begin
        elts_2_pc <= elts_3_pc;
      end else begin
        elts_2_pc <= io_enq_bits_pc;
      end
    end
    if (metaReset) begin
      elts_2_data <= 32'h0;
    end else if (wen_2) begin
      if (valid_3) begin
        elts_2_data <= elts_3_data;
      end else begin
        elts_2_data <= io_enq_bits_data;
      end
    end
    if (metaReset) begin
      elts_2_xcpt_pf_inst <= 1'h0;
    end else if (wen_2) begin
      if (valid_3) begin
        elts_2_xcpt_pf_inst <= elts_3_xcpt_pf_inst;
      end else begin
        elts_2_xcpt_pf_inst <= io_enq_bits_xcpt_pf_inst;
      end
    end
    if (metaReset) begin
      elts_2_xcpt_ae_inst <= 1'h0;
    end else if (wen_2) begin
      if (valid_3) begin
        elts_2_xcpt_ae_inst <= elts_3_xcpt_ae_inst;
      end else begin
        elts_2_xcpt_ae_inst <= io_enq_bits_xcpt_ae_inst;
      end
    end
    if (metaReset) begin
      elts_2_replay <= 1'h0;
    end else if (wen_2) begin
      if (valid_3) begin
        elts_2_replay <= elts_3_replay;
      end else begin
        elts_2_replay <= io_enq_bits_replay;
      end
    end
    if (metaReset) begin
      elts_3_btb_taken <= 1'h0;
    end else if (wen_3) begin
      if (valid_4) begin
        elts_3_btb_taken <= elts_4_btb_taken;
      end else begin
        elts_3_btb_taken <= io_enq_bits_btb_taken;
      end
    end
    if (metaReset) begin
      elts_3_btb_bridx <= 1'h0;
    end else if (wen_3) begin
      if (valid_4) begin
        elts_3_btb_bridx <= elts_4_btb_bridx;
      end else begin
        elts_3_btb_bridx <= io_enq_bits_btb_bridx;
      end
    end
    if (metaReset) begin
      elts_3_btb_entry <= 5'h0;
    end else if (wen_3) begin
      if (valid_4) begin
        elts_3_btb_entry <= elts_4_btb_entry;
      end else begin
        elts_3_btb_entry <= io_enq_bits_btb_entry;
      end
    end
    if (metaReset) begin
      elts_3_btb_bht_history <= 8'h0;
    end else if (wen_3) begin
      if (valid_4) begin
        elts_3_btb_bht_history <= elts_4_btb_bht_history;
      end else begin
        elts_3_btb_bht_history <= io_enq_bits_btb_bht_history;
      end
    end
    if (metaReset) begin
      elts_3_pc <= 40'h0;
    end else if (wen_3) begin
      if (valid_4) begin
        elts_3_pc <= elts_4_pc;
      end else begin
        elts_3_pc <= io_enq_bits_pc;
      end
    end
    if (metaReset) begin
      elts_3_data <= 32'h0;
    end else if (wen_3) begin
      if (valid_4) begin
        elts_3_data <= elts_4_data;
      end else begin
        elts_3_data <= io_enq_bits_data;
      end
    end
    if (metaReset) begin
      elts_3_xcpt_pf_inst <= 1'h0;
    end else if (wen_3) begin
      if (valid_4) begin
        elts_3_xcpt_pf_inst <= elts_4_xcpt_pf_inst;
      end else begin
        elts_3_xcpt_pf_inst <= io_enq_bits_xcpt_pf_inst;
      end
    end
    if (metaReset) begin
      elts_3_xcpt_ae_inst <= 1'h0;
    end else if (wen_3) begin
      if (valid_4) begin
        elts_3_xcpt_ae_inst <= elts_4_xcpt_ae_inst;
      end else begin
        elts_3_xcpt_ae_inst <= io_enq_bits_xcpt_ae_inst;
      end
    end
    if (metaReset) begin
      elts_3_replay <= 1'h0;
    end else if (wen_3) begin
      if (valid_4) begin
        elts_3_replay <= elts_4_replay;
      end else begin
        elts_3_replay <= io_enq_bits_replay;
      end
    end
    if (metaReset) begin
      elts_4_btb_taken <= 1'h0;
    end else if (wen_4) begin
      elts_4_btb_taken <= io_enq_bits_btb_taken;
    end
    if (metaReset) begin
      elts_4_btb_bridx <= 1'h0;
    end else if (wen_4) begin
      elts_4_btb_bridx <= io_enq_bits_btb_bridx;
    end
    if (metaReset) begin
      elts_4_btb_entry <= 5'h0;
    end else if (wen_4) begin
      elts_4_btb_entry <= io_enq_bits_btb_entry;
    end
    if (metaReset) begin
      elts_4_btb_bht_history <= 8'h0;
    end else if (wen_4) begin
      elts_4_btb_bht_history <= io_enq_bits_btb_bht_history;
    end
    if (metaReset) begin
      elts_4_pc <= 40'h0;
    end else if (wen_4) begin
      elts_4_pc <= io_enq_bits_pc;
    end
    if (metaReset) begin
      elts_4_data <= 32'h0;
    end else if (wen_4) begin
      elts_4_data <= io_enq_bits_data;
    end
    if (metaReset) begin
      elts_4_xcpt_pf_inst <= 1'h0;
    end else if (wen_4) begin
      elts_4_xcpt_pf_inst <= io_enq_bits_xcpt_pf_inst;
    end
    if (metaReset) begin
      elts_4_xcpt_ae_inst <= 1'h0;
    end else if (wen_4) begin
      elts_4_xcpt_ae_inst <= io_enq_bits_xcpt_ae_inst;
    end
    if (metaReset) begin
      elts_4_replay <= 1'h0;
    end else if (wen_4) begin
      elts_4_replay <= io_enq_bits_replay;
    end
    ShiftQueue_state <= ShiftQueue_xor0;
    if (!(ShiftQueue_cov_read_data)) begin
      ShiftQueue_covSum <= ShiftQueue_covSum + 1'h1;
    end
  end
  always @(posedge clock) begin
    if(ShiftQueue_cov_write_en & ShiftQueue_cov_write_mask) begin
      ShiftQueue_cov[ShiftQueue_cov_write_addr] <= ShiftQueue_cov_write_data; // @[Coverage map for ShiftQueue]
    end
  end
endmodule
module TLB_1(
  input         clock,
  input         reset,
  output        io_req_ready,
  input         io_req_valid,
  input  [39:0] io_req_bits_vaddr,
  output        io_resp_miss,
  output [31:0] io_resp_paddr,
  output        io_resp_pf_inst,
  output        io_resp_ae_inst,
  output        io_resp_cacheable,
  input         io_sfence_valid,
  input         io_sfence_bits_rs1,
  input         io_sfence_bits_rs2,
  input  [38:0] io_sfence_bits_addr,
  input         io_ptw_req_ready,
  output        io_ptw_req_valid,
  output        io_ptw_req_bits_valid,
  output [26:0] io_ptw_req_bits_bits_addr,
  input         io_ptw_resp_valid,
  input         io_ptw_resp_bits_ae,
  input  [53:0] io_ptw_resp_bits_pte_ppn,
  input         io_ptw_resp_bits_pte_d,
  input         io_ptw_resp_bits_pte_a,
  input         io_ptw_resp_bits_pte_g,
  input         io_ptw_resp_bits_pte_u,
  input         io_ptw_resp_bits_pte_x,
  input         io_ptw_resp_bits_pte_w,
  input         io_ptw_resp_bits_pte_r,
  input         io_ptw_resp_bits_pte_v,
  input  [1:0]  io_ptw_resp_bits_level,
  input         io_ptw_resp_bits_homogeneous,
  input  [3:0]  io_ptw_ptbr_mode,
  input         io_ptw_status_debug,
  input  [1:0]  io_ptw_status_prv,
  input         io_ptw_pmp_0_cfg_l,
  input  [1:0]  io_ptw_pmp_0_cfg_a,
  input         io_ptw_pmp_0_cfg_x,
  input         io_ptw_pmp_0_cfg_w,
  input         io_ptw_pmp_0_cfg_r,
  input  [29:0] io_ptw_pmp_0_addr,
  input  [31:0] io_ptw_pmp_0_mask,
  input         io_ptw_pmp_1_cfg_l,
  input  [1:0]  io_ptw_pmp_1_cfg_a,
  input         io_ptw_pmp_1_cfg_x,
  input         io_ptw_pmp_1_cfg_w,
  input         io_ptw_pmp_1_cfg_r,
  input  [29:0] io_ptw_pmp_1_addr,
  input  [31:0] io_ptw_pmp_1_mask,
  input         io_ptw_pmp_2_cfg_l,
  input  [1:0]  io_ptw_pmp_2_cfg_a,
  input         io_ptw_pmp_2_cfg_x,
  input         io_ptw_pmp_2_cfg_w,
  input         io_ptw_pmp_2_cfg_r,
  input  [29:0] io_ptw_pmp_2_addr,
  input  [31:0] io_ptw_pmp_2_mask,
  input         io_ptw_pmp_3_cfg_l,
  input  [1:0]  io_ptw_pmp_3_cfg_a,
  input         io_ptw_pmp_3_cfg_x,
  input         io_ptw_pmp_3_cfg_w,
  input         io_ptw_pmp_3_cfg_r,
  input  [29:0] io_ptw_pmp_3_addr,
  input  [31:0] io_ptw_pmp_3_mask,
  input         io_ptw_pmp_4_cfg_l,
  input  [1:0]  io_ptw_pmp_4_cfg_a,
  input         io_ptw_pmp_4_cfg_x,
  input         io_ptw_pmp_4_cfg_w,
  input         io_ptw_pmp_4_cfg_r,
  input  [29:0] io_ptw_pmp_4_addr,
  input  [31:0] io_ptw_pmp_4_mask,
  input         io_ptw_pmp_5_cfg_l,
  input  [1:0]  io_ptw_pmp_5_cfg_a,
  input         io_ptw_pmp_5_cfg_x,
  input         io_ptw_pmp_5_cfg_w,
  input         io_ptw_pmp_5_cfg_r,
  input  [29:0] io_ptw_pmp_5_addr,
  input  [31:0] io_ptw_pmp_5_mask,
  input         io_ptw_pmp_6_cfg_l,
  input  [1:0]  io_ptw_pmp_6_cfg_a,
  input         io_ptw_pmp_6_cfg_x,
  input         io_ptw_pmp_6_cfg_w,
  input         io_ptw_pmp_6_cfg_r,
  input  [29:0] io_ptw_pmp_6_addr,
  input  [31:0] io_ptw_pmp_6_mask,
  input         io_ptw_pmp_7_cfg_l,
  input  [1:0]  io_ptw_pmp_7_cfg_a,
  input         io_ptw_pmp_7_cfg_x,
  input         io_ptw_pmp_7_cfg_w,
  input         io_ptw_pmp_7_cfg_r,
  input  [29:0] io_ptw_pmp_7_addr,
  input  [31:0] io_ptw_pmp_7_mask,
  input         io_kill,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  wire [19:0] mpu_ppn_barrier_io_x_ppn; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_x_u; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_x_ae; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_x_sw; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_x_sx; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_x_sr; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_x_pw; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_x_px; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_x_pr; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_x_ppp; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_x_pal; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_x_paa; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_x_eff; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_x_c; // @[package.scala 258:25]
  wire [19:0] mpu_ppn_barrier_io_y_ppn; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_y_u; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_y_ae; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_y_sw; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_y_sx; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_y_sr; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_y_pw; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_y_px; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_y_pr; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_y_ppp; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_y_pal; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_y_paa; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_y_eff; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_io_y_c; // @[package.scala 258:25]
  wire [29:0] mpu_ppn_barrier_io_covSum; // @[package.scala 258:25]
  wire  mpu_ppn_barrier_metaAssert; // @[package.scala 258:25]
  wire [1:0] pmp_io_prv; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_0_cfg_l; // @[TLB.scala 192:19]
  wire [1:0] pmp_io_pmp_0_cfg_a; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_0_cfg_x; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_0_cfg_w; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_0_cfg_r; // @[TLB.scala 192:19]
  wire [29:0] pmp_io_pmp_0_addr; // @[TLB.scala 192:19]
  wire [31:0] pmp_io_pmp_0_mask; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_1_cfg_l; // @[TLB.scala 192:19]
  wire [1:0] pmp_io_pmp_1_cfg_a; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_1_cfg_x; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_1_cfg_w; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_1_cfg_r; // @[TLB.scala 192:19]
  wire [29:0] pmp_io_pmp_1_addr; // @[TLB.scala 192:19]
  wire [31:0] pmp_io_pmp_1_mask; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_2_cfg_l; // @[TLB.scala 192:19]
  wire [1:0] pmp_io_pmp_2_cfg_a; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_2_cfg_x; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_2_cfg_w; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_2_cfg_r; // @[TLB.scala 192:19]
  wire [29:0] pmp_io_pmp_2_addr; // @[TLB.scala 192:19]
  wire [31:0] pmp_io_pmp_2_mask; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_3_cfg_l; // @[TLB.scala 192:19]
  wire [1:0] pmp_io_pmp_3_cfg_a; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_3_cfg_x; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_3_cfg_w; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_3_cfg_r; // @[TLB.scala 192:19]
  wire [29:0] pmp_io_pmp_3_addr; // @[TLB.scala 192:19]
  wire [31:0] pmp_io_pmp_3_mask; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_4_cfg_l; // @[TLB.scala 192:19]
  wire [1:0] pmp_io_pmp_4_cfg_a; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_4_cfg_x; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_4_cfg_w; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_4_cfg_r; // @[TLB.scala 192:19]
  wire [29:0] pmp_io_pmp_4_addr; // @[TLB.scala 192:19]
  wire [31:0] pmp_io_pmp_4_mask; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_5_cfg_l; // @[TLB.scala 192:19]
  wire [1:0] pmp_io_pmp_5_cfg_a; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_5_cfg_x; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_5_cfg_w; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_5_cfg_r; // @[TLB.scala 192:19]
  wire [29:0] pmp_io_pmp_5_addr; // @[TLB.scala 192:19]
  wire [31:0] pmp_io_pmp_5_mask; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_6_cfg_l; // @[TLB.scala 192:19]
  wire [1:0] pmp_io_pmp_6_cfg_a; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_6_cfg_x; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_6_cfg_w; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_6_cfg_r; // @[TLB.scala 192:19]
  wire [29:0] pmp_io_pmp_6_addr; // @[TLB.scala 192:19]
  wire [31:0] pmp_io_pmp_6_mask; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_7_cfg_l; // @[TLB.scala 192:19]
  wire [1:0] pmp_io_pmp_7_cfg_a; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_7_cfg_x; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_7_cfg_w; // @[TLB.scala 192:19]
  wire  pmp_io_pmp_7_cfg_r; // @[TLB.scala 192:19]
  wire [29:0] pmp_io_pmp_7_addr; // @[TLB.scala 192:19]
  wire [31:0] pmp_io_pmp_7_mask; // @[TLB.scala 192:19]
  wire [31:0] pmp_io_addr; // @[TLB.scala 192:19]
  wire  pmp_io_r; // @[TLB.scala 192:19]
  wire  pmp_io_w; // @[TLB.scala 192:19]
  wire  pmp_io_x; // @[TLB.scala 192:19]
  wire [29:0] pmp_io_covSum; // @[TLB.scala 192:19]
  wire  pmp_metaAssert; // @[TLB.scala 192:19]
  wire [19:0] entries_barrier_io_x_ppn; // @[package.scala 258:25]
  wire  entries_barrier_io_x_u; // @[package.scala 258:25]
  wire  entries_barrier_io_x_ae; // @[package.scala 258:25]
  wire  entries_barrier_io_x_sw; // @[package.scala 258:25]
  wire  entries_barrier_io_x_sx; // @[package.scala 258:25]
  wire  entries_barrier_io_x_sr; // @[package.scala 258:25]
  wire  entries_barrier_io_x_pw; // @[package.scala 258:25]
  wire  entries_barrier_io_x_px; // @[package.scala 258:25]
  wire  entries_barrier_io_x_pr; // @[package.scala 258:25]
  wire  entries_barrier_io_x_ppp; // @[package.scala 258:25]
  wire  entries_barrier_io_x_pal; // @[package.scala 258:25]
  wire  entries_barrier_io_x_paa; // @[package.scala 258:25]
  wire  entries_barrier_io_x_eff; // @[package.scala 258:25]
  wire  entries_barrier_io_x_c; // @[package.scala 258:25]
  wire [19:0] entries_barrier_io_y_ppn; // @[package.scala 258:25]
  wire  entries_barrier_io_y_u; // @[package.scala 258:25]
  wire  entries_barrier_io_y_ae; // @[package.scala 258:25]
  wire  entries_barrier_io_y_sw; // @[package.scala 258:25]
  wire  entries_barrier_io_y_sx; // @[package.scala 258:25]
  wire  entries_barrier_io_y_sr; // @[package.scala 258:25]
  wire  entries_barrier_io_y_pw; // @[package.scala 258:25]
  wire  entries_barrier_io_y_px; // @[package.scala 258:25]
  wire  entries_barrier_io_y_pr; // @[package.scala 258:25]
  wire  entries_barrier_io_y_ppp; // @[package.scala 258:25]
  wire  entries_barrier_io_y_pal; // @[package.scala 258:25]
  wire  entries_barrier_io_y_paa; // @[package.scala 258:25]
  wire  entries_barrier_io_y_eff; // @[package.scala 258:25]
  wire  entries_barrier_io_y_c; // @[package.scala 258:25]
  wire [29:0] entries_barrier_io_covSum; // @[package.scala 258:25]
  wire  entries_barrier_metaAssert; // @[package.scala 258:25]
  wire [19:0] entries_barrier_1_io_x_ppn; // @[package.scala 258:25]
  wire  entries_barrier_1_io_x_u; // @[package.scala 258:25]
  wire  entries_barrier_1_io_x_ae; // @[package.scala 258:25]
  wire  entries_barrier_1_io_x_sw; // @[package.scala 258:25]
  wire  entries_barrier_1_io_x_sx; // @[package.scala 258:25]
  wire  entries_barrier_1_io_x_sr; // @[package.scala 258:25]
  wire  entries_barrier_1_io_x_pw; // @[package.scala 258:25]
  wire  entries_barrier_1_io_x_px; // @[package.scala 258:25]
  wire  entries_barrier_1_io_x_pr; // @[package.scala 258:25]
  wire  entries_barrier_1_io_x_ppp; // @[package.scala 258:25]
  wire  entries_barrier_1_io_x_pal; // @[package.scala 258:25]
  wire  entries_barrier_1_io_x_paa; // @[package.scala 258:25]
  wire  entries_barrier_1_io_x_eff; // @[package.scala 258:25]
  wire  entries_barrier_1_io_x_c; // @[package.scala 258:25]
  wire [19:0] entries_barrier_1_io_y_ppn; // @[package.scala 258:25]
  wire  entries_barrier_1_io_y_u; // @[package.scala 258:25]
  wire  entries_barrier_1_io_y_ae; // @[package.scala 258:25]
  wire  entries_barrier_1_io_y_sw; // @[package.scala 258:25]
  wire  entries_barrier_1_io_y_sx; // @[package.scala 258:25]
  wire  entries_barrier_1_io_y_sr; // @[package.scala 258:25]
  wire  entries_barrier_1_io_y_pw; // @[package.scala 258:25]
  wire  entries_barrier_1_io_y_px; // @[package.scala 258:25]
  wire  entries_barrier_1_io_y_pr; // @[package.scala 258:25]
  wire  entries_barrier_1_io_y_ppp; // @[package.scala 258:25]
  wire  entries_barrier_1_io_y_pal; // @[package.scala 258:25]
  wire  entries_barrier_1_io_y_paa; // @[package.scala 258:25]
  wire  entries_barrier_1_io_y_eff; // @[package.scala 258:25]
  wire  entries_barrier_1_io_y_c; // @[package.scala 258:25]
  wire [29:0] entries_barrier_1_io_covSum; // @[package.scala 258:25]
  wire  entries_barrier_1_metaAssert; // @[package.scala 258:25]
  wire [19:0] entries_barrier_2_io_x_ppn; // @[package.scala 258:25]
  wire  entries_barrier_2_io_x_u; // @[package.scala 258:25]
  wire  entries_barrier_2_io_x_ae; // @[package.scala 258:25]
  wire  entries_barrier_2_io_x_sw; // @[package.scala 258:25]
  wire  entries_barrier_2_io_x_sx; // @[package.scala 258:25]
  wire  entries_barrier_2_io_x_sr; // @[package.scala 258:25]
  wire  entries_barrier_2_io_x_pw; // @[package.scala 258:25]
  wire  entries_barrier_2_io_x_px; // @[package.scala 258:25]
  wire  entries_barrier_2_io_x_pr; // @[package.scala 258:25]
  wire  entries_barrier_2_io_x_ppp; // @[package.scala 258:25]
  wire  entries_barrier_2_io_x_pal; // @[package.scala 258:25]
  wire  entries_barrier_2_io_x_paa; // @[package.scala 258:25]
  wire  entries_barrier_2_io_x_eff; // @[package.scala 258:25]
  wire  entries_barrier_2_io_x_c; // @[package.scala 258:25]
  wire [19:0] entries_barrier_2_io_y_ppn; // @[package.scala 258:25]
  wire  entries_barrier_2_io_y_u; // @[package.scala 258:25]
  wire  entries_barrier_2_io_y_ae; // @[package.scala 258:25]
  wire  entries_barrier_2_io_y_sw; // @[package.scala 258:25]
  wire  entries_barrier_2_io_y_sx; // @[package.scala 258:25]
  wire  entries_barrier_2_io_y_sr; // @[package.scala 258:25]
  wire  entries_barrier_2_io_y_pw; // @[package.scala 258:25]
  wire  entries_barrier_2_io_y_px; // @[package.scala 258:25]
  wire  entries_barrier_2_io_y_pr; // @[package.scala 258:25]
  wire  entries_barrier_2_io_y_ppp; // @[package.scala 258:25]
  wire  entries_barrier_2_io_y_pal; // @[package.scala 258:25]
  wire  entries_barrier_2_io_y_paa; // @[package.scala 258:25]
  wire  entries_barrier_2_io_y_eff; // @[package.scala 258:25]
  wire  entries_barrier_2_io_y_c; // @[package.scala 258:25]
  wire [29:0] entries_barrier_2_io_covSum; // @[package.scala 258:25]
  wire  entries_barrier_2_metaAssert; // @[package.scala 258:25]
  wire [19:0] entries_barrier_3_io_x_ppn; // @[package.scala 258:25]
  wire  entries_barrier_3_io_x_u; // @[package.scala 258:25]
  wire  entries_barrier_3_io_x_ae; // @[package.scala 258:25]
  wire  entries_barrier_3_io_x_sw; // @[package.scala 258:25]
  wire  entries_barrier_3_io_x_sx; // @[package.scala 258:25]
  wire  entries_barrier_3_io_x_sr; // @[package.scala 258:25]
  wire  entries_barrier_3_io_x_pw; // @[package.scala 258:25]
  wire  entries_barrier_3_io_x_px; // @[package.scala 258:25]
  wire  entries_barrier_3_io_x_pr; // @[package.scala 258:25]
  wire  entries_barrier_3_io_x_ppp; // @[package.scala 258:25]
  wire  entries_barrier_3_io_x_pal; // @[package.scala 258:25]
  wire  entries_barrier_3_io_x_paa; // @[package.scala 258:25]
  wire  entries_barrier_3_io_x_eff; // @[package.scala 258:25]
  wire  entries_barrier_3_io_x_c; // @[package.scala 258:25]
  wire [19:0] entries_barrier_3_io_y_ppn; // @[package.scala 258:25]
  wire  entries_barrier_3_io_y_u; // @[package.scala 258:25]
  wire  entries_barrier_3_io_y_ae; // @[package.scala 258:25]
  wire  entries_barrier_3_io_y_sw; // @[package.scala 258:25]
  wire  entries_barrier_3_io_y_sx; // @[package.scala 258:25]
  wire  entries_barrier_3_io_y_sr; // @[package.scala 258:25]
  wire  entries_barrier_3_io_y_pw; // @[package.scala 258:25]
  wire  entries_barrier_3_io_y_px; // @[package.scala 258:25]
  wire  entries_barrier_3_io_y_pr; // @[package.scala 258:25]
  wire  entries_barrier_3_io_y_ppp; // @[package.scala 258:25]
  wire  entries_barrier_3_io_y_pal; // @[package.scala 258:25]
  wire  entries_barrier_3_io_y_paa; // @[package.scala 258:25]
  wire  entries_barrier_3_io_y_eff; // @[package.scala 258:25]
  wire  entries_barrier_3_io_y_c; // @[package.scala 258:25]
  wire [29:0] entries_barrier_3_io_covSum; // @[package.scala 258:25]
  wire  entries_barrier_3_metaAssert; // @[package.scala 258:25]
  wire [19:0] entries_barrier_4_io_x_ppn; // @[package.scala 258:25]
  wire  entries_barrier_4_io_x_u; // @[package.scala 258:25]
  wire  entries_barrier_4_io_x_ae; // @[package.scala 258:25]
  wire  entries_barrier_4_io_x_sw; // @[package.scala 258:25]
  wire  entries_barrier_4_io_x_sx; // @[package.scala 258:25]
  wire  entries_barrier_4_io_x_sr; // @[package.scala 258:25]
  wire  entries_barrier_4_io_x_pw; // @[package.scala 258:25]
  wire  entries_barrier_4_io_x_px; // @[package.scala 258:25]
  wire  entries_barrier_4_io_x_pr; // @[package.scala 258:25]
  wire  entries_barrier_4_io_x_ppp; // @[package.scala 258:25]
  wire  entries_barrier_4_io_x_pal; // @[package.scala 258:25]
  wire  entries_barrier_4_io_x_paa; // @[package.scala 258:25]
  wire  entries_barrier_4_io_x_eff; // @[package.scala 258:25]
  wire  entries_barrier_4_io_x_c; // @[package.scala 258:25]
  wire [19:0] entries_barrier_4_io_y_ppn; // @[package.scala 258:25]
  wire  entries_barrier_4_io_y_u; // @[package.scala 258:25]
  wire  entries_barrier_4_io_y_ae; // @[package.scala 258:25]
  wire  entries_barrier_4_io_y_sw; // @[package.scala 258:25]
  wire  entries_barrier_4_io_y_sx; // @[package.scala 258:25]
  wire  entries_barrier_4_io_y_sr; // @[package.scala 258:25]
  wire  entries_barrier_4_io_y_pw; // @[package.scala 258:25]
  wire  entries_barrier_4_io_y_px; // @[package.scala 258:25]
  wire  entries_barrier_4_io_y_pr; // @[package.scala 258:25]
  wire  entries_barrier_4_io_y_ppp; // @[package.scala 258:25]
  wire  entries_barrier_4_io_y_pal; // @[package.scala 258:25]
  wire  entries_barrier_4_io_y_paa; // @[package.scala 258:25]
  wire  entries_barrier_4_io_y_eff; // @[package.scala 258:25]
  wire  entries_barrier_4_io_y_c; // @[package.scala 258:25]
  wire [29:0] entries_barrier_4_io_covSum; // @[package.scala 258:25]
  wire  entries_barrier_4_metaAssert; // @[package.scala 258:25]
  wire [19:0] entries_barrier_5_io_x_ppn; // @[package.scala 258:25]
  wire  entries_barrier_5_io_x_u; // @[package.scala 258:25]
  wire  entries_barrier_5_io_x_ae; // @[package.scala 258:25]
  wire  entries_barrier_5_io_x_sw; // @[package.scala 258:25]
  wire  entries_barrier_5_io_x_sx; // @[package.scala 258:25]
  wire  entries_barrier_5_io_x_sr; // @[package.scala 258:25]
  wire  entries_barrier_5_io_x_pw; // @[package.scala 258:25]
  wire  entries_barrier_5_io_x_px; // @[package.scala 258:25]
  wire  entries_barrier_5_io_x_pr; // @[package.scala 258:25]
  wire  entries_barrier_5_io_x_ppp; // @[package.scala 258:25]
  wire  entries_barrier_5_io_x_pal; // @[package.scala 258:25]
  wire  entries_barrier_5_io_x_paa; // @[package.scala 258:25]
  wire  entries_barrier_5_io_x_eff; // @[package.scala 258:25]
  wire  entries_barrier_5_io_x_c; // @[package.scala 258:25]
  wire [19:0] entries_barrier_5_io_y_ppn; // @[package.scala 258:25]
  wire  entries_barrier_5_io_y_u; // @[package.scala 258:25]
  wire  entries_barrier_5_io_y_ae; // @[package.scala 258:25]
  wire  entries_barrier_5_io_y_sw; // @[package.scala 258:25]
  wire  entries_barrier_5_io_y_sx; // @[package.scala 258:25]
  wire  entries_barrier_5_io_y_sr; // @[package.scala 258:25]
  wire  entries_barrier_5_io_y_pw; // @[package.scala 258:25]
  wire  entries_barrier_5_io_y_px; // @[package.scala 258:25]
  wire  entries_barrier_5_io_y_pr; // @[package.scala 258:25]
  wire  entries_barrier_5_io_y_ppp; // @[package.scala 258:25]
  wire  entries_barrier_5_io_y_pal; // @[package.scala 258:25]
  wire  entries_barrier_5_io_y_paa; // @[package.scala 258:25]
  wire  entries_barrier_5_io_y_eff; // @[package.scala 258:25]
  wire  entries_barrier_5_io_y_c; // @[package.scala 258:25]
  wire [29:0] entries_barrier_5_io_covSum; // @[package.scala 258:25]
  wire  entries_barrier_5_metaAssert; // @[package.scala 258:25]
  wire [19:0] entries_barrier_6_io_x_ppn; // @[package.scala 258:25]
  wire  entries_barrier_6_io_x_u; // @[package.scala 258:25]
  wire  entries_barrier_6_io_x_ae; // @[package.scala 258:25]
  wire  entries_barrier_6_io_x_sw; // @[package.scala 258:25]
  wire  entries_barrier_6_io_x_sx; // @[package.scala 258:25]
  wire  entries_barrier_6_io_x_sr; // @[package.scala 258:25]
  wire  entries_barrier_6_io_x_pw; // @[package.scala 258:25]
  wire  entries_barrier_6_io_x_px; // @[package.scala 258:25]
  wire  entries_barrier_6_io_x_pr; // @[package.scala 258:25]
  wire  entries_barrier_6_io_x_ppp; // @[package.scala 258:25]
  wire  entries_barrier_6_io_x_pal; // @[package.scala 258:25]
  wire  entries_barrier_6_io_x_paa; // @[package.scala 258:25]
  wire  entries_barrier_6_io_x_eff; // @[package.scala 258:25]
  wire  entries_barrier_6_io_x_c; // @[package.scala 258:25]
  wire [19:0] entries_barrier_6_io_y_ppn; // @[package.scala 258:25]
  wire  entries_barrier_6_io_y_u; // @[package.scala 258:25]
  wire  entries_barrier_6_io_y_ae; // @[package.scala 258:25]
  wire  entries_barrier_6_io_y_sw; // @[package.scala 258:25]
  wire  entries_barrier_6_io_y_sx; // @[package.scala 258:25]
  wire  entries_barrier_6_io_y_sr; // @[package.scala 258:25]
  wire  entries_barrier_6_io_y_pw; // @[package.scala 258:25]
  wire  entries_barrier_6_io_y_px; // @[package.scala 258:25]
  wire  entries_barrier_6_io_y_pr; // @[package.scala 258:25]
  wire  entries_barrier_6_io_y_ppp; // @[package.scala 258:25]
  wire  entries_barrier_6_io_y_pal; // @[package.scala 258:25]
  wire  entries_barrier_6_io_y_paa; // @[package.scala 258:25]
  wire  entries_barrier_6_io_y_eff; // @[package.scala 258:25]
  wire  entries_barrier_6_io_y_c; // @[package.scala 258:25]
  wire [29:0] entries_barrier_6_io_covSum; // @[package.scala 258:25]
  wire  entries_barrier_6_metaAssert; // @[package.scala 258:25]
  wire [19:0] entries_barrier_7_io_x_ppn; // @[package.scala 258:25]
  wire  entries_barrier_7_io_x_u; // @[package.scala 258:25]
  wire  entries_barrier_7_io_x_ae; // @[package.scala 258:25]
  wire  entries_barrier_7_io_x_sw; // @[package.scala 258:25]
  wire  entries_barrier_7_io_x_sx; // @[package.scala 258:25]
  wire  entries_barrier_7_io_x_sr; // @[package.scala 258:25]
  wire  entries_barrier_7_io_x_pw; // @[package.scala 258:25]
  wire  entries_barrier_7_io_x_px; // @[package.scala 258:25]
  wire  entries_barrier_7_io_x_pr; // @[package.scala 258:25]
  wire  entries_barrier_7_io_x_ppp; // @[package.scala 258:25]
  wire  entries_barrier_7_io_x_pal; // @[package.scala 258:25]
  wire  entries_barrier_7_io_x_paa; // @[package.scala 258:25]
  wire  entries_barrier_7_io_x_eff; // @[package.scala 258:25]
  wire  entries_barrier_7_io_x_c; // @[package.scala 258:25]
  wire [19:0] entries_barrier_7_io_y_ppn; // @[package.scala 258:25]
  wire  entries_barrier_7_io_y_u; // @[package.scala 258:25]
  wire  entries_barrier_7_io_y_ae; // @[package.scala 258:25]
  wire  entries_barrier_7_io_y_sw; // @[package.scala 258:25]
  wire  entries_barrier_7_io_y_sx; // @[package.scala 258:25]
  wire  entries_barrier_7_io_y_sr; // @[package.scala 258:25]
  wire  entries_barrier_7_io_y_pw; // @[package.scala 258:25]
  wire  entries_barrier_7_io_y_px; // @[package.scala 258:25]
  wire  entries_barrier_7_io_y_pr; // @[package.scala 258:25]
  wire  entries_barrier_7_io_y_ppp; // @[package.scala 258:25]
  wire  entries_barrier_7_io_y_pal; // @[package.scala 258:25]
  wire  entries_barrier_7_io_y_paa; // @[package.scala 258:25]
  wire  entries_barrier_7_io_y_eff; // @[package.scala 258:25]
  wire  entries_barrier_7_io_y_c; // @[package.scala 258:25]
  wire [29:0] entries_barrier_7_io_covSum; // @[package.scala 258:25]
  wire  entries_barrier_7_metaAssert; // @[package.scala 258:25]
  wire [19:0] entries_barrier_8_io_x_ppn; // @[package.scala 258:25]
  wire  entries_barrier_8_io_x_u; // @[package.scala 258:25]
  wire  entries_barrier_8_io_x_ae; // @[package.scala 258:25]
  wire  entries_barrier_8_io_x_sw; // @[package.scala 258:25]
  wire  entries_barrier_8_io_x_sx; // @[package.scala 258:25]
  wire  entries_barrier_8_io_x_sr; // @[package.scala 258:25]
  wire  entries_barrier_8_io_x_pw; // @[package.scala 258:25]
  wire  entries_barrier_8_io_x_px; // @[package.scala 258:25]
  wire  entries_barrier_8_io_x_pr; // @[package.scala 258:25]
  wire  entries_barrier_8_io_x_ppp; // @[package.scala 258:25]
  wire  entries_barrier_8_io_x_pal; // @[package.scala 258:25]
  wire  entries_barrier_8_io_x_paa; // @[package.scala 258:25]
  wire  entries_barrier_8_io_x_eff; // @[package.scala 258:25]
  wire  entries_barrier_8_io_x_c; // @[package.scala 258:25]
  wire [19:0] entries_barrier_8_io_y_ppn; // @[package.scala 258:25]
  wire  entries_barrier_8_io_y_u; // @[package.scala 258:25]
  wire  entries_barrier_8_io_y_ae; // @[package.scala 258:25]
  wire  entries_barrier_8_io_y_sw; // @[package.scala 258:25]
  wire  entries_barrier_8_io_y_sx; // @[package.scala 258:25]
  wire  entries_barrier_8_io_y_sr; // @[package.scala 258:25]
  wire  entries_barrier_8_io_y_pw; // @[package.scala 258:25]
  wire  entries_barrier_8_io_y_px; // @[package.scala 258:25]
  wire  entries_barrier_8_io_y_pr; // @[package.scala 258:25]
  wire  entries_barrier_8_io_y_ppp; // @[package.scala 258:25]
  wire  entries_barrier_8_io_y_pal; // @[package.scala 258:25]
  wire  entries_barrier_8_io_y_paa; // @[package.scala 258:25]
  wire  entries_barrier_8_io_y_eff; // @[package.scala 258:25]
  wire  entries_barrier_8_io_y_c; // @[package.scala 258:25]
  wire [29:0] entries_barrier_8_io_covSum; // @[package.scala 258:25]
  wire  entries_barrier_8_metaAssert; // @[package.scala 258:25]
  wire [19:0] entries_barrier_9_io_x_ppn; // @[package.scala 258:25]
  wire  entries_barrier_9_io_x_u; // @[package.scala 258:25]
  wire  entries_barrier_9_io_x_ae; // @[package.scala 258:25]
  wire  entries_barrier_9_io_x_sw; // @[package.scala 258:25]
  wire  entries_barrier_9_io_x_sx; // @[package.scala 258:25]
  wire  entries_barrier_9_io_x_sr; // @[package.scala 258:25]
  wire  entries_barrier_9_io_x_pw; // @[package.scala 258:25]
  wire  entries_barrier_9_io_x_px; // @[package.scala 258:25]
  wire  entries_barrier_9_io_x_pr; // @[package.scala 258:25]
  wire  entries_barrier_9_io_x_ppp; // @[package.scala 258:25]
  wire  entries_barrier_9_io_x_pal; // @[package.scala 258:25]
  wire  entries_barrier_9_io_x_paa; // @[package.scala 258:25]
  wire  entries_barrier_9_io_x_eff; // @[package.scala 258:25]
  wire  entries_barrier_9_io_x_c; // @[package.scala 258:25]
  wire [19:0] entries_barrier_9_io_y_ppn; // @[package.scala 258:25]
  wire  entries_barrier_9_io_y_u; // @[package.scala 258:25]
  wire  entries_barrier_9_io_y_ae; // @[package.scala 258:25]
  wire  entries_barrier_9_io_y_sw; // @[package.scala 258:25]
  wire  entries_barrier_9_io_y_sx; // @[package.scala 258:25]
  wire  entries_barrier_9_io_y_sr; // @[package.scala 258:25]
  wire  entries_barrier_9_io_y_pw; // @[package.scala 258:25]
  wire  entries_barrier_9_io_y_px; // @[package.scala 258:25]
  wire  entries_barrier_9_io_y_pr; // @[package.scala 258:25]
  wire  entries_barrier_9_io_y_ppp; // @[package.scala 258:25]
  wire  entries_barrier_9_io_y_pal; // @[package.scala 258:25]
  wire  entries_barrier_9_io_y_paa; // @[package.scala 258:25]
  wire  entries_barrier_9_io_y_eff; // @[package.scala 258:25]
  wire  entries_barrier_9_io_y_c; // @[package.scala 258:25]
  wire [29:0] entries_barrier_9_io_covSum; // @[package.scala 258:25]
  wire  entries_barrier_9_metaAssert; // @[package.scala 258:25]
  wire [19:0] entries_barrier_10_io_x_ppn; // @[package.scala 258:25]
  wire  entries_barrier_10_io_x_u; // @[package.scala 258:25]
  wire  entries_barrier_10_io_x_ae; // @[package.scala 258:25]
  wire  entries_barrier_10_io_x_sw; // @[package.scala 258:25]
  wire  entries_barrier_10_io_x_sx; // @[package.scala 258:25]
  wire  entries_barrier_10_io_x_sr; // @[package.scala 258:25]
  wire  entries_barrier_10_io_x_pw; // @[package.scala 258:25]
  wire  entries_barrier_10_io_x_px; // @[package.scala 258:25]
  wire  entries_barrier_10_io_x_pr; // @[package.scala 258:25]
  wire  entries_barrier_10_io_x_ppp; // @[package.scala 258:25]
  wire  entries_barrier_10_io_x_pal; // @[package.scala 258:25]
  wire  entries_barrier_10_io_x_paa; // @[package.scala 258:25]
  wire  entries_barrier_10_io_x_eff; // @[package.scala 258:25]
  wire  entries_barrier_10_io_x_c; // @[package.scala 258:25]
  wire [19:0] entries_barrier_10_io_y_ppn; // @[package.scala 258:25]
  wire  entries_barrier_10_io_y_u; // @[package.scala 258:25]
  wire  entries_barrier_10_io_y_ae; // @[package.scala 258:25]
  wire  entries_barrier_10_io_y_sw; // @[package.scala 258:25]
  wire  entries_barrier_10_io_y_sx; // @[package.scala 258:25]
  wire  entries_barrier_10_io_y_sr; // @[package.scala 258:25]
  wire  entries_barrier_10_io_y_pw; // @[package.scala 258:25]
  wire  entries_barrier_10_io_y_px; // @[package.scala 258:25]
  wire  entries_barrier_10_io_y_pr; // @[package.scala 258:25]
  wire  entries_barrier_10_io_y_ppp; // @[package.scala 258:25]
  wire  entries_barrier_10_io_y_pal; // @[package.scala 258:25]
  wire  entries_barrier_10_io_y_paa; // @[package.scala 258:25]
  wire  entries_barrier_10_io_y_eff; // @[package.scala 258:25]
  wire  entries_barrier_10_io_y_c; // @[package.scala 258:25]
  wire [29:0] entries_barrier_10_io_covSum; // @[package.scala 258:25]
  wire  entries_barrier_10_metaAssert; // @[package.scala 258:25]
  wire [19:0] entries_barrier_11_io_x_ppn; // @[package.scala 258:25]
  wire  entries_barrier_11_io_x_u; // @[package.scala 258:25]
  wire  entries_barrier_11_io_x_ae; // @[package.scala 258:25]
  wire  entries_barrier_11_io_x_sw; // @[package.scala 258:25]
  wire  entries_barrier_11_io_x_sx; // @[package.scala 258:25]
  wire  entries_barrier_11_io_x_sr; // @[package.scala 258:25]
  wire  entries_barrier_11_io_x_pw; // @[package.scala 258:25]
  wire  entries_barrier_11_io_x_px; // @[package.scala 258:25]
  wire  entries_barrier_11_io_x_pr; // @[package.scala 258:25]
  wire  entries_barrier_11_io_x_ppp; // @[package.scala 258:25]
  wire  entries_barrier_11_io_x_pal; // @[package.scala 258:25]
  wire  entries_barrier_11_io_x_paa; // @[package.scala 258:25]
  wire  entries_barrier_11_io_x_eff; // @[package.scala 258:25]
  wire  entries_barrier_11_io_x_c; // @[package.scala 258:25]
  wire [19:0] entries_barrier_11_io_y_ppn; // @[package.scala 258:25]
  wire  entries_barrier_11_io_y_u; // @[package.scala 258:25]
  wire  entries_barrier_11_io_y_ae; // @[package.scala 258:25]
  wire  entries_barrier_11_io_y_sw; // @[package.scala 258:25]
  wire  entries_barrier_11_io_y_sx; // @[package.scala 258:25]
  wire  entries_barrier_11_io_y_sr; // @[package.scala 258:25]
  wire  entries_barrier_11_io_y_pw; // @[package.scala 258:25]
  wire  entries_barrier_11_io_y_px; // @[package.scala 258:25]
  wire  entries_barrier_11_io_y_pr; // @[package.scala 258:25]
  wire  entries_barrier_11_io_y_ppp; // @[package.scala 258:25]
  wire  entries_barrier_11_io_y_pal; // @[package.scala 258:25]
  wire  entries_barrier_11_io_y_paa; // @[package.scala 258:25]
  wire  entries_barrier_11_io_y_eff; // @[package.scala 258:25]
  wire  entries_barrier_11_io_y_c; // @[package.scala 258:25]
  wire [29:0] entries_barrier_11_io_covSum; // @[package.scala 258:25]
  wire  entries_barrier_11_metaAssert; // @[package.scala 258:25]
  wire [19:0] entries_barrier_12_io_x_ppn; // @[package.scala 258:25]
  wire  entries_barrier_12_io_x_u; // @[package.scala 258:25]
  wire  entries_barrier_12_io_x_ae; // @[package.scala 258:25]
  wire  entries_barrier_12_io_x_sw; // @[package.scala 258:25]
  wire  entries_barrier_12_io_x_sx; // @[package.scala 258:25]
  wire  entries_barrier_12_io_x_sr; // @[package.scala 258:25]
  wire  entries_barrier_12_io_x_pw; // @[package.scala 258:25]
  wire  entries_barrier_12_io_x_px; // @[package.scala 258:25]
  wire  entries_barrier_12_io_x_pr; // @[package.scala 258:25]
  wire  entries_barrier_12_io_x_ppp; // @[package.scala 258:25]
  wire  entries_barrier_12_io_x_pal; // @[package.scala 258:25]
  wire  entries_barrier_12_io_x_paa; // @[package.scala 258:25]
  wire  entries_barrier_12_io_x_eff; // @[package.scala 258:25]
  wire  entries_barrier_12_io_x_c; // @[package.scala 258:25]
  wire [19:0] entries_barrier_12_io_y_ppn; // @[package.scala 258:25]
  wire  entries_barrier_12_io_y_u; // @[package.scala 258:25]
  wire  entries_barrier_12_io_y_ae; // @[package.scala 258:25]
  wire  entries_barrier_12_io_y_sw; // @[package.scala 258:25]
  wire  entries_barrier_12_io_y_sx; // @[package.scala 258:25]
  wire  entries_barrier_12_io_y_sr; // @[package.scala 258:25]
  wire  entries_barrier_12_io_y_pw; // @[package.scala 258:25]
  wire  entries_barrier_12_io_y_px; // @[package.scala 258:25]
  wire  entries_barrier_12_io_y_pr; // @[package.scala 258:25]
  wire  entries_barrier_12_io_y_ppp; // @[package.scala 258:25]
  wire  entries_barrier_12_io_y_pal; // @[package.scala 258:25]
  wire  entries_barrier_12_io_y_paa; // @[package.scala 258:25]
  wire  entries_barrier_12_io_y_eff; // @[package.scala 258:25]
  wire  entries_barrier_12_io_y_c; // @[package.scala 258:25]
  wire [29:0] entries_barrier_12_io_covSum; // @[package.scala 258:25]
  wire  entries_barrier_12_metaAssert; // @[package.scala 258:25]
  wire [26:0] vpn; // @[TLB.scala 162:30]
  reg [26:0] sectored_entries_0_0_tag; // @[TLB.scala 164:29]
  reg [31:0] _RAND_0;
  reg [34:0] sectored_entries_0_0_data_0; // @[TLB.scala 164:29]
  reg [63:0] _RAND_1;
  reg [34:0] sectored_entries_0_0_data_1; // @[TLB.scala 164:29]
  reg [63:0] _RAND_2;
  reg [34:0] sectored_entries_0_0_data_2; // @[TLB.scala 164:29]
  reg [63:0] _RAND_3;
  reg [34:0] sectored_entries_0_0_data_3; // @[TLB.scala 164:29]
  reg [63:0] _RAND_4;
  reg  sectored_entries_0_0_valid_0; // @[TLB.scala 164:29]
  reg [31:0] _RAND_5;
  reg  sectored_entries_0_0_valid_1; // @[TLB.scala 164:29]
  reg [31:0] _RAND_6;
  reg  sectored_entries_0_0_valid_2; // @[TLB.scala 164:29]
  reg [31:0] _RAND_7;
  reg  sectored_entries_0_0_valid_3; // @[TLB.scala 164:29]
  reg [31:0] _RAND_8;
  reg [26:0] sectored_entries_0_1_tag; // @[TLB.scala 164:29]
  reg [31:0] _RAND_9;
  reg [34:0] sectored_entries_0_1_data_0; // @[TLB.scala 164:29]
  reg [63:0] _RAND_10;
  reg [34:0] sectored_entries_0_1_data_1; // @[TLB.scala 164:29]
  reg [63:0] _RAND_11;
  reg [34:0] sectored_entries_0_1_data_2; // @[TLB.scala 164:29]
  reg [63:0] _RAND_12;
  reg [34:0] sectored_entries_0_1_data_3; // @[TLB.scala 164:29]
  reg [63:0] _RAND_13;
  reg  sectored_entries_0_1_valid_0; // @[TLB.scala 164:29]
  reg [31:0] _RAND_14;
  reg  sectored_entries_0_1_valid_1; // @[TLB.scala 164:29]
  reg [31:0] _RAND_15;
  reg  sectored_entries_0_1_valid_2; // @[TLB.scala 164:29]
  reg [31:0] _RAND_16;
  reg  sectored_entries_0_1_valid_3; // @[TLB.scala 164:29]
  reg [31:0] _RAND_17;
  reg [26:0] sectored_entries_0_2_tag; // @[TLB.scala 164:29]
  reg [31:0] _RAND_18;
  reg [34:0] sectored_entries_0_2_data_0; // @[TLB.scala 164:29]
  reg [63:0] _RAND_19;
  reg [34:0] sectored_entries_0_2_data_1; // @[TLB.scala 164:29]
  reg [63:0] _RAND_20;
  reg [34:0] sectored_entries_0_2_data_2; // @[TLB.scala 164:29]
  reg [63:0] _RAND_21;
  reg [34:0] sectored_entries_0_2_data_3; // @[TLB.scala 164:29]
  reg [63:0] _RAND_22;
  reg  sectored_entries_0_2_valid_0; // @[TLB.scala 164:29]
  reg [31:0] _RAND_23;
  reg  sectored_entries_0_2_valid_1; // @[TLB.scala 164:29]
  reg [31:0] _RAND_24;
  reg  sectored_entries_0_2_valid_2; // @[TLB.scala 164:29]
  reg [31:0] _RAND_25;
  reg  sectored_entries_0_2_valid_3; // @[TLB.scala 164:29]
  reg [31:0] _RAND_26;
  reg [26:0] sectored_entries_0_3_tag; // @[TLB.scala 164:29]
  reg [31:0] _RAND_27;
  reg [34:0] sectored_entries_0_3_data_0; // @[TLB.scala 164:29]
  reg [63:0] _RAND_28;
  reg [34:0] sectored_entries_0_3_data_1; // @[TLB.scala 164:29]
  reg [63:0] _RAND_29;
  reg [34:0] sectored_entries_0_3_data_2; // @[TLB.scala 164:29]
  reg [63:0] _RAND_30;
  reg [34:0] sectored_entries_0_3_data_3; // @[TLB.scala 164:29]
  reg [63:0] _RAND_31;
  reg  sectored_entries_0_3_valid_0; // @[TLB.scala 164:29]
  reg [31:0] _RAND_32;
  reg  sectored_entries_0_3_valid_1; // @[TLB.scala 164:29]
  reg [31:0] _RAND_33;
  reg  sectored_entries_0_3_valid_2; // @[TLB.scala 164:29]
  reg [31:0] _RAND_34;
  reg  sectored_entries_0_3_valid_3; // @[TLB.scala 164:29]
  reg [31:0] _RAND_35;
  reg [26:0] sectored_entries_0_4_tag; // @[TLB.scala 164:29]
  reg [31:0] _RAND_36;
  reg [34:0] sectored_entries_0_4_data_0; // @[TLB.scala 164:29]
  reg [63:0] _RAND_37;
  reg [34:0] sectored_entries_0_4_data_1; // @[TLB.scala 164:29]
  reg [63:0] _RAND_38;
  reg [34:0] sectored_entries_0_4_data_2; // @[TLB.scala 164:29]
  reg [63:0] _RAND_39;
  reg [34:0] sectored_entries_0_4_data_3; // @[TLB.scala 164:29]
  reg [63:0] _RAND_40;
  reg  sectored_entries_0_4_valid_0; // @[TLB.scala 164:29]
  reg [31:0] _RAND_41;
  reg  sectored_entries_0_4_valid_1; // @[TLB.scala 164:29]
  reg [31:0] _RAND_42;
  reg  sectored_entries_0_4_valid_2; // @[TLB.scala 164:29]
  reg [31:0] _RAND_43;
  reg  sectored_entries_0_4_valid_3; // @[TLB.scala 164:29]
  reg [31:0] _RAND_44;
  reg [26:0] sectored_entries_0_5_tag; // @[TLB.scala 164:29]
  reg [31:0] _RAND_45;
  reg [34:0] sectored_entries_0_5_data_0; // @[TLB.scala 164:29]
  reg [63:0] _RAND_46;
  reg [34:0] sectored_entries_0_5_data_1; // @[TLB.scala 164:29]
  reg [63:0] _RAND_47;
  reg [34:0] sectored_entries_0_5_data_2; // @[TLB.scala 164:29]
  reg [63:0] _RAND_48;
  reg [34:0] sectored_entries_0_5_data_3; // @[TLB.scala 164:29]
  reg [63:0] _RAND_49;
  reg  sectored_entries_0_5_valid_0; // @[TLB.scala 164:29]
  reg [31:0] _RAND_50;
  reg  sectored_entries_0_5_valid_1; // @[TLB.scala 164:29]
  reg [31:0] _RAND_51;
  reg  sectored_entries_0_5_valid_2; // @[TLB.scala 164:29]
  reg [31:0] _RAND_52;
  reg  sectored_entries_0_5_valid_3; // @[TLB.scala 164:29]
  reg [31:0] _RAND_53;
  reg [26:0] sectored_entries_0_6_tag; // @[TLB.scala 164:29]
  reg [31:0] _RAND_54;
  reg [34:0] sectored_entries_0_6_data_0; // @[TLB.scala 164:29]
  reg [63:0] _RAND_55;
  reg [34:0] sectored_entries_0_6_data_1; // @[TLB.scala 164:29]
  reg [63:0] _RAND_56;
  reg [34:0] sectored_entries_0_6_data_2; // @[TLB.scala 164:29]
  reg [63:0] _RAND_57;
  reg [34:0] sectored_entries_0_6_data_3; // @[TLB.scala 164:29]
  reg [63:0] _RAND_58;
  reg  sectored_entries_0_6_valid_0; // @[TLB.scala 164:29]
  reg [31:0] _RAND_59;
  reg  sectored_entries_0_6_valid_1; // @[TLB.scala 164:29]
  reg [31:0] _RAND_60;
  reg  sectored_entries_0_6_valid_2; // @[TLB.scala 164:29]
  reg [31:0] _RAND_61;
  reg  sectored_entries_0_6_valid_3; // @[TLB.scala 164:29]
  reg [31:0] _RAND_62;
  reg [26:0] sectored_entries_0_7_tag; // @[TLB.scala 164:29]
  reg [31:0] _RAND_63;
  reg [34:0] sectored_entries_0_7_data_0; // @[TLB.scala 164:29]
  reg [63:0] _RAND_64;
  reg [34:0] sectored_entries_0_7_data_1; // @[TLB.scala 164:29]
  reg [63:0] _RAND_65;
  reg [34:0] sectored_entries_0_7_data_2; // @[TLB.scala 164:29]
  reg [63:0] _RAND_66;
  reg [34:0] sectored_entries_0_7_data_3; // @[TLB.scala 164:29]
  reg [63:0] _RAND_67;
  reg  sectored_entries_0_7_valid_0; // @[TLB.scala 164:29]
  reg [31:0] _RAND_68;
  reg  sectored_entries_0_7_valid_1; // @[TLB.scala 164:29]
  reg [31:0] _RAND_69;
  reg  sectored_entries_0_7_valid_2; // @[TLB.scala 164:29]
  reg [31:0] _RAND_70;
  reg  sectored_entries_0_7_valid_3; // @[TLB.scala 164:29]
  reg [31:0] _RAND_71;
  reg [1:0] superpage_entries_0_level; // @[TLB.scala 165:30]
  reg [31:0] _RAND_72;
  reg [26:0] superpage_entries_0_tag; // @[TLB.scala 165:30]
  reg [31:0] _RAND_73;
  reg [34:0] superpage_entries_0_data_0; // @[TLB.scala 165:30]
  reg [63:0] _RAND_74;
  reg  superpage_entries_0_valid_0; // @[TLB.scala 165:30]
  reg [31:0] _RAND_75;
  reg [1:0] superpage_entries_1_level; // @[TLB.scala 165:30]
  reg [31:0] _RAND_76;
  reg [26:0] superpage_entries_1_tag; // @[TLB.scala 165:30]
  reg [31:0] _RAND_77;
  reg [34:0] superpage_entries_1_data_0; // @[TLB.scala 165:30]
  reg [63:0] _RAND_78;
  reg  superpage_entries_1_valid_0; // @[TLB.scala 165:30]
  reg [31:0] _RAND_79;
  reg [1:0] superpage_entries_2_level; // @[TLB.scala 165:30]
  reg [31:0] _RAND_80;
  reg [26:0] superpage_entries_2_tag; // @[TLB.scala 165:30]
  reg [31:0] _RAND_81;
  reg [34:0] superpage_entries_2_data_0; // @[TLB.scala 165:30]
  reg [63:0] _RAND_82;
  reg  superpage_entries_2_valid_0; // @[TLB.scala 165:30]
  reg [31:0] _RAND_83;
  reg [1:0] superpage_entries_3_level; // @[TLB.scala 165:30]
  reg [31:0] _RAND_84;
  reg [26:0] superpage_entries_3_tag; // @[TLB.scala 165:30]
  reg [31:0] _RAND_85;
  reg [34:0] superpage_entries_3_data_0; // @[TLB.scala 165:30]
  reg [63:0] _RAND_86;
  reg  superpage_entries_3_valid_0; // @[TLB.scala 165:30]
  reg [31:0] _RAND_87;
  reg [1:0] special_entry_level; // @[TLB.scala 166:56]
  reg [31:0] _RAND_88;
  reg [26:0] special_entry_tag; // @[TLB.scala 166:56]
  reg [31:0] _RAND_89;
  reg [34:0] special_entry_data_0; // @[TLB.scala 166:56]
  reg [63:0] _RAND_90;
  reg  special_entry_valid_0; // @[TLB.scala 166:56]
  reg [31:0] _RAND_91;
  reg [1:0] state; // @[TLB.scala 172:18]
  reg [31:0] _RAND_92;
  reg [26:0] r_refill_tag; // @[TLB.scala 173:25]
  reg [31:0] _RAND_93;
  reg [1:0] r_superpage_repl_addr; // @[TLB.scala 174:34]
  reg [31:0] _RAND_94;
  reg [2:0] r_sectored_repl_addr; // @[TLB.scala 175:33]
  reg [31:0] _RAND_95;
  reg [2:0] r_sectored_hit_addr; // @[TLB.scala 176:32]
  reg [31:0] _RAND_96;
  reg  r_sectored_hit; // @[TLB.scala 177:27]
  reg [31:0] _RAND_97;
  wire  priv_s; // @[TLB.scala 180:20]
  wire  priv_uses_vm; // @[TLB.scala 181:27]
  wire  vm_enabled; // @[TLB.scala 182:83]
  wire [19:0] refill_ppn; // @[TLB.scala 185:44]
  wire  _invalidate_refill_T; // @[package.scala 15:47]
  wire  _invalidate_refill_T_1; // @[package.scala 15:47]
  wire  _invalidate_refill_T_2; // @[package.scala 72:59]
  wire  invalidate_refill; // @[TLB.scala 187:88]
  wire [1:0] mpu_ppn_hi; // @[TLB.scala 105:26]
  wire  mpu_ppn_ignore; // @[TLB.scala 107:28]
  wire [26:0] _mpu_ppn_T_17; // @[TLB.scala 108:28]
  wire [26:0] _GEN_919; // @[TLB.scala 108:47]
  wire [26:0] _mpu_ppn_T_18; // @[TLB.scala 108:47]
  wire [8:0] mpu_ppn_lo; // @[TLB.scala 108:58]
  wire  mpu_ppn_ignore_1; // @[TLB.scala 107:28]
  wire [26:0] _mpu_ppn_T_19; // @[TLB.scala 108:28]
  wire [26:0] _mpu_ppn_T_20; // @[TLB.scala 108:47]
  wire [8:0] mpu_ppn_lo_1; // @[TLB.scala 108:58]
  wire [19:0] _mpu_ppn_T_21; // @[Cat.scala 30:58]
  wire [27:0] _mpu_ppn_T_23; // @[TLB.scala 189:20]
  wire [27:0] mpu_ppn; // @[TLB.scala 188:20]
  wire [11:0] mpu_physaddr_lo; // @[TLB.scala 190:52]
  wire [39:0] mpu_physaddr; // @[Cat.scala 30:58]
  wire [2:0] _mpu_priv_T_2; // @[Cat.scala 30:58]
  wire [2:0] mpu_priv; // @[TLB.scala 191:27]
  wire [39:0] _legal_address_T; // @[Parameters.scala 137:31]
  wire [40:0] _legal_address_T_1; // @[Parameters.scala 137:49]
  wire [40:0] _legal_address_T_3; // @[Parameters.scala 137:52]
  wire  _legal_address_T_4; // @[Parameters.scala 137:67]
  wire [39:0] _legal_address_T_5; // @[Parameters.scala 137:31]
  wire [40:0] _legal_address_T_6; // @[Parameters.scala 137:49]
  wire [40:0] _legal_address_T_8; // @[Parameters.scala 137:52]
  wire  _legal_address_T_9; // @[Parameters.scala 137:67]
  wire [39:0] _legal_address_T_10; // @[Parameters.scala 137:31]
  wire [40:0] _legal_address_T_11; // @[Parameters.scala 137:49]
  wire [40:0] _legal_address_T_13; // @[Parameters.scala 137:52]
  wire  _legal_address_T_14; // @[Parameters.scala 137:67]
  wire [40:0] _legal_address_T_16; // @[Parameters.scala 137:49]
  wire [40:0] _legal_address_T_18; // @[Parameters.scala 137:52]
  wire  _legal_address_T_19; // @[Parameters.scala 137:67]
  wire [39:0] _legal_address_T_20; // @[Parameters.scala 137:31]
  wire [40:0] _legal_address_T_21; // @[Parameters.scala 137:49]
  wire [40:0] _legal_address_T_23; // @[Parameters.scala 137:52]
  wire  _legal_address_T_24; // @[Parameters.scala 137:67]
  wire [39:0] _legal_address_T_25; // @[Parameters.scala 137:31]
  wire [40:0] _legal_address_T_26; // @[Parameters.scala 137:49]
  wire [40:0] _legal_address_T_28; // @[Parameters.scala 137:52]
  wire  _legal_address_T_29; // @[Parameters.scala 137:67]
  wire [39:0] _legal_address_T_30; // @[Parameters.scala 137:31]
  wire [40:0] _legal_address_T_31; // @[Parameters.scala 137:49]
  wire [40:0] _legal_address_T_33; // @[Parameters.scala 137:52]
  wire  _legal_address_T_34; // @[Parameters.scala 137:67]
  wire  _legal_address_T_35; // @[TLB.scala 197:67]
  wire  _legal_address_T_36; // @[TLB.scala 197:67]
  wire  _legal_address_T_37; // @[TLB.scala 197:67]
  wire  _legal_address_T_38; // @[TLB.scala 197:67]
  wire  _legal_address_T_39; // @[TLB.scala 197:67]
  wire  legal_address; // @[TLB.scala 197:67]
  wire [40:0] _cacheable_T_8; // @[Parameters.scala 137:52]
  wire  _cacheable_T_9; // @[Parameters.scala 137:67]
  wire  cacheable; // @[TLB.scala 199:19]
  wire [39:0] _homogeneous_T_54; // @[Parameters.scala 137:31]
  wire [40:0] _homogeneous_T_55; // @[Parameters.scala 137:49]
  wire [40:0] _homogeneous_T_57; // @[Parameters.scala 137:52]
  wire  _homogeneous_T_58; // @[Parameters.scala 137:67]
  wire [40:0] _homogeneous_T_71; // @[Parameters.scala 137:52]
  wire  _homogeneous_T_72; // @[Parameters.scala 137:67]
  wire  _homogeneous_T_79; // @[TLBPermissions.scala 83:66]
  wire  _deny_access_to_debug_T; // @[TLB.scala 202:39]
  wire  deny_access_to_debug; // @[TLB.scala 202:48]
  wire  _prot_r_T_7; // @[TLB.scala 203:41]
  wire  prot_r; // @[TLB.scala 203:66]
  wire [39:0] _prot_w_T_10; // @[Parameters.scala 137:31]
  wire [40:0] _prot_w_T_11; // @[Parameters.scala 137:49]
  wire [40:0] _prot_w_T_13; // @[Parameters.scala 137:52]
  wire  _prot_w_T_14; // @[Parameters.scala 137:67]
  wire [40:0] _prot_w_T_18; // @[Parameters.scala 137:52]
  wire  _prot_w_T_19; // @[Parameters.scala 137:67]
  wire  _prot_w_T_21; // @[Parameters.scala 615:89]
  wire  _prot_w_T_22; // @[Parameters.scala 615:89]
  wire  _prot_w_T_31; // @[TLB.scala 199:19]
  wire  _prot_w_T_33; // @[TLB.scala 204:45]
  wire  prot_w; // @[TLB.scala 204:70]
  wire  prot_al; // @[TLB.scala 199:19]
  wire [40:0] _prot_x_T_3; // @[Parameters.scala 137:52]
  wire  _prot_x_T_4; // @[Parameters.scala 137:67]
  wire  _prot_x_T_15; // @[Parameters.scala 615:89]
  wire  _prot_x_T_16; // @[Parameters.scala 615:89]
  wire  _prot_x_T_31; // @[TLB.scala 199:19]
  wire  _prot_x_T_33; // @[TLB.scala 208:40]
  wire  prot_x; // @[TLB.scala 208:65]
  wire [40:0] _prot_eff_T_20; // @[Parameters.scala 137:52]
  wire  _prot_eff_T_21; // @[Parameters.scala 137:67]
  wire [40:0] _prot_eff_T_25; // @[Parameters.scala 137:52]
  wire  _prot_eff_T_26; // @[Parameters.scala 137:67]
  wire  _prot_eff_T_37; // @[Parameters.scala 615:89]
  wire  _prot_eff_T_38; // @[Parameters.scala 615:89]
  wire  _prot_eff_T_39; // @[Parameters.scala 615:89]
  wire  prot_eff; // @[TLB.scala 199:19]
  wire  _sector_hits_T; // @[package.scala 72:59]
  wire  _sector_hits_T_1; // @[package.scala 72:59]
  wire  _sector_hits_T_2; // @[package.scala 72:59]
  wire [26:0] _sector_hits_T_3; // @[TLB.scala 88:41]
  wire  _sector_hits_T_5; // @[TLB.scala 88:66]
  wire  sector_hits_0; // @[TLB.scala 87:40]
  wire  _sector_hits_T_6; // @[package.scala 72:59]
  wire  _sector_hits_T_7; // @[package.scala 72:59]
  wire  _sector_hits_T_8; // @[package.scala 72:59]
  wire [26:0] _sector_hits_T_9; // @[TLB.scala 88:41]
  wire  _sector_hits_T_11; // @[TLB.scala 88:66]
  wire  sector_hits_1; // @[TLB.scala 87:40]
  wire  _sector_hits_T_12; // @[package.scala 72:59]
  wire  _sector_hits_T_13; // @[package.scala 72:59]
  wire  _sector_hits_T_14; // @[package.scala 72:59]
  wire [26:0] _sector_hits_T_15; // @[TLB.scala 88:41]
  wire  _sector_hits_T_17; // @[TLB.scala 88:66]
  wire  sector_hits_2; // @[TLB.scala 87:40]
  wire  _sector_hits_T_18; // @[package.scala 72:59]
  wire  _sector_hits_T_19; // @[package.scala 72:59]
  wire  _sector_hits_T_20; // @[package.scala 72:59]
  wire [26:0] _sector_hits_T_21; // @[TLB.scala 88:41]
  wire  _sector_hits_T_23; // @[TLB.scala 88:66]
  wire  sector_hits_3; // @[TLB.scala 87:40]
  wire  _sector_hits_T_24; // @[package.scala 72:59]
  wire  _sector_hits_T_25; // @[package.scala 72:59]
  wire  _sector_hits_T_26; // @[package.scala 72:59]
  wire [26:0] _sector_hits_T_27; // @[TLB.scala 88:41]
  wire  _sector_hits_T_29; // @[TLB.scala 88:66]
  wire  sector_hits_4; // @[TLB.scala 87:40]
  wire  _sector_hits_T_30; // @[package.scala 72:59]
  wire  _sector_hits_T_31; // @[package.scala 72:59]
  wire  _sector_hits_T_32; // @[package.scala 72:59]
  wire [26:0] _sector_hits_T_33; // @[TLB.scala 88:41]
  wire  _sector_hits_T_35; // @[TLB.scala 88:66]
  wire  sector_hits_5; // @[TLB.scala 87:40]
  wire  _sector_hits_T_36; // @[package.scala 72:59]
  wire  _sector_hits_T_37; // @[package.scala 72:59]
  wire  _sector_hits_T_38; // @[package.scala 72:59]
  wire [26:0] _sector_hits_T_39; // @[TLB.scala 88:41]
  wire  _sector_hits_T_41; // @[TLB.scala 88:66]
  wire  sector_hits_6; // @[TLB.scala 87:40]
  wire  _sector_hits_T_42; // @[package.scala 72:59]
  wire  _sector_hits_T_43; // @[package.scala 72:59]
  wire  _sector_hits_T_44; // @[package.scala 72:59]
  wire [26:0] _sector_hits_T_45; // @[TLB.scala 88:41]
  wire  _sector_hits_T_47; // @[TLB.scala 88:66]
  wire  sector_hits_7; // @[TLB.scala 87:40]
  wire  _superpage_hits_T_2; // @[TLB.scala 95:77]
  wire  _superpage_hits_T_4; // @[TLB.scala 95:29]
  wire  superpage_hits_ignore_1; // @[TLB.scala 94:28]
  wire  _superpage_hits_T_7; // @[TLB.scala 95:77]
  wire  _superpage_hits_T_8; // @[TLB.scala 95:40]
  wire  superpage_hits_0; // @[TLB.scala 95:29]
  wire  _superpage_hits_T_16; // @[TLB.scala 95:77]
  wire  _superpage_hits_T_18; // @[TLB.scala 95:29]
  wire  superpage_hits_ignore_4; // @[TLB.scala 94:28]
  wire  _superpage_hits_T_21; // @[TLB.scala 95:77]
  wire  _superpage_hits_T_22; // @[TLB.scala 95:40]
  wire  superpage_hits_1; // @[TLB.scala 95:29]
  wire  _superpage_hits_T_30; // @[TLB.scala 95:77]
  wire  _superpage_hits_T_32; // @[TLB.scala 95:29]
  wire  superpage_hits_ignore_7; // @[TLB.scala 94:28]
  wire  _superpage_hits_T_35; // @[TLB.scala 95:77]
  wire  _superpage_hits_T_36; // @[TLB.scala 95:40]
  wire  superpage_hits_2; // @[TLB.scala 95:29]
  wire  _superpage_hits_T_44; // @[TLB.scala 95:77]
  wire  _superpage_hits_T_46; // @[TLB.scala 95:29]
  wire  superpage_hits_ignore_10; // @[TLB.scala 94:28]
  wire  _superpage_hits_T_49; // @[TLB.scala 95:77]
  wire  _superpage_hits_T_50; // @[TLB.scala 95:40]
  wire  superpage_hits_3; // @[TLB.scala 95:29]
  wire [1:0] hitsVec_idx; // @[package.scala 154:13]
  wire  _GEN_1; // @[TLB.scala 100:18]
  wire  _GEN_2; // @[TLB.scala 100:18]
  wire  _GEN_3; // @[TLB.scala 100:18]
  wire  _hitsVec_T_3; // @[TLB.scala 100:18]
  wire  hitsVec_0; // @[TLB.scala 213:44]
  wire  _GEN_5; // @[TLB.scala 100:18]
  wire  _GEN_6; // @[TLB.scala 100:18]
  wire  _GEN_7; // @[TLB.scala 100:18]
  wire  _hitsVec_T_7; // @[TLB.scala 100:18]
  wire  hitsVec_1; // @[TLB.scala 213:44]
  wire  _GEN_9; // @[TLB.scala 100:18]
  wire  _GEN_10; // @[TLB.scala 100:18]
  wire  _GEN_11; // @[TLB.scala 100:18]
  wire  _hitsVec_T_11; // @[TLB.scala 100:18]
  wire  hitsVec_2; // @[TLB.scala 213:44]
  wire  _GEN_13; // @[TLB.scala 100:18]
  wire  _GEN_14; // @[TLB.scala 100:18]
  wire  _GEN_15; // @[TLB.scala 100:18]
  wire  _hitsVec_T_15; // @[TLB.scala 100:18]
  wire  hitsVec_3; // @[TLB.scala 213:44]
  wire  _GEN_17; // @[TLB.scala 100:18]
  wire  _GEN_18; // @[TLB.scala 100:18]
  wire  _GEN_19; // @[TLB.scala 100:18]
  wire  _hitsVec_T_19; // @[TLB.scala 100:18]
  wire  hitsVec_4; // @[TLB.scala 213:44]
  wire  _GEN_21; // @[TLB.scala 100:18]
  wire  _GEN_22; // @[TLB.scala 100:18]
  wire  _GEN_23; // @[TLB.scala 100:18]
  wire  _hitsVec_T_23; // @[TLB.scala 100:18]
  wire  hitsVec_5; // @[TLB.scala 213:44]
  wire  _GEN_25; // @[TLB.scala 100:18]
  wire  _GEN_26; // @[TLB.scala 100:18]
  wire  _GEN_27; // @[TLB.scala 100:18]
  wire  _hitsVec_T_27; // @[TLB.scala 100:18]
  wire  hitsVec_6; // @[TLB.scala 213:44]
  wire  _GEN_29; // @[TLB.scala 100:18]
  wire  _GEN_30; // @[TLB.scala 100:18]
  wire  _GEN_31; // @[TLB.scala 100:18]
  wire  _hitsVec_T_31; // @[TLB.scala 100:18]
  wire  hitsVec_7; // @[TLB.scala 213:44]
  wire  hitsVec_8; // @[TLB.scala 213:44]
  wire  hitsVec_9; // @[TLB.scala 213:44]
  wire  hitsVec_10; // @[TLB.scala 213:44]
  wire  hitsVec_11; // @[TLB.scala 213:44]
  wire  _hitsVec_T_94; // @[TLB.scala 95:77]
  wire  _hitsVec_T_96; // @[TLB.scala 95:29]
  wire  _hitsVec_T_99; // @[TLB.scala 95:77]
  wire  _hitsVec_T_100; // @[TLB.scala 95:40]
  wire  _hitsVec_T_101; // @[TLB.scala 95:29]
  wire  _hitsVec_T_104; // @[TLB.scala 95:77]
  wire  _hitsVec_T_105; // @[TLB.scala 95:40]
  wire  _hitsVec_T_106; // @[TLB.scala 95:29]
  wire  hitsVec_12; // @[TLB.scala 213:44]
  wire [5:0] real_hits_lo; // @[Cat.scala 30:58]
  wire [12:0] real_hits; // @[Cat.scala 30:58]
  wire  hits_hi; // @[TLB.scala 215:18]
  wire [13:0] hits; // @[Cat.scala 30:58]
  wire  newEntry_g; // @[TLB.scala 224:25]
  wire  _newEntry_sr_T_1; // @[PTW.scala 73:44]
  wire  _newEntry_sr_T_2; // @[PTW.scala 73:38]
  wire  _newEntry_sr_T_3; // @[PTW.scala 73:32]
  wire  _newEntry_sr_T_4; // @[PTW.scala 73:52]
  wire  newEntry_sr; // @[PTW.scala 77:35]
  wire  _newEntry_sw_T_5; // @[PTW.scala 78:35]
  wire  newEntry_sw; // @[PTW.scala 78:40]
  wire  newEntry_sx; // @[PTW.scala 79:35]
  wire [7:0] special_entry_data_0_lo; // @[TLB.scala 122:24]
  wire [34:0] _special_entry_data_0_T; // @[TLB.scala 122:24]
  wire  _GEN_32; // @[TLB.scala 241:34]
  wire  _T_2; // @[TLB.scala 243:40]
  wire  _T_3; // @[TLB.scala 244:82]
  wire  _GEN_35; // @[TLB.scala 244:89]
  wire  _T_4; // @[TLB.scala 244:82]
  wire  _GEN_39; // @[TLB.scala 244:89]
  wire  _T_5; // @[TLB.scala 244:82]
  wire  _GEN_43; // @[TLB.scala 244:89]
  wire  _T_6; // @[TLB.scala 244:82]
  wire  _GEN_47; // @[TLB.scala 244:89]
  wire [2:0] waddr; // @[TLB.scala 250:22]
  wire  _T_7; // @[TLB.scala 251:75]
  wire  _GEN_49; // @[TLB.scala 252:32]
  wire  _GEN_50; // @[TLB.scala 252:32]
  wire  _GEN_51; // @[TLB.scala 252:32]
  wire  _GEN_52; // @[TLB.scala 252:32]
  wire [1:0] idx; // @[package.scala 154:13]
  wire  _GEN_921; // @[TLB.scala 121:16]
  wire  _GEN_53; // @[TLB.scala 121:16]
  wire  _GEN_922; // @[TLB.scala 121:16]
  wire  _GEN_54; // @[TLB.scala 121:16]
  wire  _GEN_923; // @[TLB.scala 121:16]
  wire  _GEN_55; // @[TLB.scala 121:16]
  wire  _GEN_924; // @[TLB.scala 121:16]
  wire  _GEN_56; // @[TLB.scala 121:16]
  wire  _GEN_61; // @[TLB.scala 254:34]
  wire  _GEN_62; // @[TLB.scala 254:34]
  wire  _GEN_63; // @[TLB.scala 254:34]
  wire  _GEN_64; // @[TLB.scala 254:34]
  wire  _GEN_65; // @[TLB.scala 251:82]
  wire  _GEN_66; // @[TLB.scala 251:82]
  wire  _GEN_67; // @[TLB.scala 251:82]
  wire  _GEN_68; // @[TLB.scala 251:82]
  wire  _T_9; // @[TLB.scala 251:75]
  wire  _GEN_75; // @[TLB.scala 252:32]
  wire  _GEN_76; // @[TLB.scala 252:32]
  wire  _GEN_77; // @[TLB.scala 252:32]
  wire  _GEN_78; // @[TLB.scala 252:32]
  wire  _GEN_79; // @[TLB.scala 121:16]
  wire  _GEN_80; // @[TLB.scala 121:16]
  wire  _GEN_81; // @[TLB.scala 121:16]
  wire  _GEN_82; // @[TLB.scala 121:16]
  wire  _GEN_87; // @[TLB.scala 254:34]
  wire  _GEN_88; // @[TLB.scala 254:34]
  wire  _GEN_89; // @[TLB.scala 254:34]
  wire  _GEN_90; // @[TLB.scala 254:34]
  wire  _GEN_91; // @[TLB.scala 251:82]
  wire  _GEN_92; // @[TLB.scala 251:82]
  wire  _GEN_93; // @[TLB.scala 251:82]
  wire  _GEN_94; // @[TLB.scala 251:82]
  wire  _T_11; // @[TLB.scala 251:75]
  wire  _GEN_101; // @[TLB.scala 252:32]
  wire  _GEN_102; // @[TLB.scala 252:32]
  wire  _GEN_103; // @[TLB.scala 252:32]
  wire  _GEN_104; // @[TLB.scala 252:32]
  wire  _GEN_105; // @[TLB.scala 121:16]
  wire  _GEN_106; // @[TLB.scala 121:16]
  wire  _GEN_107; // @[TLB.scala 121:16]
  wire  _GEN_108; // @[TLB.scala 121:16]
  wire  _GEN_113; // @[TLB.scala 254:34]
  wire  _GEN_114; // @[TLB.scala 254:34]
  wire  _GEN_115; // @[TLB.scala 254:34]
  wire  _GEN_116; // @[TLB.scala 254:34]
  wire  _GEN_117; // @[TLB.scala 251:82]
  wire  _GEN_118; // @[TLB.scala 251:82]
  wire  _GEN_119; // @[TLB.scala 251:82]
  wire  _GEN_120; // @[TLB.scala 251:82]
  wire  _T_13; // @[TLB.scala 251:75]
  wire  _GEN_127; // @[TLB.scala 252:32]
  wire  _GEN_128; // @[TLB.scala 252:32]
  wire  _GEN_129; // @[TLB.scala 252:32]
  wire  _GEN_130; // @[TLB.scala 252:32]
  wire  _GEN_131; // @[TLB.scala 121:16]
  wire  _GEN_132; // @[TLB.scala 121:16]
  wire  _GEN_133; // @[TLB.scala 121:16]
  wire  _GEN_134; // @[TLB.scala 121:16]
  wire  _GEN_139; // @[TLB.scala 254:34]
  wire  _GEN_140; // @[TLB.scala 254:34]
  wire  _GEN_141; // @[TLB.scala 254:34]
  wire  _GEN_142; // @[TLB.scala 254:34]
  wire  _GEN_143; // @[TLB.scala 251:82]
  wire  _GEN_144; // @[TLB.scala 251:82]
  wire  _GEN_145; // @[TLB.scala 251:82]
  wire  _GEN_146; // @[TLB.scala 251:82]
  wire  _T_15; // @[TLB.scala 251:75]
  wire  _GEN_153; // @[TLB.scala 252:32]
  wire  _GEN_154; // @[TLB.scala 252:32]
  wire  _GEN_155; // @[TLB.scala 252:32]
  wire  _GEN_156; // @[TLB.scala 252:32]
  wire  _GEN_157; // @[TLB.scala 121:16]
  wire  _GEN_158; // @[TLB.scala 121:16]
  wire  _GEN_159; // @[TLB.scala 121:16]
  wire  _GEN_160; // @[TLB.scala 121:16]
  wire  _GEN_165; // @[TLB.scala 254:34]
  wire  _GEN_166; // @[TLB.scala 254:34]
  wire  _GEN_167; // @[TLB.scala 254:34]
  wire  _GEN_168; // @[TLB.scala 254:34]
  wire  _GEN_169; // @[TLB.scala 251:82]
  wire  _GEN_170; // @[TLB.scala 251:82]
  wire  _GEN_171; // @[TLB.scala 251:82]
  wire  _GEN_172; // @[TLB.scala 251:82]
  wire  _T_17; // @[TLB.scala 251:75]
  wire  _GEN_179; // @[TLB.scala 252:32]
  wire  _GEN_180; // @[TLB.scala 252:32]
  wire  _GEN_181; // @[TLB.scala 252:32]
  wire  _GEN_182; // @[TLB.scala 252:32]
  wire  _GEN_183; // @[TLB.scala 121:16]
  wire  _GEN_184; // @[TLB.scala 121:16]
  wire  _GEN_185; // @[TLB.scala 121:16]
  wire  _GEN_186; // @[TLB.scala 121:16]
  wire  _GEN_191; // @[TLB.scala 254:34]
  wire  _GEN_192; // @[TLB.scala 254:34]
  wire  _GEN_193; // @[TLB.scala 254:34]
  wire  _GEN_194; // @[TLB.scala 254:34]
  wire  _GEN_195; // @[TLB.scala 251:82]
  wire  _GEN_196; // @[TLB.scala 251:82]
  wire  _GEN_197; // @[TLB.scala 251:82]
  wire  _GEN_198; // @[TLB.scala 251:82]
  wire  _T_19; // @[TLB.scala 251:75]
  wire  _GEN_205; // @[TLB.scala 252:32]
  wire  _GEN_206; // @[TLB.scala 252:32]
  wire  _GEN_207; // @[TLB.scala 252:32]
  wire  _GEN_208; // @[TLB.scala 252:32]
  wire  _GEN_209; // @[TLB.scala 121:16]
  wire  _GEN_210; // @[TLB.scala 121:16]
  wire  _GEN_211; // @[TLB.scala 121:16]
  wire  _GEN_212; // @[TLB.scala 121:16]
  wire  _GEN_217; // @[TLB.scala 254:34]
  wire  _GEN_218; // @[TLB.scala 254:34]
  wire  _GEN_219; // @[TLB.scala 254:34]
  wire  _GEN_220; // @[TLB.scala 254:34]
  wire  _GEN_221; // @[TLB.scala 251:82]
  wire  _GEN_222; // @[TLB.scala 251:82]
  wire  _GEN_223; // @[TLB.scala 251:82]
  wire  _GEN_224; // @[TLB.scala 251:82]
  wire  _T_21; // @[TLB.scala 251:75]
  wire  _GEN_231; // @[TLB.scala 252:32]
  wire  _GEN_232; // @[TLB.scala 252:32]
  wire  _GEN_233; // @[TLB.scala 252:32]
  wire  _GEN_234; // @[TLB.scala 252:32]
  wire  _GEN_235; // @[TLB.scala 121:16]
  wire  _GEN_236; // @[TLB.scala 121:16]
  wire  _GEN_237; // @[TLB.scala 121:16]
  wire  _GEN_238; // @[TLB.scala 121:16]
  wire  _GEN_243; // @[TLB.scala 254:34]
  wire  _GEN_244; // @[TLB.scala 254:34]
  wire  _GEN_245; // @[TLB.scala 254:34]
  wire  _GEN_246; // @[TLB.scala 254:34]
  wire  _GEN_247; // @[TLB.scala 251:82]
  wire  _GEN_248; // @[TLB.scala 251:82]
  wire  _GEN_249; // @[TLB.scala 251:82]
  wire  _GEN_250; // @[TLB.scala 251:82]
  wire  _GEN_259; // @[TLB.scala 243:54]
  wire  _GEN_263; // @[TLB.scala 243:54]
  wire  _GEN_267; // @[TLB.scala 243:54]
  wire  _GEN_271; // @[TLB.scala 243:54]
  wire  _GEN_273; // @[TLB.scala 243:54]
  wire  _GEN_274; // @[TLB.scala 243:54]
  wire  _GEN_275; // @[TLB.scala 243:54]
  wire  _GEN_276; // @[TLB.scala 243:54]
  wire  _GEN_283; // @[TLB.scala 243:54]
  wire  _GEN_284; // @[TLB.scala 243:54]
  wire  _GEN_285; // @[TLB.scala 243:54]
  wire  _GEN_286; // @[TLB.scala 243:54]
  wire  _GEN_293; // @[TLB.scala 243:54]
  wire  _GEN_294; // @[TLB.scala 243:54]
  wire  _GEN_295; // @[TLB.scala 243:54]
  wire  _GEN_296; // @[TLB.scala 243:54]
  wire  _GEN_303; // @[TLB.scala 243:54]
  wire  _GEN_304; // @[TLB.scala 243:54]
  wire  _GEN_305; // @[TLB.scala 243:54]
  wire  _GEN_306; // @[TLB.scala 243:54]
  wire  _GEN_313; // @[TLB.scala 243:54]
  wire  _GEN_314; // @[TLB.scala 243:54]
  wire  _GEN_315; // @[TLB.scala 243:54]
  wire  _GEN_316; // @[TLB.scala 243:54]
  wire  _GEN_323; // @[TLB.scala 243:54]
  wire  _GEN_324; // @[TLB.scala 243:54]
  wire  _GEN_325; // @[TLB.scala 243:54]
  wire  _GEN_326; // @[TLB.scala 243:54]
  wire  _GEN_333; // @[TLB.scala 243:54]
  wire  _GEN_334; // @[TLB.scala 243:54]
  wire  _GEN_335; // @[TLB.scala 243:54]
  wire  _GEN_336; // @[TLB.scala 243:54]
  wire  _GEN_343; // @[TLB.scala 243:54]
  wire  _GEN_344; // @[TLB.scala 243:54]
  wire  _GEN_345; // @[TLB.scala 243:54]
  wire  _GEN_346; // @[TLB.scala 243:54]
  wire  _GEN_355; // @[TLB.scala 238:68]
  wire  _GEN_359; // @[TLB.scala 238:68]
  wire  _GEN_363; // @[TLB.scala 238:68]
  wire  _GEN_367; // @[TLB.scala 238:68]
  wire  _GEN_371; // @[TLB.scala 238:68]
  wire  _GEN_373; // @[TLB.scala 238:68]
  wire  _GEN_374; // @[TLB.scala 238:68]
  wire  _GEN_375; // @[TLB.scala 238:68]
  wire  _GEN_376; // @[TLB.scala 238:68]
  wire  _GEN_383; // @[TLB.scala 238:68]
  wire  _GEN_384; // @[TLB.scala 238:68]
  wire  _GEN_385; // @[TLB.scala 238:68]
  wire  _GEN_386; // @[TLB.scala 238:68]
  wire  _GEN_393; // @[TLB.scala 238:68]
  wire  _GEN_394; // @[TLB.scala 238:68]
  wire  _GEN_395; // @[TLB.scala 238:68]
  wire  _GEN_396; // @[TLB.scala 238:68]
  wire  _GEN_403; // @[TLB.scala 238:68]
  wire  _GEN_404; // @[TLB.scala 238:68]
  wire  _GEN_405; // @[TLB.scala 238:68]
  wire  _GEN_406; // @[TLB.scala 238:68]
  wire  _GEN_413; // @[TLB.scala 238:68]
  wire  _GEN_414; // @[TLB.scala 238:68]
  wire  _GEN_415; // @[TLB.scala 238:68]
  wire  _GEN_416; // @[TLB.scala 238:68]
  wire  _GEN_423; // @[TLB.scala 238:68]
  wire  _GEN_424; // @[TLB.scala 238:68]
  wire  _GEN_425; // @[TLB.scala 238:68]
  wire  _GEN_426; // @[TLB.scala 238:68]
  wire  _GEN_433; // @[TLB.scala 238:68]
  wire  _GEN_434; // @[TLB.scala 238:68]
  wire  _GEN_435; // @[TLB.scala 238:68]
  wire  _GEN_436; // @[TLB.scala 238:68]
  wire  _GEN_443; // @[TLB.scala 238:68]
  wire  _GEN_444; // @[TLB.scala 238:68]
  wire  _GEN_445; // @[TLB.scala 238:68]
  wire  _GEN_446; // @[TLB.scala 238:68]
  wire  _GEN_455; // @[TLB.scala 218:20]
  wire  _GEN_459; // @[TLB.scala 218:20]
  wire  _GEN_463; // @[TLB.scala 218:20]
  wire  _GEN_467; // @[TLB.scala 218:20]
  wire  _GEN_471; // @[TLB.scala 218:20]
  wire  _GEN_473; // @[TLB.scala 218:20]
  wire  _GEN_474; // @[TLB.scala 218:20]
  wire  _GEN_475; // @[TLB.scala 218:20]
  wire  _GEN_476; // @[TLB.scala 218:20]
  wire  _GEN_483; // @[TLB.scala 218:20]
  wire  _GEN_484; // @[TLB.scala 218:20]
  wire  _GEN_485; // @[TLB.scala 218:20]
  wire  _GEN_486; // @[TLB.scala 218:20]
  wire  _GEN_493; // @[TLB.scala 218:20]
  wire  _GEN_494; // @[TLB.scala 218:20]
  wire  _GEN_495; // @[TLB.scala 218:20]
  wire  _GEN_496; // @[TLB.scala 218:20]
  wire  _GEN_503; // @[TLB.scala 218:20]
  wire  _GEN_504; // @[TLB.scala 218:20]
  wire  _GEN_505; // @[TLB.scala 218:20]
  wire  _GEN_506; // @[TLB.scala 218:20]
  wire  _GEN_513; // @[TLB.scala 218:20]
  wire  _GEN_514; // @[TLB.scala 218:20]
  wire  _GEN_515; // @[TLB.scala 218:20]
  wire  _GEN_516; // @[TLB.scala 218:20]
  wire  _GEN_523; // @[TLB.scala 218:20]
  wire  _GEN_524; // @[TLB.scala 218:20]
  wire  _GEN_525; // @[TLB.scala 218:20]
  wire  _GEN_526; // @[TLB.scala 218:20]
  wire  _GEN_533; // @[TLB.scala 218:20]
  wire  _GEN_534; // @[TLB.scala 218:20]
  wire  _GEN_535; // @[TLB.scala 218:20]
  wire  _GEN_536; // @[TLB.scala 218:20]
  wire  _GEN_543; // @[TLB.scala 218:20]
  wire  _GEN_544; // @[TLB.scala 218:20]
  wire  _GEN_545; // @[TLB.scala 218:20]
  wire  _GEN_546; // @[TLB.scala 218:20]
  wire [34:0] _GEN_554;
  wire [34:0] _GEN_555;
  wire [34:0] _GEN_556;
  wire [34:0] _GEN_558;
  wire [34:0] _GEN_559;
  wire [34:0] _GEN_560;
  wire [34:0] _GEN_562;
  wire [34:0] _GEN_563;
  wire [34:0] _GEN_564;
  wire [34:0] _GEN_566;
  wire [34:0] _GEN_567;
  wire [34:0] _GEN_568;
  wire [34:0] _GEN_570;
  wire [34:0] _GEN_571;
  wire [34:0] _GEN_572;
  wire [34:0] _GEN_574;
  wire [34:0] _GEN_575;
  wire [34:0] _GEN_576;
  wire [34:0] _GEN_578;
  wire [34:0] _GEN_579;
  wire [34:0] _GEN_580;
  wire [34:0] _GEN_582;
  wire [34:0] _GEN_583;
  wire [34:0] _GEN_584;
  wire [1:0] ppn_hi; // @[TLB.scala 105:26]
  wire [26:0] _ppn_T_1; // @[TLB.scala 108:28]
  wire [26:0] _GEN_953; // @[TLB.scala 108:47]
  wire [26:0] _ppn_T_2; // @[TLB.scala 108:47]
  wire [8:0] ppn_lo; // @[TLB.scala 108:58]
  wire [26:0] _ppn_T_4; // @[TLB.scala 108:47]
  wire [8:0] ppn_lo_1; // @[TLB.scala 108:58]
  wire [19:0] _ppn_T_5; // @[Cat.scala 30:58]
  wire [1:0] ppn_hi_2; // @[TLB.scala 105:26]
  wire [26:0] _ppn_T_6; // @[TLB.scala 108:28]
  wire [26:0] _GEN_955; // @[TLB.scala 108:47]
  wire [26:0] _ppn_T_7; // @[TLB.scala 108:47]
  wire [8:0] ppn_lo_2; // @[TLB.scala 108:58]
  wire [26:0] _ppn_T_9; // @[TLB.scala 108:47]
  wire [8:0] ppn_lo_3; // @[TLB.scala 108:58]
  wire [19:0] _ppn_T_10; // @[Cat.scala 30:58]
  wire [1:0] ppn_hi_4; // @[TLB.scala 105:26]
  wire [26:0] _ppn_T_11; // @[TLB.scala 108:28]
  wire [26:0] _GEN_957; // @[TLB.scala 108:47]
  wire [26:0] _ppn_T_12; // @[TLB.scala 108:47]
  wire [8:0] ppn_lo_4; // @[TLB.scala 108:58]
  wire [26:0] _ppn_T_14; // @[TLB.scala 108:47]
  wire [8:0] ppn_lo_5; // @[TLB.scala 108:58]
  wire [19:0] _ppn_T_15; // @[Cat.scala 30:58]
  wire [1:0] ppn_hi_6; // @[TLB.scala 105:26]
  wire [26:0] _ppn_T_16; // @[TLB.scala 108:28]
  wire [26:0] _GEN_959; // @[TLB.scala 108:47]
  wire [26:0] _ppn_T_17; // @[TLB.scala 108:47]
  wire [8:0] ppn_lo_6; // @[TLB.scala 108:58]
  wire [26:0] _ppn_T_19; // @[TLB.scala 108:47]
  wire [8:0] ppn_lo_7; // @[TLB.scala 108:58]
  wire [19:0] _ppn_T_20; // @[Cat.scala 30:58]
  wire [1:0] ppn_hi_8; // @[TLB.scala 105:26]
  wire [26:0] _GEN_961; // @[TLB.scala 108:47]
  wire [26:0] _ppn_T_22; // @[TLB.scala 108:47]
  wire [8:0] ppn_lo_8; // @[TLB.scala 108:58]
  wire [26:0] _ppn_T_24; // @[TLB.scala 108:47]
  wire [8:0] ppn_lo_9; // @[TLB.scala 108:58]
  wire [19:0] _ppn_T_25; // @[Cat.scala 30:58]
  wire [19:0] _ppn_T_27; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_28; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_29; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_30; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_31; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_32; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_33; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_34; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_35; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_36; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_37; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_38; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_39; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_40; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_41; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_42; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_43; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_44; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_45; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_46; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_47; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_48; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_49; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_50; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_51; // @[Mux.scala 27:72]
  wire [19:0] _ppn_T_52; // @[Mux.scala 27:72]
  wire [19:0] ppn; // @[Mux.scala 27:72]
  wire [5:0] ptw_ae_array_lo; // @[Cat.scala 30:58]
  wire [13:0] ptw_ae_array; // @[Cat.scala 30:58]
  wire [5:0] priv_rw_ok_lo; // @[Cat.scala 30:58]
  wire [12:0] _priv_rw_ok_T_2; // @[Cat.scala 30:58]
  wire [12:0] priv_x_ok; // @[TLB.scala 266:22]
  wire [5:0] r_array_lo_1; // @[Cat.scala 30:58]
  wire [12:0] _r_array_T_1; // @[Cat.scala 30:58]
  wire [12:0] x_array_lo_1; // @[TLB.scala 269:39]
  wire [13:0] x_array; // @[Cat.scala 30:58]
  wire [1:0] px_array_hi; // @[Bitwise.scala 72:12]
  wire [5:0] px_array_lo; // @[Cat.scala 30:58]
  wire [13:0] _px_array_T_1; // @[Cat.scala 30:58]
  wire [13:0] px_array; // @[TLB.scala 272:87]
  wire [1:0] c_array_hi; // @[Bitwise.scala 72:12]
  wire [5:0] c_array_lo; // @[Cat.scala 30:58]
  wire [13:0] c_array; // @[Cat.scala 30:58]
  wire [39:0] bad_va_maskedVAddr; // @[TLB.scala 289:43]
  wire  _bad_va_T_1; // @[TLB.scala 290:61]
  wire  _bad_va_T_2; // @[TLB.scala 290:82]
  wire  _bad_va_T_3; // @[TLB.scala 290:67]
  wire  bad_va; // @[TLB.scala 284:117]
  wire [13:0] _pf_inst_array_T; // @[TLB.scala 322:33]
  wire [13:0] pf_inst_array; // @[TLB.scala 322:23]
  wire  tlb_hit; // @[TLB.scala 324:27]
  wire  _tlb_miss_T_1; // @[TLB.scala 325:29]
  wire  tlb_miss; // @[TLB.scala 325:40]
  reg [6:0] state_vec_0; // @[Replacement.scala 305:17]
  reg [31:0] _RAND_98;
  reg [2:0] state_reg_1; // @[Replacement.scala 168:70]
  reg [31:0] _RAND_99;
  wire  _T_23; // @[TLB.scala 329:22]
  wire  _T_24; // @[package.scala 72:59]
  wire  _T_25; // @[package.scala 72:59]
  wire  _T_26; // @[package.scala 72:59]
  wire  _T_27; // @[package.scala 72:59]
  wire  _T_28; // @[package.scala 72:59]
  wire  _T_29; // @[package.scala 72:59]
  wire  _T_30; // @[package.scala 72:59]
  wire [7:0] _T_31; // @[Cat.scala 30:58]
  wire [3:0] hi_1; // @[OneHot.scala 30:18]
  wire [3:0] lo_1; // @[OneHot.scala 31:18]
  wire  hi_2; // @[OneHot.scala 32:14]
  wire [3:0] _T_32; // @[OneHot.scala 32:28]
  wire [1:0] hi_3; // @[OneHot.scala 30:18]
  wire [1:0] lo_2; // @[OneHot.scala 31:18]
  wire  hi_4; // @[OneHot.scala 32:14]
  wire [1:0] _T_33; // @[OneHot.scala 32:28]
  wire  lo_3; // @[CircuitMath.scala 30:8]
  wire [2:0] state_vec_0_touch_way_sized; // @[Cat.scala 30:58]
  wire  state_vec_0_hi_hi; // @[Replacement.scala 196:33]
  wire [2:0] state_vec_0_left_subtree_state; // @[package.scala 154:13]
  wire [2:0] state_vec_0_right_subtree_state; // @[Replacement.scala 198:38]
  wire  state_vec_0_hi_hi_1; // @[Replacement.scala 196:33]
  wire  state_vec_0_left_subtree_state_1; // @[package.scala 154:13]
  wire  state_vec_0_right_subtree_state_1; // @[Replacement.scala 198:38]
  wire  state_vec_0_hi_lo; // @[Replacement.scala 203:16]
  wire  state_vec_0_lo; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_0_T_7; // @[Cat.scala 30:58]
  wire [2:0] state_vec_0_hi_lo_1; // @[Replacement.scala 203:16]
  wire  state_vec_0_left_subtree_state_2; // @[package.scala 154:13]
  wire  state_vec_0_right_subtree_state_2; // @[Replacement.scala 198:38]
  wire  state_vec_0_hi_lo_2; // @[Replacement.scala 203:16]
  wire  state_vec_0_lo_1; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_0_T_15; // @[Cat.scala 30:58]
  wire [2:0] state_vec_0_lo_2; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_0_T_16; // @[Cat.scala 30:58]
  wire  _T_35; // @[package.scala 72:59]
  wire  _T_36; // @[package.scala 72:59]
  wire  _T_37; // @[package.scala 72:59]
  wire [3:0] _T_38; // @[Cat.scala 30:58]
  wire [1:0] hi_6; // @[OneHot.scala 30:18]
  wire [1:0] lo_6; // @[OneHot.scala 31:18]
  wire  hi_7; // @[OneHot.scala 32:14]
  wire [1:0] _T_39; // @[OneHot.scala 32:28]
  wire  lo_7; // @[CircuitMath.scala 30:8]
  wire [1:0] state_reg_touch_way_sized; // @[Cat.scala 30:58]
  wire  state_reg_hi_hi; // @[Replacement.scala 196:33]
  wire  state_reg_left_subtree_state; // @[package.scala 154:13]
  wire  state_reg_right_subtree_state; // @[Replacement.scala 198:38]
  wire  state_reg_hi_lo; // @[Replacement.scala 203:16]
  wire  state_reg_lo; // @[Replacement.scala 206:16]
  wire [2:0] _state_reg_T_6; // @[Cat.scala 30:58]
  wire  multipleHits_leftOne; // @[Misc.scala 180:37]
  wire  multipleHits_leftOne_1; // @[Misc.scala 180:37]
  wire  multipleHits_rightOne; // @[Misc.scala 181:39]
  wire  multipleHits_rightOne_1; // @[Misc.scala 182:16]
  wire  multipleHits_rightTwo; // @[Misc.scala 182:61]
  wire  multipleHits_leftOne_2; // @[Misc.scala 182:16]
  wire  _multipleHits_T_9; // @[Misc.scala 182:61]
  wire  multipleHits_leftTwo; // @[Misc.scala 182:49]
  wire  multipleHits_leftOne_3; // @[Misc.scala 180:37]
  wire  multipleHits_leftOne_4; // @[Misc.scala 180:37]
  wire  multipleHits_rightOne_2; // @[Misc.scala 181:39]
  wire  multipleHits_rightOne_3; // @[Misc.scala 182:16]
  wire  multipleHits_rightTwo_1; // @[Misc.scala 182:61]
  wire  multipleHits_rightOne_4; // @[Misc.scala 182:16]
  wire  _multipleHits_T_18; // @[Misc.scala 182:61]
  wire  multipleHits_rightTwo_2; // @[Misc.scala 182:49]
  wire  multipleHits_leftOne_5; // @[Misc.scala 182:16]
  wire  _multipleHits_T_19; // @[Misc.scala 182:37]
  wire  _multipleHits_T_20; // @[Misc.scala 182:61]
  wire  multipleHits_leftTwo_1; // @[Misc.scala 182:49]
  wire  multipleHits_leftOne_6; // @[Misc.scala 180:37]
  wire  multipleHits_leftOne_7; // @[Misc.scala 180:37]
  wire  multipleHits_rightOne_5; // @[Misc.scala 181:39]
  wire  multipleHits_rightOne_6; // @[Misc.scala 182:16]
  wire  multipleHits_rightTwo_3; // @[Misc.scala 182:61]
  wire  multipleHits_leftOne_8; // @[Misc.scala 182:16]
  wire  _multipleHits_T_30; // @[Misc.scala 182:61]
  wire  multipleHits_leftTwo_2; // @[Misc.scala 182:49]
  wire  multipleHits_leftOne_9; // @[Misc.scala 180:37]
  wire  multipleHits_rightOne_7; // @[Misc.scala 181:39]
  wire  multipleHits_leftOne_10; // @[Misc.scala 182:16]
  wire  multipleHits_leftTwo_3; // @[Misc.scala 182:61]
  wire  multipleHits_leftOne_11; // @[Misc.scala 180:37]
  wire  multipleHits_rightOne_8; // @[Misc.scala 181:39]
  wire  multipleHits_rightOne_9; // @[Misc.scala 182:16]
  wire  multipleHits_rightTwo_4; // @[Misc.scala 182:61]
  wire  multipleHits_rightOne_10; // @[Misc.scala 182:16]
  wire  _multipleHits_T_42; // @[Misc.scala 182:37]
  wire  _multipleHits_T_43; // @[Misc.scala 182:61]
  wire  multipleHits_rightTwo_5; // @[Misc.scala 182:49]
  wire  multipleHits_rightOne_11; // @[Misc.scala 182:16]
  wire  _multipleHits_T_44; // @[Misc.scala 182:37]
  wire  _multipleHits_T_45; // @[Misc.scala 182:61]
  wire  multipleHits_rightTwo_6; // @[Misc.scala 182:49]
  wire  _multipleHits_T_47; // @[Misc.scala 182:37]
  wire  _multipleHits_T_48; // @[Misc.scala 182:61]
  wire  multipleHits; // @[Misc.scala 182:49]
  wire [13:0] _io_resp_pf_inst_T; // @[TLB.scala 344:47]
  wire  _io_resp_pf_inst_T_1; // @[TLB.scala 344:55]
  wire [13:0] _io_resp_ae_inst_T_1; // @[TLB.scala 347:33]
  wire [13:0] _io_resp_cacheable_T; // @[TLB.scala 351:33]
  wire  _io_resp_miss_T; // @[TLB.scala 354:29]
  wire  _T_41; // @[Decoupled.scala 40:37]
  wire  _T_42; // @[TLB.scala 363:25]
  wire  r_superpage_repl_addr_hi; // @[Replacement.scala 243:38]
  wire  r_superpage_repl_addr_lo; // @[Replacement.scala 250:16]
  wire [1:0] _r_superpage_repl_addr_T_2; // @[Cat.scala 30:58]
  wire [3:0] r_superpage_repl_addr_valids; // @[Cat.scala 30:58]
  wire  _r_superpage_repl_addr_T_3; // @[TLB.scala 411:16]
  wire  _r_superpage_repl_addr_T_5; // @[OneHot.scala 47:40]
  wire  _r_superpage_repl_addr_T_6; // @[OneHot.scala 47:40]
  wire  _r_superpage_repl_addr_T_7; // @[OneHot.scala 47:40]
  wire  r_sectored_repl_addr_hi; // @[Replacement.scala 243:38]
  wire  r_sectored_repl_addr_hi_1; // @[Replacement.scala 243:38]
  wire  r_sectored_repl_addr_lo; // @[Replacement.scala 250:16]
  wire [1:0] _r_sectored_repl_addr_T_2; // @[Cat.scala 30:58]
  wire  r_sectored_repl_addr_hi_2; // @[Replacement.scala 243:38]
  wire  r_sectored_repl_addr_lo_1; // @[Replacement.scala 250:16]
  wire [1:0] _r_sectored_repl_addr_T_5; // @[Cat.scala 30:58]
  wire [1:0] r_sectored_repl_addr_lo_2; // @[Replacement.scala 250:16]
  wire [2:0] _r_sectored_repl_addr_T_6; // @[Cat.scala 30:58]
  wire [7:0] r_sectored_repl_addr_valids; // @[Cat.scala 30:58]
  wire  _r_sectored_repl_addr_T_7; // @[TLB.scala 411:16]
  wire  _r_sectored_repl_addr_T_9; // @[OneHot.scala 47:40]
  wire  _r_sectored_repl_addr_T_10; // @[OneHot.scala 47:40]
  wire  _r_sectored_repl_addr_T_11; // @[OneHot.scala 47:40]
  wire  _r_sectored_repl_addr_T_12; // @[OneHot.scala 47:40]
  wire  _r_sectored_repl_addr_T_13; // @[OneHot.scala 47:40]
  wire  _r_sectored_repl_addr_T_14; // @[OneHot.scala 47:40]
  wire  _r_sectored_repl_addr_T_15; // @[OneHot.scala 47:40]
  wire  _T_44; // @[TLB.scala 377:17]
  wire  _T_45; // @[TLB.scala 377:28]
  wire  _T_48; // @[TLB.scala 385:72]
  wire  _T_49; // @[TLB.scala 385:34]
  wire  _T_51; // @[TLB.scala 385:13]
  wire  _T_59; // @[TLB.scala 134:61]
  wire  _GEN_617; // @[TLB.scala 142:19]
  wire  _GEN_618; // @[TLB.scala 142:19]
  wire  _GEN_619; // @[TLB.scala 142:19]
  wire  _GEN_620; // @[TLB.scala 142:19]
  wire  _GEN_621; // @[TLB.scala 388:40]
  wire  _GEN_622; // @[TLB.scala 388:40]
  wire  _GEN_623; // @[TLB.scala 388:40]
  wire  _GEN_624; // @[TLB.scala 388:40]
  wire  _T_198; // @[TLB.scala 134:61]
  wire  _GEN_645; // @[TLB.scala 142:19]
  wire  _GEN_646; // @[TLB.scala 142:19]
  wire  _GEN_647; // @[TLB.scala 142:19]
  wire  _GEN_648; // @[TLB.scala 142:19]
  wire  _GEN_649; // @[TLB.scala 388:40]
  wire  _GEN_650; // @[TLB.scala 388:40]
  wire  _GEN_651; // @[TLB.scala 388:40]
  wire  _GEN_652; // @[TLB.scala 388:40]
  wire  _T_337; // @[TLB.scala 134:61]
  wire  _GEN_673; // @[TLB.scala 142:19]
  wire  _GEN_674; // @[TLB.scala 142:19]
  wire  _GEN_675; // @[TLB.scala 142:19]
  wire  _GEN_676; // @[TLB.scala 142:19]
  wire  _GEN_677; // @[TLB.scala 388:40]
  wire  _GEN_678; // @[TLB.scala 388:40]
  wire  _GEN_679; // @[TLB.scala 388:40]
  wire  _GEN_680; // @[TLB.scala 388:40]
  wire  _T_476; // @[TLB.scala 134:61]
  wire  _GEN_701; // @[TLB.scala 142:19]
  wire  _GEN_702; // @[TLB.scala 142:19]
  wire  _GEN_703; // @[TLB.scala 142:19]
  wire  _GEN_704; // @[TLB.scala 142:19]
  wire  _GEN_705; // @[TLB.scala 388:40]
  wire  _GEN_706; // @[TLB.scala 388:40]
  wire  _GEN_707; // @[TLB.scala 388:40]
  wire  _GEN_708; // @[TLB.scala 388:40]
  wire  _T_615; // @[TLB.scala 134:61]
  wire  _GEN_729; // @[TLB.scala 142:19]
  wire  _GEN_730; // @[TLB.scala 142:19]
  wire  _GEN_731; // @[TLB.scala 142:19]
  wire  _GEN_732; // @[TLB.scala 142:19]
  wire  _GEN_733; // @[TLB.scala 388:40]
  wire  _GEN_734; // @[TLB.scala 388:40]
  wire  _GEN_735; // @[TLB.scala 388:40]
  wire  _GEN_736; // @[TLB.scala 388:40]
  wire  _T_754; // @[TLB.scala 134:61]
  wire  _GEN_757; // @[TLB.scala 142:19]
  wire  _GEN_758; // @[TLB.scala 142:19]
  wire  _GEN_759; // @[TLB.scala 142:19]
  wire  _GEN_760; // @[TLB.scala 142:19]
  wire  _GEN_761; // @[TLB.scala 388:40]
  wire  _GEN_762; // @[TLB.scala 388:40]
  wire  _GEN_763; // @[TLB.scala 388:40]
  wire  _GEN_764; // @[TLB.scala 388:40]
  wire  _T_893; // @[TLB.scala 134:61]
  wire  _GEN_785; // @[TLB.scala 142:19]
  wire  _GEN_786; // @[TLB.scala 142:19]
  wire  _GEN_787; // @[TLB.scala 142:19]
  wire  _GEN_788; // @[TLB.scala 142:19]
  wire  _GEN_789; // @[TLB.scala 388:40]
  wire  _GEN_790; // @[TLB.scala 388:40]
  wire  _GEN_791; // @[TLB.scala 388:40]
  wire  _GEN_792; // @[TLB.scala 388:40]
  wire  _T_1032; // @[TLB.scala 134:61]
  wire  _GEN_813; // @[TLB.scala 142:19]
  wire  _GEN_814; // @[TLB.scala 142:19]
  wire  _GEN_815; // @[TLB.scala 142:19]
  wire  _GEN_816; // @[TLB.scala 142:19]
  wire  _GEN_817; // @[TLB.scala 388:40]
  wire  _GEN_818; // @[TLB.scala 388:40]
  wire  _GEN_819; // @[TLB.scala 388:40]
  wire  _GEN_820; // @[TLB.scala 388:40]
  wire  _GEN_826; // @[TLB.scala 142:19]
  wire  _GEN_827; // @[TLB.scala 388:40]
  wire  _GEN_830; // @[TLB.scala 142:19]
  wire  _GEN_831; // @[TLB.scala 388:40]
  wire  _GEN_834; // @[TLB.scala 142:19]
  wire  _GEN_835; // @[TLB.scala 388:40]
  wire  _GEN_838; // @[TLB.scala 142:19]
  wire  _GEN_839; // @[TLB.scala 388:40]
  wire  _GEN_842; // @[TLB.scala 142:19]
  wire  _GEN_843; // @[TLB.scala 388:40]
  wire  _T_1326; // @[TLB.scala 392:24]
  reg [19:0] TLB_1_state; // @[Register tracking TLB_1 state]
  reg [31:0] _RAND_100;
  reg  TLB_1_cov [0:1048575]; // @[Coverage map for TLB_1]
  reg [31:0] _RAND_101;
  wire  TLB_1_cov_read_data; // @[Coverage map for TLB_1]
  wire [19:0] TLB_1_cov_read_addr; // @[Coverage map for TLB_1]
  wire  TLB_1_cov_write_data; // @[Coverage map for TLB_1]
  wire [19:0] TLB_1_cov_write_addr; // @[Coverage map for TLB_1]
  wire  TLB_1_cov_write_mask; // @[Coverage map for TLB_1]
  wire  TLB_1_cov_write_en; // @[Coverage map for TLB_1]
  reg [29:0] TLB_1_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_102;
  wire  mux_cond_0;
  wire  mux_cond_1;
  wire  mux_cond_2;
  wire  mux_cond_3;
  wire  mux_cond_4;
  wire  mux_cond_5;
  wire  mux_cond_6;
  wire  mux_cond_7;
  wire  mux_cond_8;
  wire  mux_cond_9;
  wire  mux_cond_10;
  wire  mux_cond_11;
  wire  mux_cond_12;
  wire  mux_cond_13;
  wire  mux_cond_14;
  wire  mux_cond_15;
  wire  mux_cond_16;
  wire  mux_cond_17;
  wire  mux_cond_18;
  wire  mux_cond_19;
  wire  mux_cond_20;
  wire  mux_cond_21;
  wire  mux_cond_22;
  wire  mux_cond_23;
  wire  mux_cond_24;
  wire  mux_cond_25;
  wire  mux_cond_26;
  wire  mux_cond_27;
  wire  mux_cond_28;
  wire  mux_cond_29;
  wire  mux_cond_30;
  wire  mux_cond_31;
  wire  mux_cond_32;
  wire  mux_cond_33;
  wire  mux_cond_34;
  wire  mux_cond_35;
  wire  mux_cond_36;
  wire  mux_cond_37;
  wire  mux_cond_38;
  wire  mux_cond_39;
  wire  mux_cond_40;
  wire  mux_cond_41;
  wire  mux_cond_42;
  wire  mux_cond_43;
  wire  mux_cond_44;
  wire  mux_cond_45;
  wire  mux_cond_46;
  wire  mux_cond_47;
  wire  mux_cond_48;
  wire  mux_cond_49;
  wire  mux_cond_50;
  wire  mux_cond_51;
  wire  mux_cond_52;
  wire  mux_cond_53;
  wire  mux_cond_54;
  wire  mux_cond_55;
  wire  mux_cond_56;
  wire  mux_cond_57;
  wire  mux_cond_58;
  wire  mux_cond_59;
  wire  mux_cond_60;
  wire  mux_cond_61;
  wire  mux_cond_62;
  wire  mux_cond_63;
  wire  mux_cond_64;
  wire  mux_cond_65;
  wire  mux_cond_66;
  wire  mux_cond_67;
  wire  mux_cond_68;
  wire  r_sectored_hit_shl;
  wire [19:0] r_sectored_hit_pad;
  wire [10:0] r_sectored_repl_addr_shl;
  wire [19:0] r_sectored_repl_addr_pad;
  wire [1:0] r_superpage_repl_addr_shl;
  wire [19:0] r_superpage_repl_addr_pad;
  wire [13:0] special_entry_valid_0_shl;
  wire [19:0] special_entry_valid_0_pad;
  wire [13:0] special_entry_level_shl;
  wire [19:0] special_entry_level_pad;
  wire [13:0] state_shl;
  wire [19:0] state_pad;
  wire [3:0] r_sectored_hit_addr_shl;
  wire [19:0] r_sectored_hit_addr_pad;
  wire [16:0] mux_cond_0_shl;
  wire [19:0] mux_cond_0_pad;
  wire [10:0] mux_cond_1_shl;
  wire [19:0] mux_cond_1_pad;
  wire [2:0] mux_cond_2_shl;
  wire [19:0] mux_cond_2_pad;
  wire [15:0] mux_cond_3_shl;
  wire [19:0] mux_cond_3_pad;
  wire [4:0] mux_cond_4_shl;
  wire [19:0] mux_cond_4_pad;
  wire [13:0] mux_cond_5_shl;
  wire [19:0] mux_cond_5_pad;
  wire [9:0] mux_cond_6_shl;
  wire [19:0] mux_cond_6_pad;
  wire [8:0] mux_cond_7_shl;
  wire [19:0] mux_cond_7_pad;
  wire [12:0] mux_cond_8_shl;
  wire [19:0] mux_cond_8_pad;
  wire [19:0] mux_cond_9_shl;
  wire [19:0] mux_cond_9_pad;
  wire [18:0] mux_cond_10_shl;
  wire [19:0] mux_cond_10_pad;
  wire [9:0] mux_cond_11_shl;
  wire [19:0] mux_cond_11_pad;
  wire [19:0] mux_cond_12_shl;
  wire [19:0] mux_cond_12_pad;
  wire [7:0] mux_cond_13_shl;
  wire [19:0] mux_cond_13_pad;
  wire [11:0] mux_cond_14_shl;
  wire [19:0] mux_cond_14_pad;
  wire  mux_cond_15_shl;
  wire [19:0] mux_cond_15_pad;
  wire [4:0] mux_cond_16_shl;
  wire [19:0] mux_cond_16_pad;
  wire [19:0] mux_cond_17_shl;
  wire [19:0] mux_cond_17_pad;
  wire [9:0] mux_cond_18_shl;
  wire [19:0] mux_cond_18_pad;
  wire [8:0] mux_cond_19_shl;
  wire [19:0] mux_cond_19_pad;
  wire [4:0] mux_cond_20_shl;
  wire [19:0] mux_cond_20_pad;
  wire [6:0] mux_cond_21_shl;
  wire [19:0] mux_cond_21_pad;
  wire [11:0] mux_cond_22_shl;
  wire [19:0] mux_cond_22_pad;
  wire [14:0] mux_cond_23_shl;
  wire [19:0] mux_cond_23_pad;
  wire [7:0] mux_cond_24_shl;
  wire [19:0] mux_cond_24_pad;
  wire [7:0] mux_cond_25_shl;
  wire [19:0] mux_cond_25_pad;
  wire [19:0] mux_cond_26_shl;
  wire [19:0] mux_cond_26_pad;
  wire [10:0] mux_cond_27_shl;
  wire [19:0] mux_cond_27_pad;
  wire [17:0] mux_cond_28_shl;
  wire [19:0] mux_cond_28_pad;
  wire [3:0] mux_cond_29_shl;
  wire [19:0] mux_cond_29_pad;
  wire [9:0] mux_cond_30_shl;
  wire [19:0] mux_cond_30_pad;
  wire [15:0] mux_cond_31_shl;
  wire [19:0] mux_cond_31_pad;
  wire  mux_cond_32_shl;
  wire [19:0] mux_cond_32_pad;
  wire [12:0] mux_cond_33_shl;
  wire [19:0] mux_cond_33_pad;
  wire [17:0] mux_cond_34_shl;
  wire [19:0] mux_cond_34_pad;
  wire [9:0] mux_cond_35_shl;
  wire [19:0] mux_cond_35_pad;
  wire [12:0] mux_cond_36_shl;
  wire [19:0] mux_cond_36_pad;
  wire  mux_cond_37_shl;
  wire [19:0] mux_cond_37_pad;
  wire [5:0] mux_cond_38_shl;
  wire [19:0] mux_cond_38_pad;
  wire [2:0] mux_cond_39_shl;
  wire [19:0] mux_cond_39_pad;
  wire [18:0] mux_cond_40_shl;
  wire [19:0] mux_cond_40_pad;
  wire [13:0] mux_cond_41_shl;
  wire [19:0] mux_cond_41_pad;
  wire [5:0] mux_cond_42_shl;
  wire [19:0] mux_cond_42_pad;
  wire [18:0] mux_cond_43_shl;
  wire [19:0] mux_cond_43_pad;
  wire [18:0] mux_cond_44_shl;
  wire [19:0] mux_cond_44_pad;
  wire [2:0] mux_cond_45_shl;
  wire [19:0] mux_cond_45_pad;
  wire [12:0] mux_cond_46_shl;
  wire [19:0] mux_cond_46_pad;
  wire [18:0] mux_cond_47_shl;
  wire [19:0] mux_cond_47_pad;
  wire [16:0] mux_cond_48_shl;
  wire [19:0] mux_cond_48_pad;
  wire  mux_cond_49_shl;
  wire [19:0] mux_cond_49_pad;
  wire [4:0] mux_cond_50_shl;
  wire [19:0] mux_cond_50_pad;
  wire [9:0] mux_cond_51_shl;
  wire [19:0] mux_cond_51_pad;
  wire [13:0] mux_cond_52_shl;
  wire [19:0] mux_cond_52_pad;
  wire [4:0] mux_cond_53_shl;
  wire [19:0] mux_cond_53_pad;
  wire [5:0] mux_cond_54_shl;
  wire [19:0] mux_cond_54_pad;
  wire [10:0] mux_cond_55_shl;
  wire [19:0] mux_cond_55_pad;
  wire [12:0] mux_cond_56_shl;
  wire [19:0] mux_cond_56_pad;
  wire [4:0] mux_cond_57_shl;
  wire [19:0] mux_cond_57_pad;
  wire [19:0] mux_cond_58_shl;
  wire [19:0] mux_cond_58_pad;
  wire [8:0] mux_cond_59_shl;
  wire [19:0] mux_cond_59_pad;
  wire [12:0] mux_cond_60_shl;
  wire [19:0] mux_cond_60_pad;
  wire [13:0] mux_cond_61_shl;
  wire [19:0] mux_cond_61_pad;
  wire [19:0] mux_cond_62_shl;
  wire [19:0] mux_cond_62_pad;
  wire [7:0] mux_cond_63_shl;
  wire [19:0] mux_cond_63_pad;
  wire [1:0] mux_cond_64_shl;
  wire [19:0] mux_cond_64_pad;
  wire [3:0] mux_cond_65_shl;
  wire [19:0] mux_cond_65_pad;
  wire [1:0] mux_cond_66_shl;
  wire [19:0] mux_cond_66_pad;
  wire [15:0] mux_cond_67_shl;
  wire [19:0] mux_cond_67_pad;
  wire [15:0] mux_cond_68_shl;
  wire [19:0] mux_cond_68_pad;
  wire [5:0] sectored_entries_0_0_valid_3_shl;
  wire [19:0] sectored_entries_0_0_valid_3_pad;
  wire [4:0] sectored_entries_0_0_valid_2_shl;
  wire [19:0] sectored_entries_0_0_valid_2_pad;
  wire [5:0] sectored_entries_0_2_valid_0_shl;
  wire [19:0] sectored_entries_0_2_valid_0_pad;
  wire [5:0] sectored_entries_0_3_valid_0_shl;
  wire [19:0] sectored_entries_0_3_valid_0_pad;
  wire [14:0] superpage_entries_2_level_shl;
  wire [19:0] superpage_entries_2_level_pad;
  wire [4:0] sectored_entries_0_7_valid_1_shl;
  wire [19:0] sectored_entries_0_7_valid_1_pad;
  wire [5:0] sectored_entries_0_4_valid_0_shl;
  wire [19:0] sectored_entries_0_4_valid_0_pad;
  wire [5:0] sectored_entries_0_1_valid_3_shl;
  wire [19:0] sectored_entries_0_1_valid_3_pad;
  wire [4:0] sectored_entries_0_1_valid_1_shl;
  wire [19:0] sectored_entries_0_1_valid_1_pad;
  wire [5:0] sectored_entries_0_2_valid_3_shl;
  wire [19:0] sectored_entries_0_2_valid_3_pad;
  wire [4:0] sectored_entries_0_2_valid_1_shl;
  wire [19:0] sectored_entries_0_2_valid_1_pad;
  wire [1:0] superpage_entries_1_valid_0_shl;
  wire [19:0] superpage_entries_1_valid_0_pad;
  wire [5:0] sectored_entries_0_7_valid_0_shl;
  wire [19:0] sectored_entries_0_7_valid_0_pad;
  wire [1:0] superpage_entries_3_valid_0_shl;
  wire [19:0] superpage_entries_3_valid_0_pad;
  wire [5:0] sectored_entries_0_5_valid_3_shl;
  wire [19:0] sectored_entries_0_5_valid_3_pad;
  wire [4:0] sectored_entries_0_5_valid_1_shl;
  wire [19:0] sectored_entries_0_5_valid_1_pad;
  wire [5:0] sectored_entries_0_4_valid_3_shl;
  wire [19:0] sectored_entries_0_4_valid_3_pad;
  wire [4:0] sectored_entries_0_5_valid_2_shl;
  wire [19:0] sectored_entries_0_5_valid_2_pad;
  wire [4:0] sectored_entries_0_1_valid_2_shl;
  wire [19:0] sectored_entries_0_1_valid_2_pad;
  wire [4:0] sectored_entries_0_3_valid_1_shl;
  wire [19:0] sectored_entries_0_3_valid_1_pad;
  wire [5:0] sectored_entries_0_1_valid_0_shl;
  wire [19:0] sectored_entries_0_1_valid_0_pad;
  wire [4:0] sectored_entries_0_4_valid_2_shl;
  wire [19:0] sectored_entries_0_4_valid_2_pad;
  wire [4:0] sectored_entries_0_4_valid_1_shl;
  wire [19:0] sectored_entries_0_4_valid_1_pad;
  wire [14:0] superpage_entries_3_level_shl;
  wire [19:0] superpage_entries_3_level_pad;
  wire [4:0] sectored_entries_0_0_valid_1_shl;
  wire [19:0] sectored_entries_0_0_valid_1_pad;
  wire [4:0] sectored_entries_0_3_valid_2_shl;
  wire [19:0] sectored_entries_0_3_valid_2_pad;
  wire [4:0] sectored_entries_0_6_valid_1_shl;
  wire [19:0] sectored_entries_0_6_valid_1_pad;
  wire [5:0] sectored_entries_0_7_valid_3_shl;
  wire [19:0] sectored_entries_0_7_valid_3_pad;
  wire [5:0] sectored_entries_0_3_valid_3_shl;
  wire [19:0] sectored_entries_0_3_valid_3_pad;
  wire [5:0] sectored_entries_0_0_valid_0_shl;
  wire [19:0] sectored_entries_0_0_valid_0_pad;
  wire [1:0] superpage_entries_0_valid_0_shl;
  wire [19:0] superpage_entries_0_valid_0_pad;
  wire [4:0] sectored_entries_0_2_valid_2_shl;
  wire [19:0] sectored_entries_0_2_valid_2_pad;
  wire [4:0] sectored_entries_0_6_valid_2_shl;
  wire [19:0] sectored_entries_0_6_valid_2_pad;
  wire [1:0] superpage_entries_2_valid_0_shl;
  wire [19:0] superpage_entries_2_valid_0_pad;
  wire [5:0] sectored_entries_0_6_valid_3_shl;
  wire [19:0] sectored_entries_0_6_valid_3_pad;
  wire [5:0] sectored_entries_0_6_valid_0_shl;
  wire [19:0] sectored_entries_0_6_valid_0_pad;
  wire [4:0] sectored_entries_0_7_valid_2_shl;
  wire [19:0] sectored_entries_0_7_valid_2_pad;
  wire [14:0] superpage_entries_0_level_shl;
  wire [19:0] superpage_entries_0_level_pad;
  wire [14:0] superpage_entries_1_level_shl;
  wire [19:0] superpage_entries_1_level_pad;
  wire [5:0] sectored_entries_0_5_valid_0_shl;
  wire [19:0] sectored_entries_0_5_valid_0_pad;
  wire [19:0] TLB_1_xor64;
  wire [19:0] TLB_1_xor31;
  wire [19:0] TLB_1_xor65;
  wire [19:0] TLB_1_xor66;
  wire [19:0] TLB_1_xor32;
  wire [19:0] TLB_1_xor15;
  wire [19:0] TLB_1_xor68;
  wire [19:0] TLB_1_xor33;
  wire [19:0] TLB_1_xor69;
  wire [19:0] TLB_1_xor70;
  wire [19:0] TLB_1_xor34;
  wire [19:0] TLB_1_xor16;
  wire [19:0] TLB_1_xor7;
  wire [19:0] TLB_1_xor72;
  wire [19:0] TLB_1_xor35;
  wire [19:0] TLB_1_xor73;
  wire [19:0] TLB_1_xor74;
  wire [19:0] TLB_1_xor36;
  wire [19:0] TLB_1_xor17;
  wire [19:0] TLB_1_xor75;
  wire [19:0] TLB_1_xor76;
  wire [19:0] TLB_1_xor37;
  wire [19:0] TLB_1_xor77;
  wire [19:0] TLB_1_xor78;
  wire [19:0] TLB_1_xor38;
  wire [19:0] TLB_1_xor18;
  wire [19:0] TLB_1_xor8;
  wire [19:0] TLB_1_xor3;
  wire [19:0] TLB_1_xor80;
  wire [19:0] TLB_1_xor39;
  wire [19:0] TLB_1_xor81;
  wire [19:0] TLB_1_xor82;
  wire [19:0] TLB_1_xor40;
  wire [19:0] TLB_1_xor19;
  wire [19:0] TLB_1_xor84;
  wire [19:0] TLB_1_xor41;
  wire [19:0] TLB_1_xor85;
  wire [19:0] TLB_1_xor86;
  wire [19:0] TLB_1_xor42;
  wire [19:0] TLB_1_xor20;
  wire [19:0] TLB_1_xor9;
  wire [19:0] TLB_1_xor88;
  wire [19:0] TLB_1_xor43;
  wire [19:0] TLB_1_xor89;
  wire [19:0] TLB_1_xor90;
  wire [19:0] TLB_1_xor44;
  wire [19:0] TLB_1_xor21;
  wire [19:0] TLB_1_xor91;
  wire [19:0] TLB_1_xor92;
  wire [19:0] TLB_1_xor45;
  wire [19:0] TLB_1_xor93;
  wire [19:0] TLB_1_xor94;
  wire [19:0] TLB_1_xor46;
  wire [19:0] TLB_1_xor22;
  wire [19:0] TLB_1_xor10;
  wire [19:0] TLB_1_xor4;
  wire [19:0] TLB_1_xor1;
  wire [19:0] TLB_1_xor96;
  wire [19:0] TLB_1_xor47;
  wire [19:0] TLB_1_xor97;
  wire [19:0] TLB_1_xor98;
  wire [19:0] TLB_1_xor48;
  wire [19:0] TLB_1_xor23;
  wire [19:0] TLB_1_xor100;
  wire [19:0] TLB_1_xor49;
  wire [19:0] TLB_1_xor101;
  wire [19:0] TLB_1_xor102;
  wire [19:0] TLB_1_xor50;
  wire [19:0] TLB_1_xor24;
  wire [19:0] TLB_1_xor11;
  wire [19:0] TLB_1_xor104;
  wire [19:0] TLB_1_xor51;
  wire [19:0] TLB_1_xor105;
  wire [19:0] TLB_1_xor106;
  wire [19:0] TLB_1_xor52;
  wire [19:0] TLB_1_xor25;
  wire [19:0] TLB_1_xor107;
  wire [19:0] TLB_1_xor108;
  wire [19:0] TLB_1_xor53;
  wire [19:0] TLB_1_xor109;
  wire [19:0] TLB_1_xor110;
  wire [19:0] TLB_1_xor54;
  wire [19:0] TLB_1_xor26;
  wire [19:0] TLB_1_xor12;
  wire [19:0] TLB_1_xor5;
  wire [19:0] TLB_1_xor112;
  wire [19:0] TLB_1_xor55;
  wire [19:0] TLB_1_xor113;
  wire [19:0] TLB_1_xor114;
  wire [19:0] TLB_1_xor56;
  wire [19:0] TLB_1_xor27;
  wire [19:0] TLB_1_xor116;
  wire [19:0] TLB_1_xor57;
  wire [19:0] TLB_1_xor117;
  wire [19:0] TLB_1_xor118;
  wire [19:0] TLB_1_xor58;
  wire [19:0] TLB_1_xor28;
  wire [19:0] TLB_1_xor13;
  wire [19:0] TLB_1_xor120;
  wire [19:0] TLB_1_xor59;
  wire [19:0] TLB_1_xor121;
  wire [19:0] TLB_1_xor122;
  wire [19:0] TLB_1_xor60;
  wire [19:0] TLB_1_xor29;
  wire [19:0] TLB_1_xor123;
  wire [19:0] TLB_1_xor124;
  wire [19:0] TLB_1_xor61;
  wire [19:0] TLB_1_xor125;
  wire [19:0] TLB_1_xor126;
  wire [19:0] TLB_1_xor62;
  wire [19:0] TLB_1_xor30;
  wire [19:0] TLB_1_xor14;
  wire [19:0] TLB_1_xor6;
  wire [19:0] TLB_1_xor2;
  wire [19:0] TLB_1_xor0;
  wire [29:0] mpu_ppn_barrier_sum;
  wire [29:0] entries_barrier_10_sum;
  wire [29:0] entries_barrier_9_sum;
  wire [29:0] entries_barrier_7_sum;
  wire [29:0] entries_barrier_sum;
  wire [29:0] pmp_sum;
  wire [29:0] entries_barrier_6_sum;
  wire [29:0] entries_barrier_12_sum;
  wire [29:0] entries_barrier_1_sum;
  wire [29:0] entries_barrier_11_sum;
  wire [29:0] entries_barrier_8_sum;
  wire [29:0] entries_barrier_2_sum;
  wire [29:0] entries_barrier_4_sum;
  wire [29:0] entries_barrier_5_sum;
  wire [29:0] entries_barrier_3_sum;
  wire  stopEn0;
  wire  entries_barrier_11_metaAssert_wire;
  wire  entries_barrier_8_metaAssert_wire;
  wire  entries_barrier_3_metaAssert_wire;
  wire  pmp_metaAssert_wire;
  wire  entries_barrier_6_metaAssert_wire;
  wire  entries_barrier_12_metaAssert_wire;
  wire  entries_barrier_9_metaAssert_wire;
  wire  mpu_ppn_barrier_metaAssert_wire;
  wire  entries_barrier_7_metaAssert_wire;
  wire  entries_barrier_metaAssert_wire;
  wire  entries_barrier_5_metaAssert_wire;
  wire  entries_barrier_2_metaAssert_wire;
  wire  entries_barrier_4_metaAssert_wire;
  wire  entries_barrier_1_metaAssert_wire;
  wire  entries_barrier_10_metaAssert_wire;
  wire  TLB_1_or7;
  wire  TLB_1_or8;
  wire  TLB_1_or3;
  wire  TLB_1_or9;
  wire  TLB_1_or10;
  wire  TLB_1_or4;
  wire  TLB_1_or1;
  wire  TLB_1_or11;
  wire  TLB_1_or12;
  wire  TLB_1_or5;
  wire  TLB_1_or13;
  wire  TLB_1_or14;
  wire  TLB_1_or6;
  wire  TLB_1_or2;
  wire  TLB_1_or0;
  reg  TLB_1_metaAssert;
  reg [31:0] _RAND_103;
  OptimizationBarrier mpu_ppn_barrier ( // @[package.scala 258:25]
    .io_x_ppn(mpu_ppn_barrier_io_x_ppn),
    .io_x_u(mpu_ppn_barrier_io_x_u),
    .io_x_ae(mpu_ppn_barrier_io_x_ae),
    .io_x_sw(mpu_ppn_barrier_io_x_sw),
    .io_x_sx(mpu_ppn_barrier_io_x_sx),
    .io_x_sr(mpu_ppn_barrier_io_x_sr),
    .io_x_pw(mpu_ppn_barrier_io_x_pw),
    .io_x_px(mpu_ppn_barrier_io_x_px),
    .io_x_pr(mpu_ppn_barrier_io_x_pr),
    .io_x_ppp(mpu_ppn_barrier_io_x_ppp),
    .io_x_pal(mpu_ppn_barrier_io_x_pal),
    .io_x_paa(mpu_ppn_barrier_io_x_paa),
    .io_x_eff(mpu_ppn_barrier_io_x_eff),
    .io_x_c(mpu_ppn_barrier_io_x_c),
    .io_y_ppn(mpu_ppn_barrier_io_y_ppn),
    .io_y_u(mpu_ppn_barrier_io_y_u),
    .io_y_ae(mpu_ppn_barrier_io_y_ae),
    .io_y_sw(mpu_ppn_barrier_io_y_sw),
    .io_y_sx(mpu_ppn_barrier_io_y_sx),
    .io_y_sr(mpu_ppn_barrier_io_y_sr),
    .io_y_pw(mpu_ppn_barrier_io_y_pw),
    .io_y_px(mpu_ppn_barrier_io_y_px),
    .io_y_pr(mpu_ppn_barrier_io_y_pr),
    .io_y_ppp(mpu_ppn_barrier_io_y_ppp),
    .io_y_pal(mpu_ppn_barrier_io_y_pal),
    .io_y_paa(mpu_ppn_barrier_io_y_paa),
    .io_y_eff(mpu_ppn_barrier_io_y_eff),
    .io_y_c(mpu_ppn_barrier_io_y_c),
    .io_covSum(mpu_ppn_barrier_io_covSum),
    .metaAssert(mpu_ppn_barrier_metaAssert)
  );
  PMPChecker_2 pmp ( // @[TLB.scala 192:19]
    .io_prv(pmp_io_prv),
    .io_pmp_0_cfg_l(pmp_io_pmp_0_cfg_l),
    .io_pmp_0_cfg_a(pmp_io_pmp_0_cfg_a),
    .io_pmp_0_cfg_x(pmp_io_pmp_0_cfg_x),
    .io_pmp_0_cfg_w(pmp_io_pmp_0_cfg_w),
    .io_pmp_0_cfg_r(pmp_io_pmp_0_cfg_r),
    .io_pmp_0_addr(pmp_io_pmp_0_addr),
    .io_pmp_0_mask(pmp_io_pmp_0_mask),
    .io_pmp_1_cfg_l(pmp_io_pmp_1_cfg_l),
    .io_pmp_1_cfg_a(pmp_io_pmp_1_cfg_a),
    .io_pmp_1_cfg_x(pmp_io_pmp_1_cfg_x),
    .io_pmp_1_cfg_w(pmp_io_pmp_1_cfg_w),
    .io_pmp_1_cfg_r(pmp_io_pmp_1_cfg_r),
    .io_pmp_1_addr(pmp_io_pmp_1_addr),
    .io_pmp_1_mask(pmp_io_pmp_1_mask),
    .io_pmp_2_cfg_l(pmp_io_pmp_2_cfg_l),
    .io_pmp_2_cfg_a(pmp_io_pmp_2_cfg_a),
    .io_pmp_2_cfg_x(pmp_io_pmp_2_cfg_x),
    .io_pmp_2_cfg_w(pmp_io_pmp_2_cfg_w),
    .io_pmp_2_cfg_r(pmp_io_pmp_2_cfg_r),
    .io_pmp_2_addr(pmp_io_pmp_2_addr),
    .io_pmp_2_mask(pmp_io_pmp_2_mask),
    .io_pmp_3_cfg_l(pmp_io_pmp_3_cfg_l),
    .io_pmp_3_cfg_a(pmp_io_pmp_3_cfg_a),
    .io_pmp_3_cfg_x(pmp_io_pmp_3_cfg_x),
    .io_pmp_3_cfg_w(pmp_io_pmp_3_cfg_w),
    .io_pmp_3_cfg_r(pmp_io_pmp_3_cfg_r),
    .io_pmp_3_addr(pmp_io_pmp_3_addr),
    .io_pmp_3_mask(pmp_io_pmp_3_mask),
    .io_pmp_4_cfg_l(pmp_io_pmp_4_cfg_l),
    .io_pmp_4_cfg_a(pmp_io_pmp_4_cfg_a),
    .io_pmp_4_cfg_x(pmp_io_pmp_4_cfg_x),
    .io_pmp_4_cfg_w(pmp_io_pmp_4_cfg_w),
    .io_pmp_4_cfg_r(pmp_io_pmp_4_cfg_r),
    .io_pmp_4_addr(pmp_io_pmp_4_addr),
    .io_pmp_4_mask(pmp_io_pmp_4_mask),
    .io_pmp_5_cfg_l(pmp_io_pmp_5_cfg_l),
    .io_pmp_5_cfg_a(pmp_io_pmp_5_cfg_a),
    .io_pmp_5_cfg_x(pmp_io_pmp_5_cfg_x),
    .io_pmp_5_cfg_w(pmp_io_pmp_5_cfg_w),
    .io_pmp_5_cfg_r(pmp_io_pmp_5_cfg_r),
    .io_pmp_5_addr(pmp_io_pmp_5_addr),
    .io_pmp_5_mask(pmp_io_pmp_5_mask),
    .io_pmp_6_cfg_l(pmp_io_pmp_6_cfg_l),
    .io_pmp_6_cfg_a(pmp_io_pmp_6_cfg_a),
    .io_pmp_6_cfg_x(pmp_io_pmp_6_cfg_x),
    .io_pmp_6_cfg_w(pmp_io_pmp_6_cfg_w),
    .io_pmp_6_cfg_r(pmp_io_pmp_6_cfg_r),
    .io_pmp_6_addr(pmp_io_pmp_6_addr),
    .io_pmp_6_mask(pmp_io_pmp_6_mask),
    .io_pmp_7_cfg_l(pmp_io_pmp_7_cfg_l),
    .io_pmp_7_cfg_a(pmp_io_pmp_7_cfg_a),
    .io_pmp_7_cfg_x(pmp_io_pmp_7_cfg_x),
    .io_pmp_7_cfg_w(pmp_io_pmp_7_cfg_w),
    .io_pmp_7_cfg_r(pmp_io_pmp_7_cfg_r),
    .io_pmp_7_addr(pmp_io_pmp_7_addr),
    .io_pmp_7_mask(pmp_io_pmp_7_mask),
    .io_addr(pmp_io_addr),
    .io_r(pmp_io_r),
    .io_w(pmp_io_w),
    .io_x(pmp_io_x),
    .io_covSum(pmp_io_covSum),
    .metaAssert(pmp_metaAssert)
  );
  OptimizationBarrier entries_barrier ( // @[package.scala 258:25]
    .io_x_ppn(entries_barrier_io_x_ppn),
    .io_x_u(entries_barrier_io_x_u),
    .io_x_ae(entries_barrier_io_x_ae),
    .io_x_sw(entries_barrier_io_x_sw),
    .io_x_sx(entries_barrier_io_x_sx),
    .io_x_sr(entries_barrier_io_x_sr),
    .io_x_pw(entries_barrier_io_x_pw),
    .io_x_px(entries_barrier_io_x_px),
    .io_x_pr(entries_barrier_io_x_pr),
    .io_x_ppp(entries_barrier_io_x_ppp),
    .io_x_pal(entries_barrier_io_x_pal),
    .io_x_paa(entries_barrier_io_x_paa),
    .io_x_eff(entries_barrier_io_x_eff),
    .io_x_c(entries_barrier_io_x_c),
    .io_y_ppn(entries_barrier_io_y_ppn),
    .io_y_u(entries_barrier_io_y_u),
    .io_y_ae(entries_barrier_io_y_ae),
    .io_y_sw(entries_barrier_io_y_sw),
    .io_y_sx(entries_barrier_io_y_sx),
    .io_y_sr(entries_barrier_io_y_sr),
    .io_y_pw(entries_barrier_io_y_pw),
    .io_y_px(entries_barrier_io_y_px),
    .io_y_pr(entries_barrier_io_y_pr),
    .io_y_ppp(entries_barrier_io_y_ppp),
    .io_y_pal(entries_barrier_io_y_pal),
    .io_y_paa(entries_barrier_io_y_paa),
    .io_y_eff(entries_barrier_io_y_eff),
    .io_y_c(entries_barrier_io_y_c),
    .io_covSum(entries_barrier_io_covSum),
    .metaAssert(entries_barrier_metaAssert)
  );
  OptimizationBarrier entries_barrier_1 ( // @[package.scala 258:25]
    .io_x_ppn(entries_barrier_1_io_x_ppn),
    .io_x_u(entries_barrier_1_io_x_u),
    .io_x_ae(entries_barrier_1_io_x_ae),
    .io_x_sw(entries_barrier_1_io_x_sw),
    .io_x_sx(entries_barrier_1_io_x_sx),
    .io_x_sr(entries_barrier_1_io_x_sr),
    .io_x_pw(entries_barrier_1_io_x_pw),
    .io_x_px(entries_barrier_1_io_x_px),
    .io_x_pr(entries_barrier_1_io_x_pr),
    .io_x_ppp(entries_barrier_1_io_x_ppp),
    .io_x_pal(entries_barrier_1_io_x_pal),
    .io_x_paa(entries_barrier_1_io_x_paa),
    .io_x_eff(entries_barrier_1_io_x_eff),
    .io_x_c(entries_barrier_1_io_x_c),
    .io_y_ppn(entries_barrier_1_io_y_ppn),
    .io_y_u(entries_barrier_1_io_y_u),
    .io_y_ae(entries_barrier_1_io_y_ae),
    .io_y_sw(entries_barrier_1_io_y_sw),
    .io_y_sx(entries_barrier_1_io_y_sx),
    .io_y_sr(entries_barrier_1_io_y_sr),
    .io_y_pw(entries_barrier_1_io_y_pw),
    .io_y_px(entries_barrier_1_io_y_px),
    .io_y_pr(entries_barrier_1_io_y_pr),
    .io_y_ppp(entries_barrier_1_io_y_ppp),
    .io_y_pal(entries_barrier_1_io_y_pal),
    .io_y_paa(entries_barrier_1_io_y_paa),
    .io_y_eff(entries_barrier_1_io_y_eff),
    .io_y_c(entries_barrier_1_io_y_c),
    .io_covSum(entries_barrier_1_io_covSum),
    .metaAssert(entries_barrier_1_metaAssert)
  );
  OptimizationBarrier entries_barrier_2 ( // @[package.scala 258:25]
    .io_x_ppn(entries_barrier_2_io_x_ppn),
    .io_x_u(entries_barrier_2_io_x_u),
    .io_x_ae(entries_barrier_2_io_x_ae),
    .io_x_sw(entries_barrier_2_io_x_sw),
    .io_x_sx(entries_barrier_2_io_x_sx),
    .io_x_sr(entries_barrier_2_io_x_sr),
    .io_x_pw(entries_barrier_2_io_x_pw),
    .io_x_px(entries_barrier_2_io_x_px),
    .io_x_pr(entries_barrier_2_io_x_pr),
    .io_x_ppp(entries_barrier_2_io_x_ppp),
    .io_x_pal(entries_barrier_2_io_x_pal),
    .io_x_paa(entries_barrier_2_io_x_paa),
    .io_x_eff(entries_barrier_2_io_x_eff),
    .io_x_c(entries_barrier_2_io_x_c),
    .io_y_ppn(entries_barrier_2_io_y_ppn),
    .io_y_u(entries_barrier_2_io_y_u),
    .io_y_ae(entries_barrier_2_io_y_ae),
    .io_y_sw(entries_barrier_2_io_y_sw),
    .io_y_sx(entries_barrier_2_io_y_sx),
    .io_y_sr(entries_barrier_2_io_y_sr),
    .io_y_pw(entries_barrier_2_io_y_pw),
    .io_y_px(entries_barrier_2_io_y_px),
    .io_y_pr(entries_barrier_2_io_y_pr),
    .io_y_ppp(entries_barrier_2_io_y_ppp),
    .io_y_pal(entries_barrier_2_io_y_pal),
    .io_y_paa(entries_barrier_2_io_y_paa),
    .io_y_eff(entries_barrier_2_io_y_eff),
    .io_y_c(entries_barrier_2_io_y_c),
    .io_covSum(entries_barrier_2_io_covSum),
    .metaAssert(entries_barrier_2_metaAssert)
  );
  OptimizationBarrier entries_barrier_3 ( // @[package.scala 258:25]
    .io_x_ppn(entries_barrier_3_io_x_ppn),
    .io_x_u(entries_barrier_3_io_x_u),
    .io_x_ae(entries_barrier_3_io_x_ae),
    .io_x_sw(entries_barrier_3_io_x_sw),
    .io_x_sx(entries_barrier_3_io_x_sx),
    .io_x_sr(entries_barrier_3_io_x_sr),
    .io_x_pw(entries_barrier_3_io_x_pw),
    .io_x_px(entries_barrier_3_io_x_px),
    .io_x_pr(entries_barrier_3_io_x_pr),
    .io_x_ppp(entries_barrier_3_io_x_ppp),
    .io_x_pal(entries_barrier_3_io_x_pal),
    .io_x_paa(entries_barrier_3_io_x_paa),
    .io_x_eff(entries_barrier_3_io_x_eff),
    .io_x_c(entries_barrier_3_io_x_c),
    .io_y_ppn(entries_barrier_3_io_y_ppn),
    .io_y_u(entries_barrier_3_io_y_u),
    .io_y_ae(entries_barrier_3_io_y_ae),
    .io_y_sw(entries_barrier_3_io_y_sw),
    .io_y_sx(entries_barrier_3_io_y_sx),
    .io_y_sr(entries_barrier_3_io_y_sr),
    .io_y_pw(entries_barrier_3_io_y_pw),
    .io_y_px(entries_barrier_3_io_y_px),
    .io_y_pr(entries_barrier_3_io_y_pr),
    .io_y_ppp(entries_barrier_3_io_y_ppp),
    .io_y_pal(entries_barrier_3_io_y_pal),
    .io_y_paa(entries_barrier_3_io_y_paa),
    .io_y_eff(entries_barrier_3_io_y_eff),
    .io_y_c(entries_barrier_3_io_y_c),
    .io_covSum(entries_barrier_3_io_covSum),
    .metaAssert(entries_barrier_3_metaAssert)
  );
  OptimizationBarrier entries_barrier_4 ( // @[package.scala 258:25]
    .io_x_ppn(entries_barrier_4_io_x_ppn),
    .io_x_u(entries_barrier_4_io_x_u),
    .io_x_ae(entries_barrier_4_io_x_ae),
    .io_x_sw(entries_barrier_4_io_x_sw),
    .io_x_sx(entries_barrier_4_io_x_sx),
    .io_x_sr(entries_barrier_4_io_x_sr),
    .io_x_pw(entries_barrier_4_io_x_pw),
    .io_x_px(entries_barrier_4_io_x_px),
    .io_x_pr(entries_barrier_4_io_x_pr),
    .io_x_ppp(entries_barrier_4_io_x_ppp),
    .io_x_pal(entries_barrier_4_io_x_pal),
    .io_x_paa(entries_barrier_4_io_x_paa),
    .io_x_eff(entries_barrier_4_io_x_eff),
    .io_x_c(entries_barrier_4_io_x_c),
    .io_y_ppn(entries_barrier_4_io_y_ppn),
    .io_y_u(entries_barrier_4_io_y_u),
    .io_y_ae(entries_barrier_4_io_y_ae),
    .io_y_sw(entries_barrier_4_io_y_sw),
    .io_y_sx(entries_barrier_4_io_y_sx),
    .io_y_sr(entries_barrier_4_io_y_sr),
    .io_y_pw(entries_barrier_4_io_y_pw),
    .io_y_px(entries_barrier_4_io_y_px),
    .io_y_pr(entries_barrier_4_io_y_pr),
    .io_y_ppp(entries_barrier_4_io_y_ppp),
    .io_y_pal(entries_barrier_4_io_y_pal),
    .io_y_paa(entries_barrier_4_io_y_paa),
    .io_y_eff(entries_barrier_4_io_y_eff),
    .io_y_c(entries_barrier_4_io_y_c),
    .io_covSum(entries_barrier_4_io_covSum),
    .metaAssert(entries_barrier_4_metaAssert)
  );
  OptimizationBarrier entries_barrier_5 ( // @[package.scala 258:25]
    .io_x_ppn(entries_barrier_5_io_x_ppn),
    .io_x_u(entries_barrier_5_io_x_u),
    .io_x_ae(entries_barrier_5_io_x_ae),
    .io_x_sw(entries_barrier_5_io_x_sw),
    .io_x_sx(entries_barrier_5_io_x_sx),
    .io_x_sr(entries_barrier_5_io_x_sr),
    .io_x_pw(entries_barrier_5_io_x_pw),
    .io_x_px(entries_barrier_5_io_x_px),
    .io_x_pr(entries_barrier_5_io_x_pr),
    .io_x_ppp(entries_barrier_5_io_x_ppp),
    .io_x_pal(entries_barrier_5_io_x_pal),
    .io_x_paa(entries_barrier_5_io_x_paa),
    .io_x_eff(entries_barrier_5_io_x_eff),
    .io_x_c(entries_barrier_5_io_x_c),
    .io_y_ppn(entries_barrier_5_io_y_ppn),
    .io_y_u(entries_barrier_5_io_y_u),
    .io_y_ae(entries_barrier_5_io_y_ae),
    .io_y_sw(entries_barrier_5_io_y_sw),
    .io_y_sx(entries_barrier_5_io_y_sx),
    .io_y_sr(entries_barrier_5_io_y_sr),
    .io_y_pw(entries_barrier_5_io_y_pw),
    .io_y_px(entries_barrier_5_io_y_px),
    .io_y_pr(entries_barrier_5_io_y_pr),
    .io_y_ppp(entries_barrier_5_io_y_ppp),
    .io_y_pal(entries_barrier_5_io_y_pal),
    .io_y_paa(entries_barrier_5_io_y_paa),
    .io_y_eff(entries_barrier_5_io_y_eff),
    .io_y_c(entries_barrier_5_io_y_c),
    .io_covSum(entries_barrier_5_io_covSum),
    .metaAssert(entries_barrier_5_metaAssert)
  );
  OptimizationBarrier entries_barrier_6 ( // @[package.scala 258:25]
    .io_x_ppn(entries_barrier_6_io_x_ppn),
    .io_x_u(entries_barrier_6_io_x_u),
    .io_x_ae(entries_barrier_6_io_x_ae),
    .io_x_sw(entries_barrier_6_io_x_sw),
    .io_x_sx(entries_barrier_6_io_x_sx),
    .io_x_sr(entries_barrier_6_io_x_sr),
    .io_x_pw(entries_barrier_6_io_x_pw),
    .io_x_px(entries_barrier_6_io_x_px),
    .io_x_pr(entries_barrier_6_io_x_pr),
    .io_x_ppp(entries_barrier_6_io_x_ppp),
    .io_x_pal(entries_barrier_6_io_x_pal),
    .io_x_paa(entries_barrier_6_io_x_paa),
    .io_x_eff(entries_barrier_6_io_x_eff),
    .io_x_c(entries_barrier_6_io_x_c),
    .io_y_ppn(entries_barrier_6_io_y_ppn),
    .io_y_u(entries_barrier_6_io_y_u),
    .io_y_ae(entries_barrier_6_io_y_ae),
    .io_y_sw(entries_barrier_6_io_y_sw),
    .io_y_sx(entries_barrier_6_io_y_sx),
    .io_y_sr(entries_barrier_6_io_y_sr),
    .io_y_pw(entries_barrier_6_io_y_pw),
    .io_y_px(entries_barrier_6_io_y_px),
    .io_y_pr(entries_barrier_6_io_y_pr),
    .io_y_ppp(entries_barrier_6_io_y_ppp),
    .io_y_pal(entries_barrier_6_io_y_pal),
    .io_y_paa(entries_barrier_6_io_y_paa),
    .io_y_eff(entries_barrier_6_io_y_eff),
    .io_y_c(entries_barrier_6_io_y_c),
    .io_covSum(entries_barrier_6_io_covSum),
    .metaAssert(entries_barrier_6_metaAssert)
  );
  OptimizationBarrier entries_barrier_7 ( // @[package.scala 258:25]
    .io_x_ppn(entries_barrier_7_io_x_ppn),
    .io_x_u(entries_barrier_7_io_x_u),
    .io_x_ae(entries_barrier_7_io_x_ae),
    .io_x_sw(entries_barrier_7_io_x_sw),
    .io_x_sx(entries_barrier_7_io_x_sx),
    .io_x_sr(entries_barrier_7_io_x_sr),
    .io_x_pw(entries_barrier_7_io_x_pw),
    .io_x_px(entries_barrier_7_io_x_px),
    .io_x_pr(entries_barrier_7_io_x_pr),
    .io_x_ppp(entries_barrier_7_io_x_ppp),
    .io_x_pal(entries_barrier_7_io_x_pal),
    .io_x_paa(entries_barrier_7_io_x_paa),
    .io_x_eff(entries_barrier_7_io_x_eff),
    .io_x_c(entries_barrier_7_io_x_c),
    .io_y_ppn(entries_barrier_7_io_y_ppn),
    .io_y_u(entries_barrier_7_io_y_u),
    .io_y_ae(entries_barrier_7_io_y_ae),
    .io_y_sw(entries_barrier_7_io_y_sw),
    .io_y_sx(entries_barrier_7_io_y_sx),
    .io_y_sr(entries_barrier_7_io_y_sr),
    .io_y_pw(entries_barrier_7_io_y_pw),
    .io_y_px(entries_barrier_7_io_y_px),
    .io_y_pr(entries_barrier_7_io_y_pr),
    .io_y_ppp(entries_barrier_7_io_y_ppp),
    .io_y_pal(entries_barrier_7_io_y_pal),
    .io_y_paa(entries_barrier_7_io_y_paa),
    .io_y_eff(entries_barrier_7_io_y_eff),
    .io_y_c(entries_barrier_7_io_y_c),
    .io_covSum(entries_barrier_7_io_covSum),
    .metaAssert(entries_barrier_7_metaAssert)
  );
  OptimizationBarrier entries_barrier_8 ( // @[package.scala 258:25]
    .io_x_ppn(entries_barrier_8_io_x_ppn),
    .io_x_u(entries_barrier_8_io_x_u),
    .io_x_ae(entries_barrier_8_io_x_ae),
    .io_x_sw(entries_barrier_8_io_x_sw),
    .io_x_sx(entries_barrier_8_io_x_sx),
    .io_x_sr(entries_barrier_8_io_x_sr),
    .io_x_pw(entries_barrier_8_io_x_pw),
    .io_x_px(entries_barrier_8_io_x_px),
    .io_x_pr(entries_barrier_8_io_x_pr),
    .io_x_ppp(entries_barrier_8_io_x_ppp),
    .io_x_pal(entries_barrier_8_io_x_pal),
    .io_x_paa(entries_barrier_8_io_x_paa),
    .io_x_eff(entries_barrier_8_io_x_eff),
    .io_x_c(entries_barrier_8_io_x_c),
    .io_y_ppn(entries_barrier_8_io_y_ppn),
    .io_y_u(entries_barrier_8_io_y_u),
    .io_y_ae(entries_barrier_8_io_y_ae),
    .io_y_sw(entries_barrier_8_io_y_sw),
    .io_y_sx(entries_barrier_8_io_y_sx),
    .io_y_sr(entries_barrier_8_io_y_sr),
    .io_y_pw(entries_barrier_8_io_y_pw),
    .io_y_px(entries_barrier_8_io_y_px),
    .io_y_pr(entries_barrier_8_io_y_pr),
    .io_y_ppp(entries_barrier_8_io_y_ppp),
    .io_y_pal(entries_barrier_8_io_y_pal),
    .io_y_paa(entries_barrier_8_io_y_paa),
    .io_y_eff(entries_barrier_8_io_y_eff),
    .io_y_c(entries_barrier_8_io_y_c),
    .io_covSum(entries_barrier_8_io_covSum),
    .metaAssert(entries_barrier_8_metaAssert)
  );
  OptimizationBarrier entries_barrier_9 ( // @[package.scala 258:25]
    .io_x_ppn(entries_barrier_9_io_x_ppn),
    .io_x_u(entries_barrier_9_io_x_u),
    .io_x_ae(entries_barrier_9_io_x_ae),
    .io_x_sw(entries_barrier_9_io_x_sw),
    .io_x_sx(entries_barrier_9_io_x_sx),
    .io_x_sr(entries_barrier_9_io_x_sr),
    .io_x_pw(entries_barrier_9_io_x_pw),
    .io_x_px(entries_barrier_9_io_x_px),
    .io_x_pr(entries_barrier_9_io_x_pr),
    .io_x_ppp(entries_barrier_9_io_x_ppp),
    .io_x_pal(entries_barrier_9_io_x_pal),
    .io_x_paa(entries_barrier_9_io_x_paa),
    .io_x_eff(entries_barrier_9_io_x_eff),
    .io_x_c(entries_barrier_9_io_x_c),
    .io_y_ppn(entries_barrier_9_io_y_ppn),
    .io_y_u(entries_barrier_9_io_y_u),
    .io_y_ae(entries_barrier_9_io_y_ae),
    .io_y_sw(entries_barrier_9_io_y_sw),
    .io_y_sx(entries_barrier_9_io_y_sx),
    .io_y_sr(entries_barrier_9_io_y_sr),
    .io_y_pw(entries_barrier_9_io_y_pw),
    .io_y_px(entries_barrier_9_io_y_px),
    .io_y_pr(entries_barrier_9_io_y_pr),
    .io_y_ppp(entries_barrier_9_io_y_ppp),
    .io_y_pal(entries_barrier_9_io_y_pal),
    .io_y_paa(entries_barrier_9_io_y_paa),
    .io_y_eff(entries_barrier_9_io_y_eff),
    .io_y_c(entries_barrier_9_io_y_c),
    .io_covSum(entries_barrier_9_io_covSum),
    .metaAssert(entries_barrier_9_metaAssert)
  );
  OptimizationBarrier entries_barrier_10 ( // @[package.scala 258:25]
    .io_x_ppn(entries_barrier_10_io_x_ppn),
    .io_x_u(entries_barrier_10_io_x_u),
    .io_x_ae(entries_barrier_10_io_x_ae),
    .io_x_sw(entries_barrier_10_io_x_sw),
    .io_x_sx(entries_barrier_10_io_x_sx),
    .io_x_sr(entries_barrier_10_io_x_sr),
    .io_x_pw(entries_barrier_10_io_x_pw),
    .io_x_px(entries_barrier_10_io_x_px),
    .io_x_pr(entries_barrier_10_io_x_pr),
    .io_x_ppp(entries_barrier_10_io_x_ppp),
    .io_x_pal(entries_barrier_10_io_x_pal),
    .io_x_paa(entries_barrier_10_io_x_paa),
    .io_x_eff(entries_barrier_10_io_x_eff),
    .io_x_c(entries_barrier_10_io_x_c),
    .io_y_ppn(entries_barrier_10_io_y_ppn),
    .io_y_u(entries_barrier_10_io_y_u),
    .io_y_ae(entries_barrier_10_io_y_ae),
    .io_y_sw(entries_barrier_10_io_y_sw),
    .io_y_sx(entries_barrier_10_io_y_sx),
    .io_y_sr(entries_barrier_10_io_y_sr),
    .io_y_pw(entries_barrier_10_io_y_pw),
    .io_y_px(entries_barrier_10_io_y_px),
    .io_y_pr(entries_barrier_10_io_y_pr),
    .io_y_ppp(entries_barrier_10_io_y_ppp),
    .io_y_pal(entries_barrier_10_io_y_pal),
    .io_y_paa(entries_barrier_10_io_y_paa),
    .io_y_eff(entries_barrier_10_io_y_eff),
    .io_y_c(entries_barrier_10_io_y_c),
    .io_covSum(entries_barrier_10_io_covSum),
    .metaAssert(entries_barrier_10_metaAssert)
  );
  OptimizationBarrier entries_barrier_11 ( // @[package.scala 258:25]
    .io_x_ppn(entries_barrier_11_io_x_ppn),
    .io_x_u(entries_barrier_11_io_x_u),
    .io_x_ae(entries_barrier_11_io_x_ae),
    .io_x_sw(entries_barrier_11_io_x_sw),
    .io_x_sx(entries_barrier_11_io_x_sx),
    .io_x_sr(entries_barrier_11_io_x_sr),
    .io_x_pw(entries_barrier_11_io_x_pw),
    .io_x_px(entries_barrier_11_io_x_px),
    .io_x_pr(entries_barrier_11_io_x_pr),
    .io_x_ppp(entries_barrier_11_io_x_ppp),
    .io_x_pal(entries_barrier_11_io_x_pal),
    .io_x_paa(entries_barrier_11_io_x_paa),
    .io_x_eff(entries_barrier_11_io_x_eff),
    .io_x_c(entries_barrier_11_io_x_c),
    .io_y_ppn(entries_barrier_11_io_y_ppn),
    .io_y_u(entries_barrier_11_io_y_u),
    .io_y_ae(entries_barrier_11_io_y_ae),
    .io_y_sw(entries_barrier_11_io_y_sw),
    .io_y_sx(entries_barrier_11_io_y_sx),
    .io_y_sr(entries_barrier_11_io_y_sr),
    .io_y_pw(entries_barrier_11_io_y_pw),
    .io_y_px(entries_barrier_11_io_y_px),
    .io_y_pr(entries_barrier_11_io_y_pr),
    .io_y_ppp(entries_barrier_11_io_y_ppp),
    .io_y_pal(entries_barrier_11_io_y_pal),
    .io_y_paa(entries_barrier_11_io_y_paa),
    .io_y_eff(entries_barrier_11_io_y_eff),
    .io_y_c(entries_barrier_11_io_y_c),
    .io_covSum(entries_barrier_11_io_covSum),
    .metaAssert(entries_barrier_11_metaAssert)
  );
  OptimizationBarrier entries_barrier_12 ( // @[package.scala 258:25]
    .io_x_ppn(entries_barrier_12_io_x_ppn),
    .io_x_u(entries_barrier_12_io_x_u),
    .io_x_ae(entries_barrier_12_io_x_ae),
    .io_x_sw(entries_barrier_12_io_x_sw),
    .io_x_sx(entries_barrier_12_io_x_sx),
    .io_x_sr(entries_barrier_12_io_x_sr),
    .io_x_pw(entries_barrier_12_io_x_pw),
    .io_x_px(entries_barrier_12_io_x_px),
    .io_x_pr(entries_barrier_12_io_x_pr),
    .io_x_ppp(entries_barrier_12_io_x_ppp),
    .io_x_pal(entries_barrier_12_io_x_pal),
    .io_x_paa(entries_barrier_12_io_x_paa),
    .io_x_eff(entries_barrier_12_io_x_eff),
    .io_x_c(entries_barrier_12_io_x_c),
    .io_y_ppn(entries_barrier_12_io_y_ppn),
    .io_y_u(entries_barrier_12_io_y_u),
    .io_y_ae(entries_barrier_12_io_y_ae),
    .io_y_sw(entries_barrier_12_io_y_sw),
    .io_y_sx(entries_barrier_12_io_y_sx),
    .io_y_sr(entries_barrier_12_io_y_sr),
    .io_y_pw(entries_barrier_12_io_y_pw),
    .io_y_px(entries_barrier_12_io_y_px),
    .io_y_pr(entries_barrier_12_io_y_pr),
    .io_y_ppp(entries_barrier_12_io_y_ppp),
    .io_y_pal(entries_barrier_12_io_y_pal),
    .io_y_paa(entries_barrier_12_io_y_paa),
    .io_y_eff(entries_barrier_12_io_y_eff),
    .io_y_c(entries_barrier_12_io_y_c),
    .io_covSum(entries_barrier_12_io_covSum),
    .metaAssert(entries_barrier_12_metaAssert)
  );
  assign vpn = io_req_bits_vaddr[38:12]; // @[TLB.scala 162:30]
  assign priv_s = io_ptw_status_prv[0]; // @[TLB.scala 180:20]
  assign priv_uses_vm = io_ptw_status_prv <= 2'h1; // @[TLB.scala 181:27]
  assign vm_enabled = io_ptw_ptbr_mode[3] & priv_uses_vm; // @[TLB.scala 182:83]
  assign refill_ppn = io_ptw_resp_bits_pte_ppn[19:0]; // @[TLB.scala 185:44]
  assign _invalidate_refill_T = state == 2'h1; // @[package.scala 15:47]
  assign _invalidate_refill_T_1 = state == 2'h3; // @[package.scala 15:47]
  assign _invalidate_refill_T_2 = _invalidate_refill_T | _invalidate_refill_T_1; // @[package.scala 72:59]
  assign invalidate_refill = _invalidate_refill_T_2 | io_sfence_valid; // @[TLB.scala 187:88]
  assign mpu_ppn_hi = mpu_ppn_barrier_io_y_ppn[19:18]; // @[TLB.scala 105:26]
  assign mpu_ppn_ignore = special_entry_level < 2'h1; // @[TLB.scala 107:28]
  assign _mpu_ppn_T_17 = mpu_ppn_ignore ? vpn : 27'h0; // @[TLB.scala 108:28]
  assign _GEN_919 = {{7'd0}, mpu_ppn_barrier_io_y_ppn}; // @[TLB.scala 108:47]
  assign _mpu_ppn_T_18 = _mpu_ppn_T_17 | _GEN_919; // @[TLB.scala 108:47]
  assign mpu_ppn_lo = _mpu_ppn_T_18[17:9]; // @[TLB.scala 108:58]
  assign mpu_ppn_ignore_1 = special_entry_level < 2'h2; // @[TLB.scala 107:28]
  assign _mpu_ppn_T_19 = mpu_ppn_ignore_1 ? vpn : 27'h0; // @[TLB.scala 108:28]
  assign _mpu_ppn_T_20 = _mpu_ppn_T_19 | _GEN_919; // @[TLB.scala 108:47]
  assign mpu_ppn_lo_1 = _mpu_ppn_T_20[8:0]; // @[TLB.scala 108:58]
  assign _mpu_ppn_T_21 = {mpu_ppn_hi,mpu_ppn_lo,mpu_ppn_lo_1}; // @[Cat.scala 30:58]
  assign _mpu_ppn_T_23 = vm_enabled ? {{8'd0}, _mpu_ppn_T_21} : io_req_bits_vaddr[39:12]; // @[TLB.scala 189:20]
  assign mpu_ppn = io_ptw_resp_valid ? {{8'd0}, refill_ppn} : _mpu_ppn_T_23; // @[TLB.scala 188:20]
  assign mpu_physaddr_lo = io_req_bits_vaddr[11:0]; // @[TLB.scala 190:52]
  assign mpu_physaddr = {mpu_ppn,mpu_physaddr_lo}; // @[Cat.scala 30:58]
  assign _mpu_priv_T_2 = {io_ptw_status_debug,io_ptw_status_prv}; // @[Cat.scala 30:58]
  assign mpu_priv = io_ptw_resp_valid ? 3'h1 : _mpu_priv_T_2; // @[TLB.scala 191:27]
  assign _legal_address_T = mpu_physaddr ^ 40'h3000; // @[Parameters.scala 137:31]
  assign _legal_address_T_1 = {1'b0,$signed(_legal_address_T)}; // @[Parameters.scala 137:49]
  assign _legal_address_T_3 = $signed(_legal_address_T_1) & -41'sh1000; // @[Parameters.scala 137:52]
  assign _legal_address_T_4 = $signed(_legal_address_T_3) == 41'sh0; // @[Parameters.scala 137:67]
  assign _legal_address_T_5 = mpu_physaddr ^ 40'hc000000; // @[Parameters.scala 137:31]
  assign _legal_address_T_6 = {1'b0,$signed(_legal_address_T_5)}; // @[Parameters.scala 137:49]
  assign _legal_address_T_8 = $signed(_legal_address_T_6) & -41'sh4000000; // @[Parameters.scala 137:52]
  assign _legal_address_T_9 = $signed(_legal_address_T_8) == 41'sh0; // @[Parameters.scala 137:67]
  assign _legal_address_T_10 = mpu_physaddr ^ 40'h2000000; // @[Parameters.scala 137:31]
  assign _legal_address_T_11 = {1'b0,$signed(_legal_address_T_10)}; // @[Parameters.scala 137:49]
  assign _legal_address_T_13 = $signed(_legal_address_T_11) & -41'sh10000; // @[Parameters.scala 137:52]
  assign _legal_address_T_14 = $signed(_legal_address_T_13) == 41'sh0; // @[Parameters.scala 137:67]
  assign _legal_address_T_16 = {1'b0,$signed(mpu_physaddr)}; // @[Parameters.scala 137:49]
  assign _legal_address_T_18 = $signed(_legal_address_T_16) & -41'sh1000; // @[Parameters.scala 137:52]
  assign _legal_address_T_19 = $signed(_legal_address_T_18) == 41'sh0; // @[Parameters.scala 137:67]
  assign _legal_address_T_20 = mpu_physaddr ^ 40'h10000; // @[Parameters.scala 137:31]
  assign _legal_address_T_21 = {1'b0,$signed(_legal_address_T_20)}; // @[Parameters.scala 137:49]
  assign _legal_address_T_23 = $signed(_legal_address_T_21) & -41'sh10000; // @[Parameters.scala 137:52]
  assign _legal_address_T_24 = $signed(_legal_address_T_23) == 41'sh0; // @[Parameters.scala 137:67]
  assign _legal_address_T_25 = mpu_physaddr ^ 40'h80000000; // @[Parameters.scala 137:31]
  assign _legal_address_T_26 = {1'b0,$signed(_legal_address_T_25)}; // @[Parameters.scala 137:49]
  assign _legal_address_T_28 = $signed(_legal_address_T_26) & -41'sh10000000; // @[Parameters.scala 137:52]
  assign _legal_address_T_29 = $signed(_legal_address_T_28) == 41'sh0; // @[Parameters.scala 137:67]
  assign _legal_address_T_30 = mpu_physaddr ^ 40'h60000000; // @[Parameters.scala 137:31]
  assign _legal_address_T_31 = {1'b0,$signed(_legal_address_T_30)}; // @[Parameters.scala 137:49]
  assign _legal_address_T_33 = $signed(_legal_address_T_31) & -41'sh20000000; // @[Parameters.scala 137:52]
  assign _legal_address_T_34 = $signed(_legal_address_T_33) == 41'sh0; // @[Parameters.scala 137:67]
  assign _legal_address_T_35 = _legal_address_T_4 | _legal_address_T_9; // @[TLB.scala 197:67]
  assign _legal_address_T_36 = _legal_address_T_35 | _legal_address_T_14; // @[TLB.scala 197:67]
  assign _legal_address_T_37 = _legal_address_T_36 | _legal_address_T_19; // @[TLB.scala 197:67]
  assign _legal_address_T_38 = _legal_address_T_37 | _legal_address_T_24; // @[TLB.scala 197:67]
  assign _legal_address_T_39 = _legal_address_T_38 | _legal_address_T_29; // @[TLB.scala 197:67]
  assign legal_address = _legal_address_T_39 | _legal_address_T_34; // @[TLB.scala 197:67]
  assign _cacheable_T_8 = $signed(_legal_address_T_26) & 41'sh80000000; // @[Parameters.scala 137:52]
  assign _cacheable_T_9 = $signed(_cacheable_T_8) == 41'sh0; // @[Parameters.scala 137:67]
  assign cacheable = legal_address & _cacheable_T_9; // @[TLB.scala 199:19]
  assign _homogeneous_T_54 = mpu_physaddr ^ 40'h8000000; // @[Parameters.scala 137:31]
  assign _homogeneous_T_55 = {1'b0,$signed(_homogeneous_T_54)}; // @[Parameters.scala 137:49]
  assign _homogeneous_T_57 = $signed(_homogeneous_T_55) & 41'shc8000000; // @[Parameters.scala 137:52]
  assign _homogeneous_T_58 = $signed(_homogeneous_T_57) == 41'sh0; // @[Parameters.scala 137:67]
  assign _homogeneous_T_71 = $signed(_legal_address_T_16) & 41'shc8010000; // @[Parameters.scala 137:52]
  assign _homogeneous_T_72 = $signed(_homogeneous_T_71) == 41'sh0; // @[Parameters.scala 137:67]
  assign _homogeneous_T_79 = _homogeneous_T_72 | _homogeneous_T_58; // @[TLBPermissions.scala 83:66]
  assign _deny_access_to_debug_T = mpu_priv <= 3'h3; // @[TLB.scala 202:39]
  assign deny_access_to_debug = _deny_access_to_debug_T & _legal_address_T_19; // @[TLB.scala 202:48]
  assign _prot_r_T_7 = legal_address & ~deny_access_to_debug; // @[TLB.scala 203:41]
  assign prot_r = _prot_r_T_7 & pmp_io_r; // @[TLB.scala 203:66]
  assign _prot_w_T_10 = mpu_physaddr ^ 40'h40000000; // @[Parameters.scala 137:31]
  assign _prot_w_T_11 = {1'b0,$signed(_prot_w_T_10)}; // @[Parameters.scala 137:49]
  assign _prot_w_T_13 = $signed(_prot_w_T_11) & 41'shc0000000; // @[Parameters.scala 137:52]
  assign _prot_w_T_14 = $signed(_prot_w_T_13) == 41'sh0; // @[Parameters.scala 137:67]
  assign _prot_w_T_18 = $signed(_legal_address_T_26) & 41'shc0000000; // @[Parameters.scala 137:52]
  assign _prot_w_T_19 = $signed(_prot_w_T_18) == 41'sh0; // @[Parameters.scala 137:67]
  assign _prot_w_T_21 = _homogeneous_T_79 | _prot_w_T_14; // @[Parameters.scala 615:89]
  assign _prot_w_T_22 = _prot_w_T_21 | _prot_w_T_19; // @[Parameters.scala 615:89]
  assign _prot_w_T_31 = legal_address & _prot_w_T_22; // @[TLB.scala 199:19]
  assign _prot_w_T_33 = _prot_w_T_31 & ~deny_access_to_debug; // @[TLB.scala 204:45]
  assign prot_w = _prot_w_T_33 & pmp_io_w; // @[TLB.scala 204:70]
  assign prot_al = legal_address & _homogeneous_T_79; // @[TLB.scala 199:19]
  assign _prot_x_T_3 = $signed(_legal_address_T_16) & 41'shca000000; // @[Parameters.scala 137:52]
  assign _prot_x_T_4 = $signed(_prot_x_T_3) == 41'sh0; // @[Parameters.scala 137:67]
  assign _prot_x_T_15 = _prot_x_T_4 | _prot_w_T_14; // @[Parameters.scala 615:89]
  assign _prot_x_T_16 = _prot_x_T_15 | _prot_w_T_19; // @[Parameters.scala 615:89]
  assign _prot_x_T_31 = legal_address & _prot_x_T_16; // @[TLB.scala 199:19]
  assign _prot_x_T_33 = _prot_x_T_31 & ~deny_access_to_debug; // @[TLB.scala 208:40]
  assign prot_x = _prot_x_T_33 & pmp_io_x; // @[TLB.scala 208:65]
  assign _prot_eff_T_20 = $signed(_legal_address_T_16) & 41'shca012000; // @[Parameters.scala 137:52]
  assign _prot_eff_T_21 = $signed(_prot_eff_T_20) == 41'sh0; // @[Parameters.scala 137:67]
  assign _prot_eff_T_25 = $signed(_legal_address_T_11) & 41'shca010000; // @[Parameters.scala 137:52]
  assign _prot_eff_T_26 = $signed(_prot_eff_T_25) == 41'sh0; // @[Parameters.scala 137:67]
  assign _prot_eff_T_37 = _prot_eff_T_21 | _prot_eff_T_26; // @[Parameters.scala 615:89]
  assign _prot_eff_T_38 = _prot_eff_T_37 | _homogeneous_T_58; // @[Parameters.scala 615:89]
  assign _prot_eff_T_39 = _prot_eff_T_38 | _prot_w_T_14; // @[Parameters.scala 615:89]
  assign prot_eff = legal_address & _prot_eff_T_39; // @[TLB.scala 199:19]
  assign _sector_hits_T = sectored_entries_0_0_valid_0 | sectored_entries_0_0_valid_1; // @[package.scala 72:59]
  assign _sector_hits_T_1 = _sector_hits_T | sectored_entries_0_0_valid_2; // @[package.scala 72:59]
  assign _sector_hits_T_2 = _sector_hits_T_1 | sectored_entries_0_0_valid_3; // @[package.scala 72:59]
  assign _sector_hits_T_3 = sectored_entries_0_0_tag ^ vpn; // @[TLB.scala 88:41]
  assign _sector_hits_T_5 = _sector_hits_T_3[26:2] == 25'h0; // @[TLB.scala 88:66]
  assign sector_hits_0 = _sector_hits_T_2 & _sector_hits_T_5; // @[TLB.scala 87:40]
  assign _sector_hits_T_6 = sectored_entries_0_1_valid_0 | sectored_entries_0_1_valid_1; // @[package.scala 72:59]
  assign _sector_hits_T_7 = _sector_hits_T_6 | sectored_entries_0_1_valid_2; // @[package.scala 72:59]
  assign _sector_hits_T_8 = _sector_hits_T_7 | sectored_entries_0_1_valid_3; // @[package.scala 72:59]
  assign _sector_hits_T_9 = sectored_entries_0_1_tag ^ vpn; // @[TLB.scala 88:41]
  assign _sector_hits_T_11 = _sector_hits_T_9[26:2] == 25'h0; // @[TLB.scala 88:66]
  assign sector_hits_1 = _sector_hits_T_8 & _sector_hits_T_11; // @[TLB.scala 87:40]
  assign _sector_hits_T_12 = sectored_entries_0_2_valid_0 | sectored_entries_0_2_valid_1; // @[package.scala 72:59]
  assign _sector_hits_T_13 = _sector_hits_T_12 | sectored_entries_0_2_valid_2; // @[package.scala 72:59]
  assign _sector_hits_T_14 = _sector_hits_T_13 | sectored_entries_0_2_valid_3; // @[package.scala 72:59]
  assign _sector_hits_T_15 = sectored_entries_0_2_tag ^ vpn; // @[TLB.scala 88:41]
  assign _sector_hits_T_17 = _sector_hits_T_15[26:2] == 25'h0; // @[TLB.scala 88:66]
  assign sector_hits_2 = _sector_hits_T_14 & _sector_hits_T_17; // @[TLB.scala 87:40]
  assign _sector_hits_T_18 = sectored_entries_0_3_valid_0 | sectored_entries_0_3_valid_1; // @[package.scala 72:59]
  assign _sector_hits_T_19 = _sector_hits_T_18 | sectored_entries_0_3_valid_2; // @[package.scala 72:59]
  assign _sector_hits_T_20 = _sector_hits_T_19 | sectored_entries_0_3_valid_3; // @[package.scala 72:59]
  assign _sector_hits_T_21 = sectored_entries_0_3_tag ^ vpn; // @[TLB.scala 88:41]
  assign _sector_hits_T_23 = _sector_hits_T_21[26:2] == 25'h0; // @[TLB.scala 88:66]
  assign sector_hits_3 = _sector_hits_T_20 & _sector_hits_T_23; // @[TLB.scala 87:40]
  assign _sector_hits_T_24 = sectored_entries_0_4_valid_0 | sectored_entries_0_4_valid_1; // @[package.scala 72:59]
  assign _sector_hits_T_25 = _sector_hits_T_24 | sectored_entries_0_4_valid_2; // @[package.scala 72:59]
  assign _sector_hits_T_26 = _sector_hits_T_25 | sectored_entries_0_4_valid_3; // @[package.scala 72:59]
  assign _sector_hits_T_27 = sectored_entries_0_4_tag ^ vpn; // @[TLB.scala 88:41]
  assign _sector_hits_T_29 = _sector_hits_T_27[26:2] == 25'h0; // @[TLB.scala 88:66]
  assign sector_hits_4 = _sector_hits_T_26 & _sector_hits_T_29; // @[TLB.scala 87:40]
  assign _sector_hits_T_30 = sectored_entries_0_5_valid_0 | sectored_entries_0_5_valid_1; // @[package.scala 72:59]
  assign _sector_hits_T_31 = _sector_hits_T_30 | sectored_entries_0_5_valid_2; // @[package.scala 72:59]
  assign _sector_hits_T_32 = _sector_hits_T_31 | sectored_entries_0_5_valid_3; // @[package.scala 72:59]
  assign _sector_hits_T_33 = sectored_entries_0_5_tag ^ vpn; // @[TLB.scala 88:41]
  assign _sector_hits_T_35 = _sector_hits_T_33[26:2] == 25'h0; // @[TLB.scala 88:66]
  assign sector_hits_5 = _sector_hits_T_32 & _sector_hits_T_35; // @[TLB.scala 87:40]
  assign _sector_hits_T_36 = sectored_entries_0_6_valid_0 | sectored_entries_0_6_valid_1; // @[package.scala 72:59]
  assign _sector_hits_T_37 = _sector_hits_T_36 | sectored_entries_0_6_valid_2; // @[package.scala 72:59]
  assign _sector_hits_T_38 = _sector_hits_T_37 | sectored_entries_0_6_valid_3; // @[package.scala 72:59]
  assign _sector_hits_T_39 = sectored_entries_0_6_tag ^ vpn; // @[TLB.scala 88:41]
  assign _sector_hits_T_41 = _sector_hits_T_39[26:2] == 25'h0; // @[TLB.scala 88:66]
  assign sector_hits_6 = _sector_hits_T_38 & _sector_hits_T_41; // @[TLB.scala 87:40]
  assign _sector_hits_T_42 = sectored_entries_0_7_valid_0 | sectored_entries_0_7_valid_1; // @[package.scala 72:59]
  assign _sector_hits_T_43 = _sector_hits_T_42 | sectored_entries_0_7_valid_2; // @[package.scala 72:59]
  assign _sector_hits_T_44 = _sector_hits_T_43 | sectored_entries_0_7_valid_3; // @[package.scala 72:59]
  assign _sector_hits_T_45 = sectored_entries_0_7_tag ^ vpn; // @[TLB.scala 88:41]
  assign _sector_hits_T_47 = _sector_hits_T_45[26:2] == 25'h0; // @[TLB.scala 88:66]
  assign sector_hits_7 = _sector_hits_T_44 & _sector_hits_T_47; // @[TLB.scala 87:40]
  assign _superpage_hits_T_2 = superpage_entries_0_tag[26:18] == vpn[26:18]; // @[TLB.scala 95:77]
  assign _superpage_hits_T_4 = superpage_entries_0_valid_0 & _superpage_hits_T_2; // @[TLB.scala 95:29]
  assign superpage_hits_ignore_1 = superpage_entries_0_level < 2'h1; // @[TLB.scala 94:28]
  assign _superpage_hits_T_7 = superpage_entries_0_tag[17:9] == vpn[17:9]; // @[TLB.scala 95:77]
  assign _superpage_hits_T_8 = superpage_hits_ignore_1 | _superpage_hits_T_7; // @[TLB.scala 95:40]
  assign superpage_hits_0 = _superpage_hits_T_4 & _superpage_hits_T_8; // @[TLB.scala 95:29]
  assign _superpage_hits_T_16 = superpage_entries_1_tag[26:18] == vpn[26:18]; // @[TLB.scala 95:77]
  assign _superpage_hits_T_18 = superpage_entries_1_valid_0 & _superpage_hits_T_16; // @[TLB.scala 95:29]
  assign superpage_hits_ignore_4 = superpage_entries_1_level < 2'h1; // @[TLB.scala 94:28]
  assign _superpage_hits_T_21 = superpage_entries_1_tag[17:9] == vpn[17:9]; // @[TLB.scala 95:77]
  assign _superpage_hits_T_22 = superpage_hits_ignore_4 | _superpage_hits_T_21; // @[TLB.scala 95:40]
  assign superpage_hits_1 = _superpage_hits_T_18 & _superpage_hits_T_22; // @[TLB.scala 95:29]
  assign _superpage_hits_T_30 = superpage_entries_2_tag[26:18] == vpn[26:18]; // @[TLB.scala 95:77]
  assign _superpage_hits_T_32 = superpage_entries_2_valid_0 & _superpage_hits_T_30; // @[TLB.scala 95:29]
  assign superpage_hits_ignore_7 = superpage_entries_2_level < 2'h1; // @[TLB.scala 94:28]
  assign _superpage_hits_T_35 = superpage_entries_2_tag[17:9] == vpn[17:9]; // @[TLB.scala 95:77]
  assign _superpage_hits_T_36 = superpage_hits_ignore_7 | _superpage_hits_T_35; // @[TLB.scala 95:40]
  assign superpage_hits_2 = _superpage_hits_T_32 & _superpage_hits_T_36; // @[TLB.scala 95:29]
  assign _superpage_hits_T_44 = superpage_entries_3_tag[26:18] == vpn[26:18]; // @[TLB.scala 95:77]
  assign _superpage_hits_T_46 = superpage_entries_3_valid_0 & _superpage_hits_T_44; // @[TLB.scala 95:29]
  assign superpage_hits_ignore_10 = superpage_entries_3_level < 2'h1; // @[TLB.scala 94:28]
  assign _superpage_hits_T_49 = superpage_entries_3_tag[17:9] == vpn[17:9]; // @[TLB.scala 95:77]
  assign _superpage_hits_T_50 = superpage_hits_ignore_10 | _superpage_hits_T_49; // @[TLB.scala 95:40]
  assign superpage_hits_3 = _superpage_hits_T_46 & _superpage_hits_T_50; // @[TLB.scala 95:29]
  assign hitsVec_idx = vpn[1:0]; // @[package.scala 154:13]
  assign _GEN_1 = 2'h1 == hitsVec_idx ? sectored_entries_0_0_valid_1 : sectored_entries_0_0_valid_0; // @[TLB.scala 100:18]
  assign _GEN_2 = 2'h2 == hitsVec_idx ? sectored_entries_0_0_valid_2 : _GEN_1; // @[TLB.scala 100:18]
  assign _GEN_3 = 2'h3 == hitsVec_idx ? sectored_entries_0_0_valid_3 : _GEN_2; // @[TLB.scala 100:18]
  assign _hitsVec_T_3 = _GEN_3 & _sector_hits_T_5; // @[TLB.scala 100:18]
  assign hitsVec_0 = vm_enabled & _hitsVec_T_3; // @[TLB.scala 213:44]
  assign _GEN_5 = 2'h1 == hitsVec_idx ? sectored_entries_0_1_valid_1 : sectored_entries_0_1_valid_0; // @[TLB.scala 100:18]
  assign _GEN_6 = 2'h2 == hitsVec_idx ? sectored_entries_0_1_valid_2 : _GEN_5; // @[TLB.scala 100:18]
  assign _GEN_7 = 2'h3 == hitsVec_idx ? sectored_entries_0_1_valid_3 : _GEN_6; // @[TLB.scala 100:18]
  assign _hitsVec_T_7 = _GEN_7 & _sector_hits_T_11; // @[TLB.scala 100:18]
  assign hitsVec_1 = vm_enabled & _hitsVec_T_7; // @[TLB.scala 213:44]
  assign _GEN_9 = 2'h1 == hitsVec_idx ? sectored_entries_0_2_valid_1 : sectored_entries_0_2_valid_0; // @[TLB.scala 100:18]
  assign _GEN_10 = 2'h2 == hitsVec_idx ? sectored_entries_0_2_valid_2 : _GEN_9; // @[TLB.scala 100:18]
  assign _GEN_11 = 2'h3 == hitsVec_idx ? sectored_entries_0_2_valid_3 : _GEN_10; // @[TLB.scala 100:18]
  assign _hitsVec_T_11 = _GEN_11 & _sector_hits_T_17; // @[TLB.scala 100:18]
  assign hitsVec_2 = vm_enabled & _hitsVec_T_11; // @[TLB.scala 213:44]
  assign _GEN_13 = 2'h1 == hitsVec_idx ? sectored_entries_0_3_valid_1 : sectored_entries_0_3_valid_0; // @[TLB.scala 100:18]
  assign _GEN_14 = 2'h2 == hitsVec_idx ? sectored_entries_0_3_valid_2 : _GEN_13; // @[TLB.scala 100:18]
  assign _GEN_15 = 2'h3 == hitsVec_idx ? sectored_entries_0_3_valid_3 : _GEN_14; // @[TLB.scala 100:18]
  assign _hitsVec_T_15 = _GEN_15 & _sector_hits_T_23; // @[TLB.scala 100:18]
  assign hitsVec_3 = vm_enabled & _hitsVec_T_15; // @[TLB.scala 213:44]
  assign _GEN_17 = 2'h1 == hitsVec_idx ? sectored_entries_0_4_valid_1 : sectored_entries_0_4_valid_0; // @[TLB.scala 100:18]
  assign _GEN_18 = 2'h2 == hitsVec_idx ? sectored_entries_0_4_valid_2 : _GEN_17; // @[TLB.scala 100:18]
  assign _GEN_19 = 2'h3 == hitsVec_idx ? sectored_entries_0_4_valid_3 : _GEN_18; // @[TLB.scala 100:18]
  assign _hitsVec_T_19 = _GEN_19 & _sector_hits_T_29; // @[TLB.scala 100:18]
  assign hitsVec_4 = vm_enabled & _hitsVec_T_19; // @[TLB.scala 213:44]
  assign _GEN_21 = 2'h1 == hitsVec_idx ? sectored_entries_0_5_valid_1 : sectored_entries_0_5_valid_0; // @[TLB.scala 100:18]
  assign _GEN_22 = 2'h2 == hitsVec_idx ? sectored_entries_0_5_valid_2 : _GEN_21; // @[TLB.scala 100:18]
  assign _GEN_23 = 2'h3 == hitsVec_idx ? sectored_entries_0_5_valid_3 : _GEN_22; // @[TLB.scala 100:18]
  assign _hitsVec_T_23 = _GEN_23 & _sector_hits_T_35; // @[TLB.scala 100:18]
  assign hitsVec_5 = vm_enabled & _hitsVec_T_23; // @[TLB.scala 213:44]
  assign _GEN_25 = 2'h1 == hitsVec_idx ? sectored_entries_0_6_valid_1 : sectored_entries_0_6_valid_0; // @[TLB.scala 100:18]
  assign _GEN_26 = 2'h2 == hitsVec_idx ? sectored_entries_0_6_valid_2 : _GEN_25; // @[TLB.scala 100:18]
  assign _GEN_27 = 2'h3 == hitsVec_idx ? sectored_entries_0_6_valid_3 : _GEN_26; // @[TLB.scala 100:18]
  assign _hitsVec_T_27 = _GEN_27 & _sector_hits_T_41; // @[TLB.scala 100:18]
  assign hitsVec_6 = vm_enabled & _hitsVec_T_27; // @[TLB.scala 213:44]
  assign _GEN_29 = 2'h1 == hitsVec_idx ? sectored_entries_0_7_valid_1 : sectored_entries_0_7_valid_0; // @[TLB.scala 100:18]
  assign _GEN_30 = 2'h2 == hitsVec_idx ? sectored_entries_0_7_valid_2 : _GEN_29; // @[TLB.scala 100:18]
  assign _GEN_31 = 2'h3 == hitsVec_idx ? sectored_entries_0_7_valid_3 : _GEN_30; // @[TLB.scala 100:18]
  assign _hitsVec_T_31 = _GEN_31 & _sector_hits_T_47; // @[TLB.scala 100:18]
  assign hitsVec_7 = vm_enabled & _hitsVec_T_31; // @[TLB.scala 213:44]
  assign hitsVec_8 = vm_enabled & superpage_hits_0; // @[TLB.scala 213:44]
  assign hitsVec_9 = vm_enabled & superpage_hits_1; // @[TLB.scala 213:44]
  assign hitsVec_10 = vm_enabled & superpage_hits_2; // @[TLB.scala 213:44]
  assign hitsVec_11 = vm_enabled & superpage_hits_3; // @[TLB.scala 213:44]
  assign _hitsVec_T_94 = special_entry_tag[26:18] == vpn[26:18]; // @[TLB.scala 95:77]
  assign _hitsVec_T_96 = special_entry_valid_0 & _hitsVec_T_94; // @[TLB.scala 95:29]
  assign _hitsVec_T_99 = special_entry_tag[17:9] == vpn[17:9]; // @[TLB.scala 95:77]
  assign _hitsVec_T_100 = mpu_ppn_ignore | _hitsVec_T_99; // @[TLB.scala 95:40]
  assign _hitsVec_T_101 = _hitsVec_T_96 & _hitsVec_T_100; // @[TLB.scala 95:29]
  assign _hitsVec_T_104 = special_entry_tag[8:0] == vpn[8:0]; // @[TLB.scala 95:77]
  assign _hitsVec_T_105 = mpu_ppn_ignore_1 | _hitsVec_T_104; // @[TLB.scala 95:40]
  assign _hitsVec_T_106 = _hitsVec_T_101 & _hitsVec_T_105; // @[TLB.scala 95:29]
  assign hitsVec_12 = vm_enabled & _hitsVec_T_106; // @[TLB.scala 213:44]
  assign real_hits_lo = {hitsVec_5,hitsVec_4,hitsVec_3,hitsVec_2,hitsVec_1,hitsVec_0}; // @[Cat.scala 30:58]
  assign real_hits = {hitsVec_12,hitsVec_11,hitsVec_10,hitsVec_9,hitsVec_8,hitsVec_7,hitsVec_6,real_hits_lo}; // @[Cat.scala 30:58]
  assign hits_hi = ~vm_enabled; // @[TLB.scala 215:18]
  assign hits = {hits_hi,hitsVec_12,hitsVec_11,hitsVec_10,hitsVec_9,hitsVec_8,hitsVec_7,hitsVec_6,real_hits_lo}; // @[Cat.scala 30:58]
  assign newEntry_g = io_ptw_resp_bits_pte_g & io_ptw_resp_bits_pte_v; // @[TLB.scala 224:25]
  assign _newEntry_sr_T_1 = io_ptw_resp_bits_pte_x & ~io_ptw_resp_bits_pte_w; // @[PTW.scala 73:44]
  assign _newEntry_sr_T_2 = io_ptw_resp_bits_pte_r | _newEntry_sr_T_1; // @[PTW.scala 73:38]
  assign _newEntry_sr_T_3 = io_ptw_resp_bits_pte_v & _newEntry_sr_T_2; // @[PTW.scala 73:32]
  assign _newEntry_sr_T_4 = _newEntry_sr_T_3 & io_ptw_resp_bits_pte_a; // @[PTW.scala 73:52]
  assign newEntry_sr = _newEntry_sr_T_4 & io_ptw_resp_bits_pte_r; // @[PTW.scala 77:35]
  assign _newEntry_sw_T_5 = _newEntry_sr_T_4 & io_ptw_resp_bits_pte_w; // @[PTW.scala 78:35]
  assign newEntry_sw = _newEntry_sw_T_5 & io_ptw_resp_bits_pte_d; // @[PTW.scala 78:40]
  assign newEntry_sx = _newEntry_sr_T_4 & io_ptw_resp_bits_pte_x; // @[PTW.scala 79:35]
  assign special_entry_data_0_lo = {prot_x,prot_r,_prot_w_T_31,prot_al,prot_al,prot_eff,cacheable,1'h0}; // @[TLB.scala 122:24]
  assign _special_entry_data_0_T = {refill_ppn,io_ptw_resp_bits_pte_u,newEntry_g,io_ptw_resp_bits_ae,newEntry_sw,newEntry_sx,newEntry_sr,prot_w,special_entry_data_0_lo}; // @[TLB.scala 122:24]
  assign _GEN_32 = invalidate_refill ? 1'h0 : 1'h1; // @[TLB.scala 241:34]
  assign _T_2 = io_ptw_resp_bits_level < 2'h2; // @[TLB.scala 243:40]
  assign _T_3 = r_superpage_repl_addr == 2'h0; // @[TLB.scala 244:82]
  assign _GEN_35 = _T_3 ? _GEN_32 : superpage_entries_0_valid_0; // @[TLB.scala 244:89]
  assign _T_4 = r_superpage_repl_addr == 2'h1; // @[TLB.scala 244:82]
  assign _GEN_39 = _T_4 ? _GEN_32 : superpage_entries_1_valid_0; // @[TLB.scala 244:89]
  assign _T_5 = r_superpage_repl_addr == 2'h2; // @[TLB.scala 244:82]
  assign _GEN_43 = _T_5 ? _GEN_32 : superpage_entries_2_valid_0; // @[TLB.scala 244:89]
  assign _T_6 = r_superpage_repl_addr == 2'h3; // @[TLB.scala 244:82]
  assign _GEN_47 = _T_6 ? _GEN_32 : superpage_entries_3_valid_0; // @[TLB.scala 244:89]
  assign waddr = r_sectored_hit ? r_sectored_hit_addr : r_sectored_repl_addr; // @[TLB.scala 250:22]
  assign _T_7 = waddr == 3'h0; // @[TLB.scala 251:75]
  assign _GEN_49 = r_sectored_hit ? sectored_entries_0_0_valid_0 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_50 = r_sectored_hit ? sectored_entries_0_0_valid_1 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_51 = r_sectored_hit ? sectored_entries_0_0_valid_2 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_52 = r_sectored_hit ? sectored_entries_0_0_valid_3 : 1'h0; // @[TLB.scala 252:32]
  assign idx = r_refill_tag[1:0]; // @[package.scala 154:13]
  assign _GEN_921 = 2'h0 == idx; // @[TLB.scala 121:16]
  assign _GEN_53 = _GEN_921 | _GEN_49; // @[TLB.scala 121:16]
  assign _GEN_922 = 2'h1 == idx; // @[TLB.scala 121:16]
  assign _GEN_54 = _GEN_922 | _GEN_50; // @[TLB.scala 121:16]
  assign _GEN_923 = 2'h2 == idx; // @[TLB.scala 121:16]
  assign _GEN_55 = _GEN_923 | _GEN_51; // @[TLB.scala 121:16]
  assign _GEN_924 = 2'h3 == idx; // @[TLB.scala 121:16]
  assign _GEN_56 = _GEN_924 | _GEN_52; // @[TLB.scala 121:16]
  assign _GEN_61 = invalidate_refill ? 1'h0 : _GEN_53; // @[TLB.scala 254:34]
  assign _GEN_62 = invalidate_refill ? 1'h0 : _GEN_54; // @[TLB.scala 254:34]
  assign _GEN_63 = invalidate_refill ? 1'h0 : _GEN_55; // @[TLB.scala 254:34]
  assign _GEN_64 = invalidate_refill ? 1'h0 : _GEN_56; // @[TLB.scala 254:34]
  assign _GEN_65 = _T_7 ? _GEN_61 : sectored_entries_0_0_valid_0; // @[TLB.scala 251:82]
  assign _GEN_66 = _T_7 ? _GEN_62 : sectored_entries_0_0_valid_1; // @[TLB.scala 251:82]
  assign _GEN_67 = _T_7 ? _GEN_63 : sectored_entries_0_0_valid_2; // @[TLB.scala 251:82]
  assign _GEN_68 = _T_7 ? _GEN_64 : sectored_entries_0_0_valid_3; // @[TLB.scala 251:82]
  assign _T_9 = waddr == 3'h1; // @[TLB.scala 251:75]
  assign _GEN_75 = r_sectored_hit ? sectored_entries_0_1_valid_0 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_76 = r_sectored_hit ? sectored_entries_0_1_valid_1 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_77 = r_sectored_hit ? sectored_entries_0_1_valid_2 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_78 = r_sectored_hit ? sectored_entries_0_1_valid_3 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_79 = _GEN_921 | _GEN_75; // @[TLB.scala 121:16]
  assign _GEN_80 = _GEN_922 | _GEN_76; // @[TLB.scala 121:16]
  assign _GEN_81 = _GEN_923 | _GEN_77; // @[TLB.scala 121:16]
  assign _GEN_82 = _GEN_924 | _GEN_78; // @[TLB.scala 121:16]
  assign _GEN_87 = invalidate_refill ? 1'h0 : _GEN_79; // @[TLB.scala 254:34]
  assign _GEN_88 = invalidate_refill ? 1'h0 : _GEN_80; // @[TLB.scala 254:34]
  assign _GEN_89 = invalidate_refill ? 1'h0 : _GEN_81; // @[TLB.scala 254:34]
  assign _GEN_90 = invalidate_refill ? 1'h0 : _GEN_82; // @[TLB.scala 254:34]
  assign _GEN_91 = _T_9 ? _GEN_87 : sectored_entries_0_1_valid_0; // @[TLB.scala 251:82]
  assign _GEN_92 = _T_9 ? _GEN_88 : sectored_entries_0_1_valid_1; // @[TLB.scala 251:82]
  assign _GEN_93 = _T_9 ? _GEN_89 : sectored_entries_0_1_valid_2; // @[TLB.scala 251:82]
  assign _GEN_94 = _T_9 ? _GEN_90 : sectored_entries_0_1_valid_3; // @[TLB.scala 251:82]
  assign _T_11 = waddr == 3'h2; // @[TLB.scala 251:75]
  assign _GEN_101 = r_sectored_hit ? sectored_entries_0_2_valid_0 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_102 = r_sectored_hit ? sectored_entries_0_2_valid_1 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_103 = r_sectored_hit ? sectored_entries_0_2_valid_2 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_104 = r_sectored_hit ? sectored_entries_0_2_valid_3 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_105 = _GEN_921 | _GEN_101; // @[TLB.scala 121:16]
  assign _GEN_106 = _GEN_922 | _GEN_102; // @[TLB.scala 121:16]
  assign _GEN_107 = _GEN_923 | _GEN_103; // @[TLB.scala 121:16]
  assign _GEN_108 = _GEN_924 | _GEN_104; // @[TLB.scala 121:16]
  assign _GEN_113 = invalidate_refill ? 1'h0 : _GEN_105; // @[TLB.scala 254:34]
  assign _GEN_114 = invalidate_refill ? 1'h0 : _GEN_106; // @[TLB.scala 254:34]
  assign _GEN_115 = invalidate_refill ? 1'h0 : _GEN_107; // @[TLB.scala 254:34]
  assign _GEN_116 = invalidate_refill ? 1'h0 : _GEN_108; // @[TLB.scala 254:34]
  assign _GEN_117 = _T_11 ? _GEN_113 : sectored_entries_0_2_valid_0; // @[TLB.scala 251:82]
  assign _GEN_118 = _T_11 ? _GEN_114 : sectored_entries_0_2_valid_1; // @[TLB.scala 251:82]
  assign _GEN_119 = _T_11 ? _GEN_115 : sectored_entries_0_2_valid_2; // @[TLB.scala 251:82]
  assign _GEN_120 = _T_11 ? _GEN_116 : sectored_entries_0_2_valid_3; // @[TLB.scala 251:82]
  assign _T_13 = waddr == 3'h3; // @[TLB.scala 251:75]
  assign _GEN_127 = r_sectored_hit ? sectored_entries_0_3_valid_0 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_128 = r_sectored_hit ? sectored_entries_0_3_valid_1 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_129 = r_sectored_hit ? sectored_entries_0_3_valid_2 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_130 = r_sectored_hit ? sectored_entries_0_3_valid_3 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_131 = _GEN_921 | _GEN_127; // @[TLB.scala 121:16]
  assign _GEN_132 = _GEN_922 | _GEN_128; // @[TLB.scala 121:16]
  assign _GEN_133 = _GEN_923 | _GEN_129; // @[TLB.scala 121:16]
  assign _GEN_134 = _GEN_924 | _GEN_130; // @[TLB.scala 121:16]
  assign _GEN_139 = invalidate_refill ? 1'h0 : _GEN_131; // @[TLB.scala 254:34]
  assign _GEN_140 = invalidate_refill ? 1'h0 : _GEN_132; // @[TLB.scala 254:34]
  assign _GEN_141 = invalidate_refill ? 1'h0 : _GEN_133; // @[TLB.scala 254:34]
  assign _GEN_142 = invalidate_refill ? 1'h0 : _GEN_134; // @[TLB.scala 254:34]
  assign _GEN_143 = _T_13 ? _GEN_139 : sectored_entries_0_3_valid_0; // @[TLB.scala 251:82]
  assign _GEN_144 = _T_13 ? _GEN_140 : sectored_entries_0_3_valid_1; // @[TLB.scala 251:82]
  assign _GEN_145 = _T_13 ? _GEN_141 : sectored_entries_0_3_valid_2; // @[TLB.scala 251:82]
  assign _GEN_146 = _T_13 ? _GEN_142 : sectored_entries_0_3_valid_3; // @[TLB.scala 251:82]
  assign _T_15 = waddr == 3'h4; // @[TLB.scala 251:75]
  assign _GEN_153 = r_sectored_hit ? sectored_entries_0_4_valid_0 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_154 = r_sectored_hit ? sectored_entries_0_4_valid_1 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_155 = r_sectored_hit ? sectored_entries_0_4_valid_2 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_156 = r_sectored_hit ? sectored_entries_0_4_valid_3 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_157 = _GEN_921 | _GEN_153; // @[TLB.scala 121:16]
  assign _GEN_158 = _GEN_922 | _GEN_154; // @[TLB.scala 121:16]
  assign _GEN_159 = _GEN_923 | _GEN_155; // @[TLB.scala 121:16]
  assign _GEN_160 = _GEN_924 | _GEN_156; // @[TLB.scala 121:16]
  assign _GEN_165 = invalidate_refill ? 1'h0 : _GEN_157; // @[TLB.scala 254:34]
  assign _GEN_166 = invalidate_refill ? 1'h0 : _GEN_158; // @[TLB.scala 254:34]
  assign _GEN_167 = invalidate_refill ? 1'h0 : _GEN_159; // @[TLB.scala 254:34]
  assign _GEN_168 = invalidate_refill ? 1'h0 : _GEN_160; // @[TLB.scala 254:34]
  assign _GEN_169 = _T_15 ? _GEN_165 : sectored_entries_0_4_valid_0; // @[TLB.scala 251:82]
  assign _GEN_170 = _T_15 ? _GEN_166 : sectored_entries_0_4_valid_1; // @[TLB.scala 251:82]
  assign _GEN_171 = _T_15 ? _GEN_167 : sectored_entries_0_4_valid_2; // @[TLB.scala 251:82]
  assign _GEN_172 = _T_15 ? _GEN_168 : sectored_entries_0_4_valid_3; // @[TLB.scala 251:82]
  assign _T_17 = waddr == 3'h5; // @[TLB.scala 251:75]
  assign _GEN_179 = r_sectored_hit ? sectored_entries_0_5_valid_0 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_180 = r_sectored_hit ? sectored_entries_0_5_valid_1 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_181 = r_sectored_hit ? sectored_entries_0_5_valid_2 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_182 = r_sectored_hit ? sectored_entries_0_5_valid_3 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_183 = _GEN_921 | _GEN_179; // @[TLB.scala 121:16]
  assign _GEN_184 = _GEN_922 | _GEN_180; // @[TLB.scala 121:16]
  assign _GEN_185 = _GEN_923 | _GEN_181; // @[TLB.scala 121:16]
  assign _GEN_186 = _GEN_924 | _GEN_182; // @[TLB.scala 121:16]
  assign _GEN_191 = invalidate_refill ? 1'h0 : _GEN_183; // @[TLB.scala 254:34]
  assign _GEN_192 = invalidate_refill ? 1'h0 : _GEN_184; // @[TLB.scala 254:34]
  assign _GEN_193 = invalidate_refill ? 1'h0 : _GEN_185; // @[TLB.scala 254:34]
  assign _GEN_194 = invalidate_refill ? 1'h0 : _GEN_186; // @[TLB.scala 254:34]
  assign _GEN_195 = _T_17 ? _GEN_191 : sectored_entries_0_5_valid_0; // @[TLB.scala 251:82]
  assign _GEN_196 = _T_17 ? _GEN_192 : sectored_entries_0_5_valid_1; // @[TLB.scala 251:82]
  assign _GEN_197 = _T_17 ? _GEN_193 : sectored_entries_0_5_valid_2; // @[TLB.scala 251:82]
  assign _GEN_198 = _T_17 ? _GEN_194 : sectored_entries_0_5_valid_3; // @[TLB.scala 251:82]
  assign _T_19 = waddr == 3'h6; // @[TLB.scala 251:75]
  assign _GEN_205 = r_sectored_hit ? sectored_entries_0_6_valid_0 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_206 = r_sectored_hit ? sectored_entries_0_6_valid_1 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_207 = r_sectored_hit ? sectored_entries_0_6_valid_2 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_208 = r_sectored_hit ? sectored_entries_0_6_valid_3 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_209 = _GEN_921 | _GEN_205; // @[TLB.scala 121:16]
  assign _GEN_210 = _GEN_922 | _GEN_206; // @[TLB.scala 121:16]
  assign _GEN_211 = _GEN_923 | _GEN_207; // @[TLB.scala 121:16]
  assign _GEN_212 = _GEN_924 | _GEN_208; // @[TLB.scala 121:16]
  assign _GEN_217 = invalidate_refill ? 1'h0 : _GEN_209; // @[TLB.scala 254:34]
  assign _GEN_218 = invalidate_refill ? 1'h0 : _GEN_210; // @[TLB.scala 254:34]
  assign _GEN_219 = invalidate_refill ? 1'h0 : _GEN_211; // @[TLB.scala 254:34]
  assign _GEN_220 = invalidate_refill ? 1'h0 : _GEN_212; // @[TLB.scala 254:34]
  assign _GEN_221 = _T_19 ? _GEN_217 : sectored_entries_0_6_valid_0; // @[TLB.scala 251:82]
  assign _GEN_222 = _T_19 ? _GEN_218 : sectored_entries_0_6_valid_1; // @[TLB.scala 251:82]
  assign _GEN_223 = _T_19 ? _GEN_219 : sectored_entries_0_6_valid_2; // @[TLB.scala 251:82]
  assign _GEN_224 = _T_19 ? _GEN_220 : sectored_entries_0_6_valid_3; // @[TLB.scala 251:82]
  assign _T_21 = waddr == 3'h7; // @[TLB.scala 251:75]
  assign _GEN_231 = r_sectored_hit ? sectored_entries_0_7_valid_0 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_232 = r_sectored_hit ? sectored_entries_0_7_valid_1 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_233 = r_sectored_hit ? sectored_entries_0_7_valid_2 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_234 = r_sectored_hit ? sectored_entries_0_7_valid_3 : 1'h0; // @[TLB.scala 252:32]
  assign _GEN_235 = _GEN_921 | _GEN_231; // @[TLB.scala 121:16]
  assign _GEN_236 = _GEN_922 | _GEN_232; // @[TLB.scala 121:16]
  assign _GEN_237 = _GEN_923 | _GEN_233; // @[TLB.scala 121:16]
  assign _GEN_238 = _GEN_924 | _GEN_234; // @[TLB.scala 121:16]
  assign _GEN_243 = invalidate_refill ? 1'h0 : _GEN_235; // @[TLB.scala 254:34]
  assign _GEN_244 = invalidate_refill ? 1'h0 : _GEN_236; // @[TLB.scala 254:34]
  assign _GEN_245 = invalidate_refill ? 1'h0 : _GEN_237; // @[TLB.scala 254:34]
  assign _GEN_246 = invalidate_refill ? 1'h0 : _GEN_238; // @[TLB.scala 254:34]
  assign _GEN_247 = _T_21 ? _GEN_243 : sectored_entries_0_7_valid_0; // @[TLB.scala 251:82]
  assign _GEN_248 = _T_21 ? _GEN_244 : sectored_entries_0_7_valid_1; // @[TLB.scala 251:82]
  assign _GEN_249 = _T_21 ? _GEN_245 : sectored_entries_0_7_valid_2; // @[TLB.scala 251:82]
  assign _GEN_250 = _T_21 ? _GEN_246 : sectored_entries_0_7_valid_3; // @[TLB.scala 251:82]
  assign _GEN_259 = _T_2 ? _GEN_35 : superpage_entries_0_valid_0; // @[TLB.scala 243:54]
  assign _GEN_263 = _T_2 ? _GEN_39 : superpage_entries_1_valid_0; // @[TLB.scala 243:54]
  assign _GEN_267 = _T_2 ? _GEN_43 : superpage_entries_2_valid_0; // @[TLB.scala 243:54]
  assign _GEN_271 = _T_2 ? _GEN_47 : superpage_entries_3_valid_0; // @[TLB.scala 243:54]
  assign _GEN_273 = _T_2 ? sectored_entries_0_0_valid_0 : _GEN_65; // @[TLB.scala 243:54]
  assign _GEN_274 = _T_2 ? sectored_entries_0_0_valid_1 : _GEN_66; // @[TLB.scala 243:54]
  assign _GEN_275 = _T_2 ? sectored_entries_0_0_valid_2 : _GEN_67; // @[TLB.scala 243:54]
  assign _GEN_276 = _T_2 ? sectored_entries_0_0_valid_3 : _GEN_68; // @[TLB.scala 243:54]
  assign _GEN_283 = _T_2 ? sectored_entries_0_1_valid_0 : _GEN_91; // @[TLB.scala 243:54]
  assign _GEN_284 = _T_2 ? sectored_entries_0_1_valid_1 : _GEN_92; // @[TLB.scala 243:54]
  assign _GEN_285 = _T_2 ? sectored_entries_0_1_valid_2 : _GEN_93; // @[TLB.scala 243:54]
  assign _GEN_286 = _T_2 ? sectored_entries_0_1_valid_3 : _GEN_94; // @[TLB.scala 243:54]
  assign _GEN_293 = _T_2 ? sectored_entries_0_2_valid_0 : _GEN_117; // @[TLB.scala 243:54]
  assign _GEN_294 = _T_2 ? sectored_entries_0_2_valid_1 : _GEN_118; // @[TLB.scala 243:54]
  assign _GEN_295 = _T_2 ? sectored_entries_0_2_valid_2 : _GEN_119; // @[TLB.scala 243:54]
  assign _GEN_296 = _T_2 ? sectored_entries_0_2_valid_3 : _GEN_120; // @[TLB.scala 243:54]
  assign _GEN_303 = _T_2 ? sectored_entries_0_3_valid_0 : _GEN_143; // @[TLB.scala 243:54]
  assign _GEN_304 = _T_2 ? sectored_entries_0_3_valid_1 : _GEN_144; // @[TLB.scala 243:54]
  assign _GEN_305 = _T_2 ? sectored_entries_0_3_valid_2 : _GEN_145; // @[TLB.scala 243:54]
  assign _GEN_306 = _T_2 ? sectored_entries_0_3_valid_3 : _GEN_146; // @[TLB.scala 243:54]
  assign _GEN_313 = _T_2 ? sectored_entries_0_4_valid_0 : _GEN_169; // @[TLB.scala 243:54]
  assign _GEN_314 = _T_2 ? sectored_entries_0_4_valid_1 : _GEN_170; // @[TLB.scala 243:54]
  assign _GEN_315 = _T_2 ? sectored_entries_0_4_valid_2 : _GEN_171; // @[TLB.scala 243:54]
  assign _GEN_316 = _T_2 ? sectored_entries_0_4_valid_3 : _GEN_172; // @[TLB.scala 243:54]
  assign _GEN_323 = _T_2 ? sectored_entries_0_5_valid_0 : _GEN_195; // @[TLB.scala 243:54]
  assign _GEN_324 = _T_2 ? sectored_entries_0_5_valid_1 : _GEN_196; // @[TLB.scala 243:54]
  assign _GEN_325 = _T_2 ? sectored_entries_0_5_valid_2 : _GEN_197; // @[TLB.scala 243:54]
  assign _GEN_326 = _T_2 ? sectored_entries_0_5_valid_3 : _GEN_198; // @[TLB.scala 243:54]
  assign _GEN_333 = _T_2 ? sectored_entries_0_6_valid_0 : _GEN_221; // @[TLB.scala 243:54]
  assign _GEN_334 = _T_2 ? sectored_entries_0_6_valid_1 : _GEN_222; // @[TLB.scala 243:54]
  assign _GEN_335 = _T_2 ? sectored_entries_0_6_valid_2 : _GEN_223; // @[TLB.scala 243:54]
  assign _GEN_336 = _T_2 ? sectored_entries_0_6_valid_3 : _GEN_224; // @[TLB.scala 243:54]
  assign _GEN_343 = _T_2 ? sectored_entries_0_7_valid_0 : _GEN_247; // @[TLB.scala 243:54]
  assign _GEN_344 = _T_2 ? sectored_entries_0_7_valid_1 : _GEN_248; // @[TLB.scala 243:54]
  assign _GEN_345 = _T_2 ? sectored_entries_0_7_valid_2 : _GEN_249; // @[TLB.scala 243:54]
  assign _GEN_346 = _T_2 ? sectored_entries_0_7_valid_3 : _GEN_250; // @[TLB.scala 243:54]
  assign _GEN_355 = io_ptw_resp_bits_homogeneous ? special_entry_valid_0 : _GEN_32; // @[TLB.scala 238:68]
  assign _GEN_359 = io_ptw_resp_bits_homogeneous ? _GEN_259 : superpage_entries_0_valid_0; // @[TLB.scala 238:68]
  assign _GEN_363 = io_ptw_resp_bits_homogeneous ? _GEN_263 : superpage_entries_1_valid_0; // @[TLB.scala 238:68]
  assign _GEN_367 = io_ptw_resp_bits_homogeneous ? _GEN_267 : superpage_entries_2_valid_0; // @[TLB.scala 238:68]
  assign _GEN_371 = io_ptw_resp_bits_homogeneous ? _GEN_271 : superpage_entries_3_valid_0; // @[TLB.scala 238:68]
  assign _GEN_373 = io_ptw_resp_bits_homogeneous ? _GEN_273 : sectored_entries_0_0_valid_0; // @[TLB.scala 238:68]
  assign _GEN_374 = io_ptw_resp_bits_homogeneous ? _GEN_274 : sectored_entries_0_0_valid_1; // @[TLB.scala 238:68]
  assign _GEN_375 = io_ptw_resp_bits_homogeneous ? _GEN_275 : sectored_entries_0_0_valid_2; // @[TLB.scala 238:68]
  assign _GEN_376 = io_ptw_resp_bits_homogeneous ? _GEN_276 : sectored_entries_0_0_valid_3; // @[TLB.scala 238:68]
  assign _GEN_383 = io_ptw_resp_bits_homogeneous ? _GEN_283 : sectored_entries_0_1_valid_0; // @[TLB.scala 238:68]
  assign _GEN_384 = io_ptw_resp_bits_homogeneous ? _GEN_284 : sectored_entries_0_1_valid_1; // @[TLB.scala 238:68]
  assign _GEN_385 = io_ptw_resp_bits_homogeneous ? _GEN_285 : sectored_entries_0_1_valid_2; // @[TLB.scala 238:68]
  assign _GEN_386 = io_ptw_resp_bits_homogeneous ? _GEN_286 : sectored_entries_0_1_valid_3; // @[TLB.scala 238:68]
  assign _GEN_393 = io_ptw_resp_bits_homogeneous ? _GEN_293 : sectored_entries_0_2_valid_0; // @[TLB.scala 238:68]
  assign _GEN_394 = io_ptw_resp_bits_homogeneous ? _GEN_294 : sectored_entries_0_2_valid_1; // @[TLB.scala 238:68]
  assign _GEN_395 = io_ptw_resp_bits_homogeneous ? _GEN_295 : sectored_entries_0_2_valid_2; // @[TLB.scala 238:68]
  assign _GEN_396 = io_ptw_resp_bits_homogeneous ? _GEN_296 : sectored_entries_0_2_valid_3; // @[TLB.scala 238:68]
  assign _GEN_403 = io_ptw_resp_bits_homogeneous ? _GEN_303 : sectored_entries_0_3_valid_0; // @[TLB.scala 238:68]
  assign _GEN_404 = io_ptw_resp_bits_homogeneous ? _GEN_304 : sectored_entries_0_3_valid_1; // @[TLB.scala 238:68]
  assign _GEN_405 = io_ptw_resp_bits_homogeneous ? _GEN_305 : sectored_entries_0_3_valid_2; // @[TLB.scala 238:68]
  assign _GEN_406 = io_ptw_resp_bits_homogeneous ? _GEN_306 : sectored_entries_0_3_valid_3; // @[TLB.scala 238:68]
  assign _GEN_413 = io_ptw_resp_bits_homogeneous ? _GEN_313 : sectored_entries_0_4_valid_0; // @[TLB.scala 238:68]
  assign _GEN_414 = io_ptw_resp_bits_homogeneous ? _GEN_314 : sectored_entries_0_4_valid_1; // @[TLB.scala 238:68]
  assign _GEN_415 = io_ptw_resp_bits_homogeneous ? _GEN_315 : sectored_entries_0_4_valid_2; // @[TLB.scala 238:68]
  assign _GEN_416 = io_ptw_resp_bits_homogeneous ? _GEN_316 : sectored_entries_0_4_valid_3; // @[TLB.scala 238:68]
  assign _GEN_423 = io_ptw_resp_bits_homogeneous ? _GEN_323 : sectored_entries_0_5_valid_0; // @[TLB.scala 238:68]
  assign _GEN_424 = io_ptw_resp_bits_homogeneous ? _GEN_324 : sectored_entries_0_5_valid_1; // @[TLB.scala 238:68]
  assign _GEN_425 = io_ptw_resp_bits_homogeneous ? _GEN_325 : sectored_entries_0_5_valid_2; // @[TLB.scala 238:68]
  assign _GEN_426 = io_ptw_resp_bits_homogeneous ? _GEN_326 : sectored_entries_0_5_valid_3; // @[TLB.scala 238:68]
  assign _GEN_433 = io_ptw_resp_bits_homogeneous ? _GEN_333 : sectored_entries_0_6_valid_0; // @[TLB.scala 238:68]
  assign _GEN_434 = io_ptw_resp_bits_homogeneous ? _GEN_334 : sectored_entries_0_6_valid_1; // @[TLB.scala 238:68]
  assign _GEN_435 = io_ptw_resp_bits_homogeneous ? _GEN_335 : sectored_entries_0_6_valid_2; // @[TLB.scala 238:68]
  assign _GEN_436 = io_ptw_resp_bits_homogeneous ? _GEN_336 : sectored_entries_0_6_valid_3; // @[TLB.scala 238:68]
  assign _GEN_443 = io_ptw_resp_bits_homogeneous ? _GEN_343 : sectored_entries_0_7_valid_0; // @[TLB.scala 238:68]
  assign _GEN_444 = io_ptw_resp_bits_homogeneous ? _GEN_344 : sectored_entries_0_7_valid_1; // @[TLB.scala 238:68]
  assign _GEN_445 = io_ptw_resp_bits_homogeneous ? _GEN_345 : sectored_entries_0_7_valid_2; // @[TLB.scala 238:68]
  assign _GEN_446 = io_ptw_resp_bits_homogeneous ? _GEN_346 : sectored_entries_0_7_valid_3; // @[TLB.scala 238:68]
  assign _GEN_455 = io_ptw_resp_valid ? _GEN_355 : special_entry_valid_0; // @[TLB.scala 218:20]
  assign _GEN_459 = io_ptw_resp_valid ? _GEN_359 : superpage_entries_0_valid_0; // @[TLB.scala 218:20]
  assign _GEN_463 = io_ptw_resp_valid ? _GEN_363 : superpage_entries_1_valid_0; // @[TLB.scala 218:20]
  assign _GEN_467 = io_ptw_resp_valid ? _GEN_367 : superpage_entries_2_valid_0; // @[TLB.scala 218:20]
  assign _GEN_471 = io_ptw_resp_valid ? _GEN_371 : superpage_entries_3_valid_0; // @[TLB.scala 218:20]
  assign _GEN_473 = io_ptw_resp_valid ? _GEN_373 : sectored_entries_0_0_valid_0; // @[TLB.scala 218:20]
  assign _GEN_474 = io_ptw_resp_valid ? _GEN_374 : sectored_entries_0_0_valid_1; // @[TLB.scala 218:20]
  assign _GEN_475 = io_ptw_resp_valid ? _GEN_375 : sectored_entries_0_0_valid_2; // @[TLB.scala 218:20]
  assign _GEN_476 = io_ptw_resp_valid ? _GEN_376 : sectored_entries_0_0_valid_3; // @[TLB.scala 218:20]
  assign _GEN_483 = io_ptw_resp_valid ? _GEN_383 : sectored_entries_0_1_valid_0; // @[TLB.scala 218:20]
  assign _GEN_484 = io_ptw_resp_valid ? _GEN_384 : sectored_entries_0_1_valid_1; // @[TLB.scala 218:20]
  assign _GEN_485 = io_ptw_resp_valid ? _GEN_385 : sectored_entries_0_1_valid_2; // @[TLB.scala 218:20]
  assign _GEN_486 = io_ptw_resp_valid ? _GEN_386 : sectored_entries_0_1_valid_3; // @[TLB.scala 218:20]
  assign _GEN_493 = io_ptw_resp_valid ? _GEN_393 : sectored_entries_0_2_valid_0; // @[TLB.scala 218:20]
  assign _GEN_494 = io_ptw_resp_valid ? _GEN_394 : sectored_entries_0_2_valid_1; // @[TLB.scala 218:20]
  assign _GEN_495 = io_ptw_resp_valid ? _GEN_395 : sectored_entries_0_2_valid_2; // @[TLB.scala 218:20]
  assign _GEN_496 = io_ptw_resp_valid ? _GEN_396 : sectored_entries_0_2_valid_3; // @[TLB.scala 218:20]
  assign _GEN_503 = io_ptw_resp_valid ? _GEN_403 : sectored_entries_0_3_valid_0; // @[TLB.scala 218:20]
  assign _GEN_504 = io_ptw_resp_valid ? _GEN_404 : sectored_entries_0_3_valid_1; // @[TLB.scala 218:20]
  assign _GEN_505 = io_ptw_resp_valid ? _GEN_405 : sectored_entries_0_3_valid_2; // @[TLB.scala 218:20]
  assign _GEN_506 = io_ptw_resp_valid ? _GEN_406 : sectored_entries_0_3_valid_3; // @[TLB.scala 218:20]
  assign _GEN_513 = io_ptw_resp_valid ? _GEN_413 : sectored_entries_0_4_valid_0; // @[TLB.scala 218:20]
  assign _GEN_514 = io_ptw_resp_valid ? _GEN_414 : sectored_entries_0_4_valid_1; // @[TLB.scala 218:20]
  assign _GEN_515 = io_ptw_resp_valid ? _GEN_415 : sectored_entries_0_4_valid_2; // @[TLB.scala 218:20]
  assign _GEN_516 = io_ptw_resp_valid ? _GEN_416 : sectored_entries_0_4_valid_3; // @[TLB.scala 218:20]
  assign _GEN_523 = io_ptw_resp_valid ? _GEN_423 : sectored_entries_0_5_valid_0; // @[TLB.scala 218:20]
  assign _GEN_524 = io_ptw_resp_valid ? _GEN_424 : sectored_entries_0_5_valid_1; // @[TLB.scala 218:20]
  assign _GEN_525 = io_ptw_resp_valid ? _GEN_425 : sectored_entries_0_5_valid_2; // @[TLB.scala 218:20]
  assign _GEN_526 = io_ptw_resp_valid ? _GEN_426 : sectored_entries_0_5_valid_3; // @[TLB.scala 218:20]
  assign _GEN_533 = io_ptw_resp_valid ? _GEN_433 : sectored_entries_0_6_valid_0; // @[TLB.scala 218:20]
  assign _GEN_534 = io_ptw_resp_valid ? _GEN_434 : sectored_entries_0_6_valid_1; // @[TLB.scala 218:20]
  assign _GEN_535 = io_ptw_resp_valid ? _GEN_435 : sectored_entries_0_6_valid_2; // @[TLB.scala 218:20]
  assign _GEN_536 = io_ptw_resp_valid ? _GEN_436 : sectored_entries_0_6_valid_3; // @[TLB.scala 218:20]
  assign _GEN_543 = io_ptw_resp_valid ? _GEN_443 : sectored_entries_0_7_valid_0; // @[TLB.scala 218:20]
  assign _GEN_544 = io_ptw_resp_valid ? _GEN_444 : sectored_entries_0_7_valid_1; // @[TLB.scala 218:20]
  assign _GEN_545 = io_ptw_resp_valid ? _GEN_445 : sectored_entries_0_7_valid_2; // @[TLB.scala 218:20]
  assign _GEN_546 = io_ptw_resp_valid ? _GEN_446 : sectored_entries_0_7_valid_3; // @[TLB.scala 218:20]
  assign _GEN_554 = 2'h1 == hitsVec_idx ? sectored_entries_0_0_data_1 : sectored_entries_0_0_data_0;
  assign _GEN_555 = 2'h2 == hitsVec_idx ? sectored_entries_0_0_data_2 : _GEN_554;
  assign _GEN_556 = 2'h3 == hitsVec_idx ? sectored_entries_0_0_data_3 : _GEN_555;
  assign _GEN_558 = 2'h1 == hitsVec_idx ? sectored_entries_0_1_data_1 : sectored_entries_0_1_data_0;
  assign _GEN_559 = 2'h2 == hitsVec_idx ? sectored_entries_0_1_data_2 : _GEN_558;
  assign _GEN_560 = 2'h3 == hitsVec_idx ? sectored_entries_0_1_data_3 : _GEN_559;
  assign _GEN_562 = 2'h1 == hitsVec_idx ? sectored_entries_0_2_data_1 : sectored_entries_0_2_data_0;
  assign _GEN_563 = 2'h2 == hitsVec_idx ? sectored_entries_0_2_data_2 : _GEN_562;
  assign _GEN_564 = 2'h3 == hitsVec_idx ? sectored_entries_0_2_data_3 : _GEN_563;
  assign _GEN_566 = 2'h1 == hitsVec_idx ? sectored_entries_0_3_data_1 : sectored_entries_0_3_data_0;
  assign _GEN_567 = 2'h2 == hitsVec_idx ? sectored_entries_0_3_data_2 : _GEN_566;
  assign _GEN_568 = 2'h3 == hitsVec_idx ? sectored_entries_0_3_data_3 : _GEN_567;
  assign _GEN_570 = 2'h1 == hitsVec_idx ? sectored_entries_0_4_data_1 : sectored_entries_0_4_data_0;
  assign _GEN_571 = 2'h2 == hitsVec_idx ? sectored_entries_0_4_data_2 : _GEN_570;
  assign _GEN_572 = 2'h3 == hitsVec_idx ? sectored_entries_0_4_data_3 : _GEN_571;
  assign _GEN_574 = 2'h1 == hitsVec_idx ? sectored_entries_0_5_data_1 : sectored_entries_0_5_data_0;
  assign _GEN_575 = 2'h2 == hitsVec_idx ? sectored_entries_0_5_data_2 : _GEN_574;
  assign _GEN_576 = 2'h3 == hitsVec_idx ? sectored_entries_0_5_data_3 : _GEN_575;
  assign _GEN_578 = 2'h1 == hitsVec_idx ? sectored_entries_0_6_data_1 : sectored_entries_0_6_data_0;
  assign _GEN_579 = 2'h2 == hitsVec_idx ? sectored_entries_0_6_data_2 : _GEN_578;
  assign _GEN_580 = 2'h3 == hitsVec_idx ? sectored_entries_0_6_data_3 : _GEN_579;
  assign _GEN_582 = 2'h1 == hitsVec_idx ? sectored_entries_0_7_data_1 : sectored_entries_0_7_data_0;
  assign _GEN_583 = 2'h2 == hitsVec_idx ? sectored_entries_0_7_data_2 : _GEN_582;
  assign _GEN_584 = 2'h3 == hitsVec_idx ? sectored_entries_0_7_data_3 : _GEN_583;
  assign ppn_hi = entries_barrier_8_io_y_ppn[19:18]; // @[TLB.scala 105:26]
  assign _ppn_T_1 = superpage_hits_ignore_1 ? vpn : 27'h0; // @[TLB.scala 108:28]
  assign _GEN_953 = {{7'd0}, entries_barrier_8_io_y_ppn}; // @[TLB.scala 108:47]
  assign _ppn_T_2 = _ppn_T_1 | _GEN_953; // @[TLB.scala 108:47]
  assign ppn_lo = _ppn_T_2[17:9]; // @[TLB.scala 108:58]
  assign _ppn_T_4 = vpn | _GEN_953; // @[TLB.scala 108:47]
  assign ppn_lo_1 = _ppn_T_4[8:0]; // @[TLB.scala 108:58]
  assign _ppn_T_5 = {ppn_hi,ppn_lo,ppn_lo_1}; // @[Cat.scala 30:58]
  assign ppn_hi_2 = entries_barrier_9_io_y_ppn[19:18]; // @[TLB.scala 105:26]
  assign _ppn_T_6 = superpage_hits_ignore_4 ? vpn : 27'h0; // @[TLB.scala 108:28]
  assign _GEN_955 = {{7'd0}, entries_barrier_9_io_y_ppn}; // @[TLB.scala 108:47]
  assign _ppn_T_7 = _ppn_T_6 | _GEN_955; // @[TLB.scala 108:47]
  assign ppn_lo_2 = _ppn_T_7[17:9]; // @[TLB.scala 108:58]
  assign _ppn_T_9 = vpn | _GEN_955; // @[TLB.scala 108:47]
  assign ppn_lo_3 = _ppn_T_9[8:0]; // @[TLB.scala 108:58]
  assign _ppn_T_10 = {ppn_hi_2,ppn_lo_2,ppn_lo_3}; // @[Cat.scala 30:58]
  assign ppn_hi_4 = entries_barrier_10_io_y_ppn[19:18]; // @[TLB.scala 105:26]
  assign _ppn_T_11 = superpage_hits_ignore_7 ? vpn : 27'h0; // @[TLB.scala 108:28]
  assign _GEN_957 = {{7'd0}, entries_barrier_10_io_y_ppn}; // @[TLB.scala 108:47]
  assign _ppn_T_12 = _ppn_T_11 | _GEN_957; // @[TLB.scala 108:47]
  assign ppn_lo_4 = _ppn_T_12[17:9]; // @[TLB.scala 108:58]
  assign _ppn_T_14 = vpn | _GEN_957; // @[TLB.scala 108:47]
  assign ppn_lo_5 = _ppn_T_14[8:0]; // @[TLB.scala 108:58]
  assign _ppn_T_15 = {ppn_hi_4,ppn_lo_4,ppn_lo_5}; // @[Cat.scala 30:58]
  assign ppn_hi_6 = entries_barrier_11_io_y_ppn[19:18]; // @[TLB.scala 105:26]
  assign _ppn_T_16 = superpage_hits_ignore_10 ? vpn : 27'h0; // @[TLB.scala 108:28]
  assign _GEN_959 = {{7'd0}, entries_barrier_11_io_y_ppn}; // @[TLB.scala 108:47]
  assign _ppn_T_17 = _ppn_T_16 | _GEN_959; // @[TLB.scala 108:47]
  assign ppn_lo_6 = _ppn_T_17[17:9]; // @[TLB.scala 108:58]
  assign _ppn_T_19 = vpn | _GEN_959; // @[TLB.scala 108:47]
  assign ppn_lo_7 = _ppn_T_19[8:0]; // @[TLB.scala 108:58]
  assign _ppn_T_20 = {ppn_hi_6,ppn_lo_6,ppn_lo_7}; // @[Cat.scala 30:58]
  assign ppn_hi_8 = entries_barrier_12_io_y_ppn[19:18]; // @[TLB.scala 105:26]
  assign _GEN_961 = {{7'd0}, entries_barrier_12_io_y_ppn}; // @[TLB.scala 108:47]
  assign _ppn_T_22 = _mpu_ppn_T_17 | _GEN_961; // @[TLB.scala 108:47]
  assign ppn_lo_8 = _ppn_T_22[17:9]; // @[TLB.scala 108:58]
  assign _ppn_T_24 = _mpu_ppn_T_19 | _GEN_961; // @[TLB.scala 108:47]
  assign ppn_lo_9 = _ppn_T_24[8:0]; // @[TLB.scala 108:58]
  assign _ppn_T_25 = {ppn_hi_8,ppn_lo_8,ppn_lo_9}; // @[Cat.scala 30:58]
  assign _ppn_T_27 = hitsVec_0 ? entries_barrier_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  assign _ppn_T_28 = hitsVec_1 ? entries_barrier_1_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  assign _ppn_T_29 = hitsVec_2 ? entries_barrier_2_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  assign _ppn_T_30 = hitsVec_3 ? entries_barrier_3_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  assign _ppn_T_31 = hitsVec_4 ? entries_barrier_4_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  assign _ppn_T_32 = hitsVec_5 ? entries_barrier_5_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  assign _ppn_T_33 = hitsVec_6 ? entries_barrier_6_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  assign _ppn_T_34 = hitsVec_7 ? entries_barrier_7_io_y_ppn : 20'h0; // @[Mux.scala 27:72]
  assign _ppn_T_35 = hitsVec_8 ? _ppn_T_5 : 20'h0; // @[Mux.scala 27:72]
  assign _ppn_T_36 = hitsVec_9 ? _ppn_T_10 : 20'h0; // @[Mux.scala 27:72]
  assign _ppn_T_37 = hitsVec_10 ? _ppn_T_15 : 20'h0; // @[Mux.scala 27:72]
  assign _ppn_T_38 = hitsVec_11 ? _ppn_T_20 : 20'h0; // @[Mux.scala 27:72]
  assign _ppn_T_39 = hitsVec_12 ? _ppn_T_25 : 20'h0; // @[Mux.scala 27:72]
  assign _ppn_T_40 = hits_hi ? vpn[19:0] : 20'h0; // @[Mux.scala 27:72]
  assign _ppn_T_41 = _ppn_T_27 | _ppn_T_28; // @[Mux.scala 27:72]
  assign _ppn_T_42 = _ppn_T_41 | _ppn_T_29; // @[Mux.scala 27:72]
  assign _ppn_T_43 = _ppn_T_42 | _ppn_T_30; // @[Mux.scala 27:72]
  assign _ppn_T_44 = _ppn_T_43 | _ppn_T_31; // @[Mux.scala 27:72]
  assign _ppn_T_45 = _ppn_T_44 | _ppn_T_32; // @[Mux.scala 27:72]
  assign _ppn_T_46 = _ppn_T_45 | _ppn_T_33; // @[Mux.scala 27:72]
  assign _ppn_T_47 = _ppn_T_46 | _ppn_T_34; // @[Mux.scala 27:72]
  assign _ppn_T_48 = _ppn_T_47 | _ppn_T_35; // @[Mux.scala 27:72]
  assign _ppn_T_49 = _ppn_T_48 | _ppn_T_36; // @[Mux.scala 27:72]
  assign _ppn_T_50 = _ppn_T_49 | _ppn_T_37; // @[Mux.scala 27:72]
  assign _ppn_T_51 = _ppn_T_50 | _ppn_T_38; // @[Mux.scala 27:72]
  assign _ppn_T_52 = _ppn_T_51 | _ppn_T_39; // @[Mux.scala 27:72]
  assign ppn = _ppn_T_52 | _ppn_T_40; // @[Mux.scala 27:72]
  assign ptw_ae_array_lo = {entries_barrier_5_io_y_ae,entries_barrier_4_io_y_ae,entries_barrier_3_io_y_ae,entries_barrier_2_io_y_ae,entries_barrier_1_io_y_ae,entries_barrier_io_y_ae}; // @[Cat.scala 30:58]
  assign ptw_ae_array = {1'h0,entries_barrier_12_io_y_ae,entries_barrier_11_io_y_ae,entries_barrier_10_io_y_ae,entries_barrier_9_io_y_ae,entries_barrier_8_io_y_ae,entries_barrier_7_io_y_ae,entries_barrier_6_io_y_ae,ptw_ae_array_lo}; // @[Cat.scala 30:58]
  assign priv_rw_ok_lo = {entries_barrier_5_io_y_u,entries_barrier_4_io_y_u,entries_barrier_3_io_y_u,entries_barrier_2_io_y_u,entries_barrier_1_io_y_u,entries_barrier_io_y_u}; // @[Cat.scala 30:58]
  assign _priv_rw_ok_T_2 = {entries_barrier_12_io_y_u,entries_barrier_11_io_y_u,entries_barrier_10_io_y_u,entries_barrier_9_io_y_u,entries_barrier_8_io_y_u,entries_barrier_7_io_y_u,entries_barrier_6_io_y_u,priv_rw_ok_lo}; // @[Cat.scala 30:58]
  assign priv_x_ok = priv_s ? ~_priv_rw_ok_T_2 : _priv_rw_ok_T_2; // @[TLB.scala 266:22]
  assign r_array_lo_1 = {entries_barrier_5_io_y_sx,entries_barrier_4_io_y_sx,entries_barrier_3_io_y_sx,entries_barrier_2_io_y_sx,entries_barrier_1_io_y_sx,entries_barrier_io_y_sx}; // @[Cat.scala 30:58]
  assign _r_array_T_1 = {entries_barrier_12_io_y_sx,entries_barrier_11_io_y_sx,entries_barrier_10_io_y_sx,entries_barrier_9_io_y_sx,entries_barrier_8_io_y_sx,entries_barrier_7_io_y_sx,entries_barrier_6_io_y_sx,r_array_lo_1}; // @[Cat.scala 30:58]
  assign x_array_lo_1 = priv_x_ok & _r_array_T_1; // @[TLB.scala 269:39]
  assign x_array = {1'h1,x_array_lo_1}; // @[Cat.scala 30:58]
  assign px_array_hi = prot_x ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  assign px_array_lo = {entries_barrier_5_io_y_px,entries_barrier_4_io_y_px,entries_barrier_3_io_y_px,entries_barrier_2_io_y_px,entries_barrier_1_io_y_px,entries_barrier_io_y_px}; // @[Cat.scala 30:58]
  assign _px_array_T_1 = {px_array_hi,entries_barrier_11_io_y_px,entries_barrier_10_io_y_px,entries_barrier_9_io_y_px,entries_barrier_8_io_y_px,entries_barrier_7_io_y_px,entries_barrier_6_io_y_px,px_array_lo}; // @[Cat.scala 30:58]
  assign px_array = _px_array_T_1 & ~ptw_ae_array; // @[TLB.scala 272:87]
  assign c_array_hi = cacheable ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  assign c_array_lo = {entries_barrier_5_io_y_c,entries_barrier_4_io_y_c,entries_barrier_3_io_y_c,entries_barrier_2_io_y_c,entries_barrier_1_io_y_c,entries_barrier_io_y_c}; // @[Cat.scala 30:58]
  assign c_array = {c_array_hi,entries_barrier_11_io_y_c,entries_barrier_10_io_y_c,entries_barrier_9_io_y_c,entries_barrier_8_io_y_c,entries_barrier_7_io_y_c,entries_barrier_6_io_y_c,c_array_lo}; // @[Cat.scala 30:58]
  assign bad_va_maskedVAddr = io_req_bits_vaddr & 40'hc000000000; // @[TLB.scala 289:43]
  assign _bad_va_T_1 = bad_va_maskedVAddr == 40'h0; // @[TLB.scala 290:61]
  assign _bad_va_T_2 = bad_va_maskedVAddr == 40'hc000000000; // @[TLB.scala 290:82]
  assign _bad_va_T_3 = _bad_va_T_1 | _bad_va_T_2; // @[TLB.scala 290:67]
  assign bad_va = vm_enabled & ~_bad_va_T_3; // @[TLB.scala 284:117]
  assign _pf_inst_array_T = x_array | ptw_ae_array; // @[TLB.scala 322:33]
  assign pf_inst_array = ~_pf_inst_array_T; // @[TLB.scala 322:23]
  assign tlb_hit = |real_hits; // @[TLB.scala 324:27]
  assign _tlb_miss_T_1 = vm_enabled & ~bad_va; // @[TLB.scala 325:29]
  assign tlb_miss = _tlb_miss_T_1 & ~tlb_hit; // @[TLB.scala 325:40]
  assign _T_23 = io_req_valid & vm_enabled; // @[TLB.scala 329:22]
  assign _T_24 = sector_hits_0 | sector_hits_1; // @[package.scala 72:59]
  assign _T_25 = _T_24 | sector_hits_2; // @[package.scala 72:59]
  assign _T_26 = _T_25 | sector_hits_3; // @[package.scala 72:59]
  assign _T_27 = _T_26 | sector_hits_4; // @[package.scala 72:59]
  assign _T_28 = _T_27 | sector_hits_5; // @[package.scala 72:59]
  assign _T_29 = _T_28 | sector_hits_6; // @[package.scala 72:59]
  assign _T_30 = _T_29 | sector_hits_7; // @[package.scala 72:59]
  assign _T_31 = {sector_hits_7,sector_hits_6,sector_hits_5,sector_hits_4,sector_hits_3,sector_hits_2,sector_hits_1,sector_hits_0}; // @[Cat.scala 30:58]
  assign hi_1 = _T_31[7:4]; // @[OneHot.scala 30:18]
  assign lo_1 = _T_31[3:0]; // @[OneHot.scala 31:18]
  assign hi_2 = |hi_1; // @[OneHot.scala 32:14]
  assign _T_32 = hi_1 | lo_1; // @[OneHot.scala 32:28]
  assign hi_3 = _T_32[3:2]; // @[OneHot.scala 30:18]
  assign lo_2 = _T_32[1:0]; // @[OneHot.scala 31:18]
  assign hi_4 = |hi_3; // @[OneHot.scala 32:14]
  assign _T_33 = hi_3 | lo_2; // @[OneHot.scala 32:28]
  assign lo_3 = _T_33[1]; // @[CircuitMath.scala 30:8]
  assign state_vec_0_touch_way_sized = {hi_2,hi_4,lo_3}; // @[Cat.scala 30:58]
  assign state_vec_0_hi_hi = ~state_vec_0_touch_way_sized[2]; // @[Replacement.scala 196:33]
  assign state_vec_0_left_subtree_state = state_vec_0[5:3]; // @[package.scala 154:13]
  assign state_vec_0_right_subtree_state = state_vec_0[2:0]; // @[Replacement.scala 198:38]
  assign state_vec_0_hi_hi_1 = ~state_vec_0_touch_way_sized[1]; // @[Replacement.scala 196:33]
  assign state_vec_0_left_subtree_state_1 = state_vec_0_left_subtree_state[1]; // @[package.scala 154:13]
  assign state_vec_0_right_subtree_state_1 = state_vec_0_left_subtree_state[0]; // @[Replacement.scala 198:38]
  assign state_vec_0_hi_lo = state_vec_0_hi_hi_1 ? state_vec_0_left_subtree_state_1 : ~state_vec_0_touch_way_sized[0]; // @[Replacement.scala 203:16]
  assign state_vec_0_lo = state_vec_0_hi_hi_1 ? ~state_vec_0_touch_way_sized[0] : state_vec_0_right_subtree_state_1; // @[Replacement.scala 206:16]
  assign _state_vec_0_T_7 = {state_vec_0_hi_hi_1,state_vec_0_hi_lo,state_vec_0_lo}; // @[Cat.scala 30:58]
  assign state_vec_0_hi_lo_1 = state_vec_0_hi_hi ? state_vec_0_left_subtree_state : _state_vec_0_T_7; // @[Replacement.scala 203:16]
  assign state_vec_0_left_subtree_state_2 = state_vec_0_right_subtree_state[1]; // @[package.scala 154:13]
  assign state_vec_0_right_subtree_state_2 = state_vec_0_right_subtree_state[0]; // @[Replacement.scala 198:38]
  assign state_vec_0_hi_lo_2 = state_vec_0_hi_hi_1 ? state_vec_0_left_subtree_state_2 : ~state_vec_0_touch_way_sized[0]; // @[Replacement.scala 203:16]
  assign state_vec_0_lo_1 = state_vec_0_hi_hi_1 ? ~state_vec_0_touch_way_sized[0] : state_vec_0_right_subtree_state_2; // @[Replacement.scala 206:16]
  assign _state_vec_0_T_15 = {state_vec_0_hi_hi_1,state_vec_0_hi_lo_2,state_vec_0_lo_1}; // @[Cat.scala 30:58]
  assign state_vec_0_lo_2 = state_vec_0_hi_hi ? _state_vec_0_T_15 : state_vec_0_right_subtree_state; // @[Replacement.scala 206:16]
  assign _state_vec_0_T_16 = {state_vec_0_hi_hi,state_vec_0_hi_lo_1,state_vec_0_lo_2}; // @[Cat.scala 30:58]
  assign _T_35 = superpage_hits_0 | superpage_hits_1; // @[package.scala 72:59]
  assign _T_36 = _T_35 | superpage_hits_2; // @[package.scala 72:59]
  assign _T_37 = _T_36 | superpage_hits_3; // @[package.scala 72:59]
  assign _T_38 = {superpage_hits_3,superpage_hits_2,superpage_hits_1,superpage_hits_0}; // @[Cat.scala 30:58]
  assign hi_6 = _T_38[3:2]; // @[OneHot.scala 30:18]
  assign lo_6 = _T_38[1:0]; // @[OneHot.scala 31:18]
  assign hi_7 = |hi_6; // @[OneHot.scala 32:14]
  assign _T_39 = hi_6 | lo_6; // @[OneHot.scala 32:28]
  assign lo_7 = _T_39[1]; // @[CircuitMath.scala 30:8]
  assign state_reg_touch_way_sized = {hi_7,lo_7}; // @[Cat.scala 30:58]
  assign state_reg_hi_hi = ~state_reg_touch_way_sized[1]; // @[Replacement.scala 196:33]
  assign state_reg_left_subtree_state = state_reg_1[1]; // @[package.scala 154:13]
  assign state_reg_right_subtree_state = state_reg_1[0]; // @[Replacement.scala 198:38]
  assign state_reg_hi_lo = state_reg_hi_hi ? state_reg_left_subtree_state : ~state_reg_touch_way_sized[0]; // @[Replacement.scala 203:16]
  assign state_reg_lo = state_reg_hi_hi ? ~state_reg_touch_way_sized[0] : state_reg_right_subtree_state; // @[Replacement.scala 206:16]
  assign _state_reg_T_6 = {state_reg_hi_hi,state_reg_hi_lo,state_reg_lo}; // @[Cat.scala 30:58]
  assign multipleHits_leftOne = real_hits[0]; // @[Misc.scala 180:37]
  assign multipleHits_leftOne_1 = real_hits[1]; // @[Misc.scala 180:37]
  assign multipleHits_rightOne = real_hits[2]; // @[Misc.scala 181:39]
  assign multipleHits_rightOne_1 = multipleHits_leftOne_1 | multipleHits_rightOne; // @[Misc.scala 182:16]
  assign multipleHits_rightTwo = multipleHits_leftOne_1 & multipleHits_rightOne; // @[Misc.scala 182:61]
  assign multipleHits_leftOne_2 = multipleHits_leftOne | multipleHits_rightOne_1; // @[Misc.scala 182:16]
  assign _multipleHits_T_9 = multipleHits_leftOne & multipleHits_rightOne_1; // @[Misc.scala 182:61]
  assign multipleHits_leftTwo = multipleHits_rightTwo | _multipleHits_T_9; // @[Misc.scala 182:49]
  assign multipleHits_leftOne_3 = real_hits[3]; // @[Misc.scala 180:37]
  assign multipleHits_leftOne_4 = real_hits[4]; // @[Misc.scala 180:37]
  assign multipleHits_rightOne_2 = real_hits[5]; // @[Misc.scala 181:39]
  assign multipleHits_rightOne_3 = multipleHits_leftOne_4 | multipleHits_rightOne_2; // @[Misc.scala 182:16]
  assign multipleHits_rightTwo_1 = multipleHits_leftOne_4 & multipleHits_rightOne_2; // @[Misc.scala 182:61]
  assign multipleHits_rightOne_4 = multipleHits_leftOne_3 | multipleHits_rightOne_3; // @[Misc.scala 182:16]
  assign _multipleHits_T_18 = multipleHits_leftOne_3 & multipleHits_rightOne_3; // @[Misc.scala 182:61]
  assign multipleHits_rightTwo_2 = multipleHits_rightTwo_1 | _multipleHits_T_18; // @[Misc.scala 182:49]
  assign multipleHits_leftOne_5 = multipleHits_leftOne_2 | multipleHits_rightOne_4; // @[Misc.scala 182:16]
  assign _multipleHits_T_19 = multipleHits_leftTwo | multipleHits_rightTwo_2; // @[Misc.scala 182:37]
  assign _multipleHits_T_20 = multipleHits_leftOne_2 & multipleHits_rightOne_4; // @[Misc.scala 182:61]
  assign multipleHits_leftTwo_1 = _multipleHits_T_19 | _multipleHits_T_20; // @[Misc.scala 182:49]
  assign multipleHits_leftOne_6 = real_hits[6]; // @[Misc.scala 180:37]
  assign multipleHits_leftOne_7 = real_hits[7]; // @[Misc.scala 180:37]
  assign multipleHits_rightOne_5 = real_hits[8]; // @[Misc.scala 181:39]
  assign multipleHits_rightOne_6 = multipleHits_leftOne_7 | multipleHits_rightOne_5; // @[Misc.scala 182:16]
  assign multipleHits_rightTwo_3 = multipleHits_leftOne_7 & multipleHits_rightOne_5; // @[Misc.scala 182:61]
  assign multipleHits_leftOne_8 = multipleHits_leftOne_6 | multipleHits_rightOne_6; // @[Misc.scala 182:16]
  assign _multipleHits_T_30 = multipleHits_leftOne_6 & multipleHits_rightOne_6; // @[Misc.scala 182:61]
  assign multipleHits_leftTwo_2 = multipleHits_rightTwo_3 | _multipleHits_T_30; // @[Misc.scala 182:49]
  assign multipleHits_leftOne_9 = real_hits[9]; // @[Misc.scala 180:37]
  assign multipleHits_rightOne_7 = real_hits[10]; // @[Misc.scala 181:39]
  assign multipleHits_leftOne_10 = multipleHits_leftOne_9 | multipleHits_rightOne_7; // @[Misc.scala 182:16]
  assign multipleHits_leftTwo_3 = multipleHits_leftOne_9 & multipleHits_rightOne_7; // @[Misc.scala 182:61]
  assign multipleHits_leftOne_11 = real_hits[11]; // @[Misc.scala 180:37]
  assign multipleHits_rightOne_8 = real_hits[12]; // @[Misc.scala 181:39]
  assign multipleHits_rightOne_9 = multipleHits_leftOne_11 | multipleHits_rightOne_8; // @[Misc.scala 182:16]
  assign multipleHits_rightTwo_4 = multipleHits_leftOne_11 & multipleHits_rightOne_8; // @[Misc.scala 182:61]
  assign multipleHits_rightOne_10 = multipleHits_leftOne_10 | multipleHits_rightOne_9; // @[Misc.scala 182:16]
  assign _multipleHits_T_42 = multipleHits_leftTwo_3 | multipleHits_rightTwo_4; // @[Misc.scala 182:37]
  assign _multipleHits_T_43 = multipleHits_leftOne_10 & multipleHits_rightOne_9; // @[Misc.scala 182:61]
  assign multipleHits_rightTwo_5 = _multipleHits_T_42 | _multipleHits_T_43; // @[Misc.scala 182:49]
  assign multipleHits_rightOne_11 = multipleHits_leftOne_8 | multipleHits_rightOne_10; // @[Misc.scala 182:16]
  assign _multipleHits_T_44 = multipleHits_leftTwo_2 | multipleHits_rightTwo_5; // @[Misc.scala 182:37]
  assign _multipleHits_T_45 = multipleHits_leftOne_8 & multipleHits_rightOne_10; // @[Misc.scala 182:61]
  assign multipleHits_rightTwo_6 = _multipleHits_T_44 | _multipleHits_T_45; // @[Misc.scala 182:49]
  assign _multipleHits_T_47 = multipleHits_leftTwo_1 | multipleHits_rightTwo_6; // @[Misc.scala 182:37]
  assign _multipleHits_T_48 = multipleHits_leftOne_5 & multipleHits_rightOne_11; // @[Misc.scala 182:61]
  assign multipleHits = _multipleHits_T_47 | _multipleHits_T_48; // @[Misc.scala 182:49]
  assign _io_resp_pf_inst_T = pf_inst_array & hits; // @[TLB.scala 344:47]
  assign _io_resp_pf_inst_T_1 = |_io_resp_pf_inst_T; // @[TLB.scala 344:55]
  assign _io_resp_ae_inst_T_1 = ~px_array & hits; // @[TLB.scala 347:33]
  assign _io_resp_cacheable_T = c_array & hits; // @[TLB.scala 351:33]
  assign _io_resp_miss_T = io_ptw_resp_valid | tlb_miss; // @[TLB.scala 354:29]
  assign _T_41 = io_req_ready & io_req_valid; // @[Decoupled.scala 40:37]
  assign _T_42 = _T_41 & tlb_miss; // @[TLB.scala 363:25]
  assign r_superpage_repl_addr_hi = state_reg_1[2]; // @[Replacement.scala 243:38]
  assign r_superpage_repl_addr_lo = r_superpage_repl_addr_hi ? state_reg_left_subtree_state : state_reg_right_subtree_state; // @[Replacement.scala 250:16]
  assign _r_superpage_repl_addr_T_2 = {r_superpage_repl_addr_hi,r_superpage_repl_addr_lo}; // @[Cat.scala 30:58]
  assign r_superpage_repl_addr_valids = {superpage_entries_3_valid_0,superpage_entries_2_valid_0,superpage_entries_1_valid_0,superpage_entries_0_valid_0}; // @[Cat.scala 30:58]
  assign _r_superpage_repl_addr_T_3 = &r_superpage_repl_addr_valids; // @[TLB.scala 411:16]
  assign _r_superpage_repl_addr_T_5 = ~r_superpage_repl_addr_valids[0]; // @[OneHot.scala 47:40]
  assign _r_superpage_repl_addr_T_6 = ~r_superpage_repl_addr_valids[1]; // @[OneHot.scala 47:40]
  assign _r_superpage_repl_addr_T_7 = ~r_superpage_repl_addr_valids[2]; // @[OneHot.scala 47:40]
  assign r_sectored_repl_addr_hi = state_vec_0[6]; // @[Replacement.scala 243:38]
  assign r_sectored_repl_addr_hi_1 = state_vec_0_left_subtree_state[2]; // @[Replacement.scala 243:38]
  assign r_sectored_repl_addr_lo = r_sectored_repl_addr_hi_1 ? state_vec_0_left_subtree_state_1 : state_vec_0_right_subtree_state_1; // @[Replacement.scala 250:16]
  assign _r_sectored_repl_addr_T_2 = {r_sectored_repl_addr_hi_1,r_sectored_repl_addr_lo}; // @[Cat.scala 30:58]
  assign r_sectored_repl_addr_hi_2 = state_vec_0_right_subtree_state[2]; // @[Replacement.scala 243:38]
  assign r_sectored_repl_addr_lo_1 = r_sectored_repl_addr_hi_2 ? state_vec_0_left_subtree_state_2 : state_vec_0_right_subtree_state_2; // @[Replacement.scala 250:16]
  assign _r_sectored_repl_addr_T_5 = {r_sectored_repl_addr_hi_2,r_sectored_repl_addr_lo_1}; // @[Cat.scala 30:58]
  assign r_sectored_repl_addr_lo_2 = r_sectored_repl_addr_hi ? _r_sectored_repl_addr_T_2 : _r_sectored_repl_addr_T_5; // @[Replacement.scala 250:16]
  assign _r_sectored_repl_addr_T_6 = {r_sectored_repl_addr_hi,r_sectored_repl_addr_lo_2}; // @[Cat.scala 30:58]
  assign r_sectored_repl_addr_valids = {_sector_hits_T_44,_sector_hits_T_38,_sector_hits_T_32,_sector_hits_T_26,_sector_hits_T_20,_sector_hits_T_14,_sector_hits_T_8,_sector_hits_T_2}; // @[Cat.scala 30:58]
  assign _r_sectored_repl_addr_T_7 = &r_sectored_repl_addr_valids; // @[TLB.scala 411:16]
  assign _r_sectored_repl_addr_T_9 = ~r_sectored_repl_addr_valids[0]; // @[OneHot.scala 47:40]
  assign _r_sectored_repl_addr_T_10 = ~r_sectored_repl_addr_valids[1]; // @[OneHot.scala 47:40]
  assign _r_sectored_repl_addr_T_11 = ~r_sectored_repl_addr_valids[2]; // @[OneHot.scala 47:40]
  assign _r_sectored_repl_addr_T_12 = ~r_sectored_repl_addr_valids[3]; // @[OneHot.scala 47:40]
  assign _r_sectored_repl_addr_T_13 = ~r_sectored_repl_addr_valids[4]; // @[OneHot.scala 47:40]
  assign _r_sectored_repl_addr_T_14 = ~r_sectored_repl_addr_valids[5]; // @[OneHot.scala 47:40]
  assign _r_sectored_repl_addr_T_15 = ~r_sectored_repl_addr_valids[6]; // @[OneHot.scala 47:40]
  assign _T_44 = state == 2'h2; // @[TLB.scala 377:17]
  assign _T_45 = _T_44 & io_sfence_valid; // @[TLB.scala 377:28]
  assign _T_48 = io_sfence_bits_addr[38:12] == vpn; // @[TLB.scala 385:72]
  assign _T_49 = ~io_sfence_bits_rs1 | _T_48; // @[TLB.scala 385:34]
  assign _T_51 = _T_49 | reset; // @[TLB.scala 385:13]
  assign _T_59 = _sector_hits_T_3[26:18] == 9'h0; // @[TLB.scala 134:61]
  assign _GEN_617 = sectored_entries_0_0_data_0[13] ? _GEN_473 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_618 = sectored_entries_0_0_data_1[13] ? _GEN_474 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_619 = sectored_entries_0_0_data_2[13] ? _GEN_475 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_620 = sectored_entries_0_0_data_3[13] ? _GEN_476 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_621 = io_sfence_bits_rs2 & _GEN_617; // @[TLB.scala 388:40]
  assign _GEN_622 = io_sfence_bits_rs2 & _GEN_618; // @[TLB.scala 388:40]
  assign _GEN_623 = io_sfence_bits_rs2 & _GEN_619; // @[TLB.scala 388:40]
  assign _GEN_624 = io_sfence_bits_rs2 & _GEN_620; // @[TLB.scala 388:40]
  assign _T_198 = _sector_hits_T_9[26:18] == 9'h0; // @[TLB.scala 134:61]
  assign _GEN_645 = sectored_entries_0_1_data_0[13] ? _GEN_483 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_646 = sectored_entries_0_1_data_1[13] ? _GEN_484 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_647 = sectored_entries_0_1_data_2[13] ? _GEN_485 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_648 = sectored_entries_0_1_data_3[13] ? _GEN_486 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_649 = io_sfence_bits_rs2 & _GEN_645; // @[TLB.scala 388:40]
  assign _GEN_650 = io_sfence_bits_rs2 & _GEN_646; // @[TLB.scala 388:40]
  assign _GEN_651 = io_sfence_bits_rs2 & _GEN_647; // @[TLB.scala 388:40]
  assign _GEN_652 = io_sfence_bits_rs2 & _GEN_648; // @[TLB.scala 388:40]
  assign _T_337 = _sector_hits_T_15[26:18] == 9'h0; // @[TLB.scala 134:61]
  assign _GEN_673 = sectored_entries_0_2_data_0[13] ? _GEN_493 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_674 = sectored_entries_0_2_data_1[13] ? _GEN_494 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_675 = sectored_entries_0_2_data_2[13] ? _GEN_495 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_676 = sectored_entries_0_2_data_3[13] ? _GEN_496 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_677 = io_sfence_bits_rs2 & _GEN_673; // @[TLB.scala 388:40]
  assign _GEN_678 = io_sfence_bits_rs2 & _GEN_674; // @[TLB.scala 388:40]
  assign _GEN_679 = io_sfence_bits_rs2 & _GEN_675; // @[TLB.scala 388:40]
  assign _GEN_680 = io_sfence_bits_rs2 & _GEN_676; // @[TLB.scala 388:40]
  assign _T_476 = _sector_hits_T_21[26:18] == 9'h0; // @[TLB.scala 134:61]
  assign _GEN_701 = sectored_entries_0_3_data_0[13] ? _GEN_503 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_702 = sectored_entries_0_3_data_1[13] ? _GEN_504 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_703 = sectored_entries_0_3_data_2[13] ? _GEN_505 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_704 = sectored_entries_0_3_data_3[13] ? _GEN_506 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_705 = io_sfence_bits_rs2 & _GEN_701; // @[TLB.scala 388:40]
  assign _GEN_706 = io_sfence_bits_rs2 & _GEN_702; // @[TLB.scala 388:40]
  assign _GEN_707 = io_sfence_bits_rs2 & _GEN_703; // @[TLB.scala 388:40]
  assign _GEN_708 = io_sfence_bits_rs2 & _GEN_704; // @[TLB.scala 388:40]
  assign _T_615 = _sector_hits_T_27[26:18] == 9'h0; // @[TLB.scala 134:61]
  assign _GEN_729 = sectored_entries_0_4_data_0[13] ? _GEN_513 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_730 = sectored_entries_0_4_data_1[13] ? _GEN_514 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_731 = sectored_entries_0_4_data_2[13] ? _GEN_515 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_732 = sectored_entries_0_4_data_3[13] ? _GEN_516 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_733 = io_sfence_bits_rs2 & _GEN_729; // @[TLB.scala 388:40]
  assign _GEN_734 = io_sfence_bits_rs2 & _GEN_730; // @[TLB.scala 388:40]
  assign _GEN_735 = io_sfence_bits_rs2 & _GEN_731; // @[TLB.scala 388:40]
  assign _GEN_736 = io_sfence_bits_rs2 & _GEN_732; // @[TLB.scala 388:40]
  assign _T_754 = _sector_hits_T_33[26:18] == 9'h0; // @[TLB.scala 134:61]
  assign _GEN_757 = sectored_entries_0_5_data_0[13] ? _GEN_523 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_758 = sectored_entries_0_5_data_1[13] ? _GEN_524 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_759 = sectored_entries_0_5_data_2[13] ? _GEN_525 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_760 = sectored_entries_0_5_data_3[13] ? _GEN_526 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_761 = io_sfence_bits_rs2 & _GEN_757; // @[TLB.scala 388:40]
  assign _GEN_762 = io_sfence_bits_rs2 & _GEN_758; // @[TLB.scala 388:40]
  assign _GEN_763 = io_sfence_bits_rs2 & _GEN_759; // @[TLB.scala 388:40]
  assign _GEN_764 = io_sfence_bits_rs2 & _GEN_760; // @[TLB.scala 388:40]
  assign _T_893 = _sector_hits_T_39[26:18] == 9'h0; // @[TLB.scala 134:61]
  assign _GEN_785 = sectored_entries_0_6_data_0[13] ? _GEN_533 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_786 = sectored_entries_0_6_data_1[13] ? _GEN_534 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_787 = sectored_entries_0_6_data_2[13] ? _GEN_535 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_788 = sectored_entries_0_6_data_3[13] ? _GEN_536 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_789 = io_sfence_bits_rs2 & _GEN_785; // @[TLB.scala 388:40]
  assign _GEN_790 = io_sfence_bits_rs2 & _GEN_786; // @[TLB.scala 388:40]
  assign _GEN_791 = io_sfence_bits_rs2 & _GEN_787; // @[TLB.scala 388:40]
  assign _GEN_792 = io_sfence_bits_rs2 & _GEN_788; // @[TLB.scala 388:40]
  assign _T_1032 = _sector_hits_T_45[26:18] == 9'h0; // @[TLB.scala 134:61]
  assign _GEN_813 = sectored_entries_0_7_data_0[13] ? _GEN_543 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_814 = sectored_entries_0_7_data_1[13] ? _GEN_544 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_815 = sectored_entries_0_7_data_2[13] ? _GEN_545 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_816 = sectored_entries_0_7_data_3[13] ? _GEN_546 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_817 = io_sfence_bits_rs2 & _GEN_813; // @[TLB.scala 388:40]
  assign _GEN_818 = io_sfence_bits_rs2 & _GEN_814; // @[TLB.scala 388:40]
  assign _GEN_819 = io_sfence_bits_rs2 & _GEN_815; // @[TLB.scala 388:40]
  assign _GEN_820 = io_sfence_bits_rs2 & _GEN_816; // @[TLB.scala 388:40]
  assign _GEN_826 = superpage_entries_0_data_0[13] ? _GEN_459 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_827 = io_sfence_bits_rs2 & _GEN_826; // @[TLB.scala 388:40]
  assign _GEN_830 = superpage_entries_1_data_0[13] ? _GEN_463 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_831 = io_sfence_bits_rs2 & _GEN_830; // @[TLB.scala 388:40]
  assign _GEN_834 = superpage_entries_2_data_0[13] ? _GEN_467 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_835 = io_sfence_bits_rs2 & _GEN_834; // @[TLB.scala 388:40]
  assign _GEN_838 = superpage_entries_3_data_0[13] ? _GEN_471 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_839 = io_sfence_bits_rs2 & _GEN_838; // @[TLB.scala 388:40]
  assign _GEN_842 = special_entry_data_0[13] ? _GEN_455 : 1'h0; // @[TLB.scala 142:19]
  assign _GEN_843 = io_sfence_bits_rs2 & _GEN_842; // @[TLB.scala 388:40]
  assign _T_1326 = multipleHits | reset; // @[TLB.scala 392:24]
  assign io_req_ready = state == 2'h0; // @[TLB.scala 341:16]
  assign io_resp_miss = _io_resp_miss_T | multipleHits; // @[TLB.scala 354:16]
  assign io_resp_paddr = {ppn,mpu_physaddr_lo}; // @[TLB.scala 355:17]
  assign io_resp_pf_inst = bad_va | _io_resp_pf_inst_T_1; // @[TLB.scala 344:19]
  assign io_resp_ae_inst = |_io_resp_ae_inst_T_1; // @[TLB.scala 347:19]
  assign io_resp_cacheable = |_io_resp_cacheable_T; // @[TLB.scala 351:21]
  assign io_ptw_req_valid = state == 2'h1; // @[TLB.scala 357:20]
  assign io_ptw_req_bits_valid = ~io_kill; // @[TLB.scala 358:25]
  assign io_ptw_req_bits_bits_addr = r_refill_tag; // @[TLB.scala 359:29]
  assign mpu_ppn_barrier_io_x_ppn = special_entry_data_0[34:15]; // @[package.scala 266:18]
  assign mpu_ppn_barrier_io_x_u = special_entry_data_0[14]; // @[package.scala 266:18]
  assign mpu_ppn_barrier_io_x_ae = special_entry_data_0[12]; // @[package.scala 266:18]
  assign mpu_ppn_barrier_io_x_sw = special_entry_data_0[11]; // @[package.scala 266:18]
  assign mpu_ppn_barrier_io_x_sx = special_entry_data_0[10]; // @[package.scala 266:18]
  assign mpu_ppn_barrier_io_x_sr = special_entry_data_0[9]; // @[package.scala 266:18]
  assign mpu_ppn_barrier_io_x_pw = special_entry_data_0[8]; // @[package.scala 266:18]
  assign mpu_ppn_barrier_io_x_px = special_entry_data_0[7]; // @[package.scala 266:18]
  assign mpu_ppn_barrier_io_x_pr = special_entry_data_0[6]; // @[package.scala 266:18]
  assign mpu_ppn_barrier_io_x_ppp = special_entry_data_0[5]; // @[package.scala 266:18]
  assign mpu_ppn_barrier_io_x_pal = special_entry_data_0[4]; // @[package.scala 266:18]
  assign mpu_ppn_barrier_io_x_paa = special_entry_data_0[3]; // @[package.scala 266:18]
  assign mpu_ppn_barrier_io_x_eff = special_entry_data_0[2]; // @[package.scala 266:18]
  assign mpu_ppn_barrier_io_x_c = special_entry_data_0[1]; // @[package.scala 266:18]
  assign pmp_io_prv = mpu_priv[1:0]; // @[TLB.scala 196:14]
  assign pmp_io_pmp_0_cfg_l = io_ptw_pmp_0_cfg_l; // @[TLB.scala 195:14]
  assign pmp_io_pmp_0_cfg_a = io_ptw_pmp_0_cfg_a; // @[TLB.scala 195:14]
  assign pmp_io_pmp_0_cfg_x = io_ptw_pmp_0_cfg_x; // @[TLB.scala 195:14]
  assign pmp_io_pmp_0_cfg_w = io_ptw_pmp_0_cfg_w; // @[TLB.scala 195:14]
  assign pmp_io_pmp_0_cfg_r = io_ptw_pmp_0_cfg_r; // @[TLB.scala 195:14]
  assign pmp_io_pmp_0_addr = io_ptw_pmp_0_addr; // @[TLB.scala 195:14]
  assign pmp_io_pmp_0_mask = io_ptw_pmp_0_mask; // @[TLB.scala 195:14]
  assign pmp_io_pmp_1_cfg_l = io_ptw_pmp_1_cfg_l; // @[TLB.scala 195:14]
  assign pmp_io_pmp_1_cfg_a = io_ptw_pmp_1_cfg_a; // @[TLB.scala 195:14]
  assign pmp_io_pmp_1_cfg_x = io_ptw_pmp_1_cfg_x; // @[TLB.scala 195:14]
  assign pmp_io_pmp_1_cfg_w = io_ptw_pmp_1_cfg_w; // @[TLB.scala 195:14]
  assign pmp_io_pmp_1_cfg_r = io_ptw_pmp_1_cfg_r; // @[TLB.scala 195:14]
  assign pmp_io_pmp_1_addr = io_ptw_pmp_1_addr; // @[TLB.scala 195:14]
  assign pmp_io_pmp_1_mask = io_ptw_pmp_1_mask; // @[TLB.scala 195:14]
  assign pmp_io_pmp_2_cfg_l = io_ptw_pmp_2_cfg_l; // @[TLB.scala 195:14]
  assign pmp_io_pmp_2_cfg_a = io_ptw_pmp_2_cfg_a; // @[TLB.scala 195:14]
  assign pmp_io_pmp_2_cfg_x = io_ptw_pmp_2_cfg_x; // @[TLB.scala 195:14]
  assign pmp_io_pmp_2_cfg_w = io_ptw_pmp_2_cfg_w; // @[TLB.scala 195:14]
  assign pmp_io_pmp_2_cfg_r = io_ptw_pmp_2_cfg_r; // @[TLB.scala 195:14]
  assign pmp_io_pmp_2_addr = io_ptw_pmp_2_addr; // @[TLB.scala 195:14]
  assign pmp_io_pmp_2_mask = io_ptw_pmp_2_mask; // @[TLB.scala 195:14]
  assign pmp_io_pmp_3_cfg_l = io_ptw_pmp_3_cfg_l; // @[TLB.scala 195:14]
  assign pmp_io_pmp_3_cfg_a = io_ptw_pmp_3_cfg_a; // @[TLB.scala 195:14]
  assign pmp_io_pmp_3_cfg_x = io_ptw_pmp_3_cfg_x; // @[TLB.scala 195:14]
  assign pmp_io_pmp_3_cfg_w = io_ptw_pmp_3_cfg_w; // @[TLB.scala 195:14]
  assign pmp_io_pmp_3_cfg_r = io_ptw_pmp_3_cfg_r; // @[TLB.scala 195:14]
  assign pmp_io_pmp_3_addr = io_ptw_pmp_3_addr; // @[TLB.scala 195:14]
  assign pmp_io_pmp_3_mask = io_ptw_pmp_3_mask; // @[TLB.scala 195:14]
  assign pmp_io_pmp_4_cfg_l = io_ptw_pmp_4_cfg_l; // @[TLB.scala 195:14]
  assign pmp_io_pmp_4_cfg_a = io_ptw_pmp_4_cfg_a; // @[TLB.scala 195:14]
  assign pmp_io_pmp_4_cfg_x = io_ptw_pmp_4_cfg_x; // @[TLB.scala 195:14]
  assign pmp_io_pmp_4_cfg_w = io_ptw_pmp_4_cfg_w; // @[TLB.scala 195:14]
  assign pmp_io_pmp_4_cfg_r = io_ptw_pmp_4_cfg_r; // @[TLB.scala 195:14]
  assign pmp_io_pmp_4_addr = io_ptw_pmp_4_addr; // @[TLB.scala 195:14]
  assign pmp_io_pmp_4_mask = io_ptw_pmp_4_mask; // @[TLB.scala 195:14]
  assign pmp_io_pmp_5_cfg_l = io_ptw_pmp_5_cfg_l; // @[TLB.scala 195:14]
  assign pmp_io_pmp_5_cfg_a = io_ptw_pmp_5_cfg_a; // @[TLB.scala 195:14]
  assign pmp_io_pmp_5_cfg_x = io_ptw_pmp_5_cfg_x; // @[TLB.scala 195:14]
  assign pmp_io_pmp_5_cfg_w = io_ptw_pmp_5_cfg_w; // @[TLB.scala 195:14]
  assign pmp_io_pmp_5_cfg_r = io_ptw_pmp_5_cfg_r; // @[TLB.scala 195:14]
  assign pmp_io_pmp_5_addr = io_ptw_pmp_5_addr; // @[TLB.scala 195:14]
  assign pmp_io_pmp_5_mask = io_ptw_pmp_5_mask; // @[TLB.scala 195:14]
  assign pmp_io_pmp_6_cfg_l = io_ptw_pmp_6_cfg_l; // @[TLB.scala 195:14]
  assign pmp_io_pmp_6_cfg_a = io_ptw_pmp_6_cfg_a; // @[TLB.scala 195:14]
  assign pmp_io_pmp_6_cfg_x = io_ptw_pmp_6_cfg_x; // @[TLB.scala 195:14]
  assign pmp_io_pmp_6_cfg_w = io_ptw_pmp_6_cfg_w; // @[TLB.scala 195:14]
  assign pmp_io_pmp_6_cfg_r = io_ptw_pmp_6_cfg_r; // @[TLB.scala 195:14]
  assign pmp_io_pmp_6_addr = io_ptw_pmp_6_addr; // @[TLB.scala 195:14]
  assign pmp_io_pmp_6_mask = io_ptw_pmp_6_mask; // @[TLB.scala 195:14]
  assign pmp_io_pmp_7_cfg_l = io_ptw_pmp_7_cfg_l; // @[TLB.scala 195:14]
  assign pmp_io_pmp_7_cfg_a = io_ptw_pmp_7_cfg_a; // @[TLB.scala 195:14]
  assign pmp_io_pmp_7_cfg_x = io_ptw_pmp_7_cfg_x; // @[TLB.scala 195:14]
  assign pmp_io_pmp_7_cfg_w = io_ptw_pmp_7_cfg_w; // @[TLB.scala 195:14]
  assign pmp_io_pmp_7_cfg_r = io_ptw_pmp_7_cfg_r; // @[TLB.scala 195:14]
  assign pmp_io_pmp_7_addr = io_ptw_pmp_7_addr; // @[TLB.scala 195:14]
  assign pmp_io_pmp_7_mask = io_ptw_pmp_7_mask; // @[TLB.scala 195:14]
  assign pmp_io_addr = mpu_physaddr[31:0]; // @[TLB.scala 193:15]
  assign entries_barrier_io_x_ppn = _GEN_556[34:15]; // @[package.scala 266:18]
  assign entries_barrier_io_x_u = _GEN_556[14]; // @[package.scala 266:18]
  assign entries_barrier_io_x_ae = _GEN_556[12]; // @[package.scala 266:18]
  assign entries_barrier_io_x_sw = _GEN_556[11]; // @[package.scala 266:18]
  assign entries_barrier_io_x_sx = _GEN_556[10]; // @[package.scala 266:18]
  assign entries_barrier_io_x_sr = _GEN_556[9]; // @[package.scala 266:18]
  assign entries_barrier_io_x_pw = _GEN_556[8]; // @[package.scala 266:18]
  assign entries_barrier_io_x_px = _GEN_556[7]; // @[package.scala 266:18]
  assign entries_barrier_io_x_pr = _GEN_556[6]; // @[package.scala 266:18]
  assign entries_barrier_io_x_ppp = _GEN_556[5]; // @[package.scala 266:18]
  assign entries_barrier_io_x_pal = _GEN_556[4]; // @[package.scala 266:18]
  assign entries_barrier_io_x_paa = _GEN_556[3]; // @[package.scala 266:18]
  assign entries_barrier_io_x_eff = _GEN_556[2]; // @[package.scala 266:18]
  assign entries_barrier_io_x_c = _GEN_556[1]; // @[package.scala 266:18]
  assign entries_barrier_1_io_x_ppn = _GEN_560[34:15]; // @[package.scala 266:18]
  assign entries_barrier_1_io_x_u = _GEN_560[14]; // @[package.scala 266:18]
  assign entries_barrier_1_io_x_ae = _GEN_560[12]; // @[package.scala 266:18]
  assign entries_barrier_1_io_x_sw = _GEN_560[11]; // @[package.scala 266:18]
  assign entries_barrier_1_io_x_sx = _GEN_560[10]; // @[package.scala 266:18]
  assign entries_barrier_1_io_x_sr = _GEN_560[9]; // @[package.scala 266:18]
  assign entries_barrier_1_io_x_pw = _GEN_560[8]; // @[package.scala 266:18]
  assign entries_barrier_1_io_x_px = _GEN_560[7]; // @[package.scala 266:18]
  assign entries_barrier_1_io_x_pr = _GEN_560[6]; // @[package.scala 266:18]
  assign entries_barrier_1_io_x_ppp = _GEN_560[5]; // @[package.scala 266:18]
  assign entries_barrier_1_io_x_pal = _GEN_560[4]; // @[package.scala 266:18]
  assign entries_barrier_1_io_x_paa = _GEN_560[3]; // @[package.scala 266:18]
  assign entries_barrier_1_io_x_eff = _GEN_560[2]; // @[package.scala 266:18]
  assign entries_barrier_1_io_x_c = _GEN_560[1]; // @[package.scala 266:18]
  assign entries_barrier_2_io_x_ppn = _GEN_564[34:15]; // @[package.scala 266:18]
  assign entries_barrier_2_io_x_u = _GEN_564[14]; // @[package.scala 266:18]
  assign entries_barrier_2_io_x_ae = _GEN_564[12]; // @[package.scala 266:18]
  assign entries_barrier_2_io_x_sw = _GEN_564[11]; // @[package.scala 266:18]
  assign entries_barrier_2_io_x_sx = _GEN_564[10]; // @[package.scala 266:18]
  assign entries_barrier_2_io_x_sr = _GEN_564[9]; // @[package.scala 266:18]
  assign entries_barrier_2_io_x_pw = _GEN_564[8]; // @[package.scala 266:18]
  assign entries_barrier_2_io_x_px = _GEN_564[7]; // @[package.scala 266:18]
  assign entries_barrier_2_io_x_pr = _GEN_564[6]; // @[package.scala 266:18]
  assign entries_barrier_2_io_x_ppp = _GEN_564[5]; // @[package.scala 266:18]
  assign entries_barrier_2_io_x_pal = _GEN_564[4]; // @[package.scala 266:18]
  assign entries_barrier_2_io_x_paa = _GEN_564[3]; // @[package.scala 266:18]
  assign entries_barrier_2_io_x_eff = _GEN_564[2]; // @[package.scala 266:18]
  assign entries_barrier_2_io_x_c = _GEN_564[1]; // @[package.scala 266:18]
  assign entries_barrier_3_io_x_ppn = _GEN_568[34:15]; // @[package.scala 266:18]
  assign entries_barrier_3_io_x_u = _GEN_568[14]; // @[package.scala 266:18]
  assign entries_barrier_3_io_x_ae = _GEN_568[12]; // @[package.scala 266:18]
  assign entries_barrier_3_io_x_sw = _GEN_568[11]; // @[package.scala 266:18]
  assign entries_barrier_3_io_x_sx = _GEN_568[10]; // @[package.scala 266:18]
  assign entries_barrier_3_io_x_sr = _GEN_568[9]; // @[package.scala 266:18]
  assign entries_barrier_3_io_x_pw = _GEN_568[8]; // @[package.scala 266:18]
  assign entries_barrier_3_io_x_px = _GEN_568[7]; // @[package.scala 266:18]
  assign entries_barrier_3_io_x_pr = _GEN_568[6]; // @[package.scala 266:18]
  assign entries_barrier_3_io_x_ppp = _GEN_568[5]; // @[package.scala 266:18]
  assign entries_barrier_3_io_x_pal = _GEN_568[4]; // @[package.scala 266:18]
  assign entries_barrier_3_io_x_paa = _GEN_568[3]; // @[package.scala 266:18]
  assign entries_barrier_3_io_x_eff = _GEN_568[2]; // @[package.scala 266:18]
  assign entries_barrier_3_io_x_c = _GEN_568[1]; // @[package.scala 266:18]
  assign entries_barrier_4_io_x_ppn = _GEN_572[34:15]; // @[package.scala 266:18]
  assign entries_barrier_4_io_x_u = _GEN_572[14]; // @[package.scala 266:18]
  assign entries_barrier_4_io_x_ae = _GEN_572[12]; // @[package.scala 266:18]
  assign entries_barrier_4_io_x_sw = _GEN_572[11]; // @[package.scala 266:18]
  assign entries_barrier_4_io_x_sx = _GEN_572[10]; // @[package.scala 266:18]
  assign entries_barrier_4_io_x_sr = _GEN_572[9]; // @[package.scala 266:18]
  assign entries_barrier_4_io_x_pw = _GEN_572[8]; // @[package.scala 266:18]
  assign entries_barrier_4_io_x_px = _GEN_572[7]; // @[package.scala 266:18]
  assign entries_barrier_4_io_x_pr = _GEN_572[6]; // @[package.scala 266:18]
  assign entries_barrier_4_io_x_ppp = _GEN_572[5]; // @[package.scala 266:18]
  assign entries_barrier_4_io_x_pal = _GEN_572[4]; // @[package.scala 266:18]
  assign entries_barrier_4_io_x_paa = _GEN_572[3]; // @[package.scala 266:18]
  assign entries_barrier_4_io_x_eff = _GEN_572[2]; // @[package.scala 266:18]
  assign entries_barrier_4_io_x_c = _GEN_572[1]; // @[package.scala 266:18]
  assign entries_barrier_5_io_x_ppn = _GEN_576[34:15]; // @[package.scala 266:18]
  assign entries_barrier_5_io_x_u = _GEN_576[14]; // @[package.scala 266:18]
  assign entries_barrier_5_io_x_ae = _GEN_576[12]; // @[package.scala 266:18]
  assign entries_barrier_5_io_x_sw = _GEN_576[11]; // @[package.scala 266:18]
  assign entries_barrier_5_io_x_sx = _GEN_576[10]; // @[package.scala 266:18]
  assign entries_barrier_5_io_x_sr = _GEN_576[9]; // @[package.scala 266:18]
  assign entries_barrier_5_io_x_pw = _GEN_576[8]; // @[package.scala 266:18]
  assign entries_barrier_5_io_x_px = _GEN_576[7]; // @[package.scala 266:18]
  assign entries_barrier_5_io_x_pr = _GEN_576[6]; // @[package.scala 266:18]
  assign entries_barrier_5_io_x_ppp = _GEN_576[5]; // @[package.scala 266:18]
  assign entries_barrier_5_io_x_pal = _GEN_576[4]; // @[package.scala 266:18]
  assign entries_barrier_5_io_x_paa = _GEN_576[3]; // @[package.scala 266:18]
  assign entries_barrier_5_io_x_eff = _GEN_576[2]; // @[package.scala 266:18]
  assign entries_barrier_5_io_x_c = _GEN_576[1]; // @[package.scala 266:18]
  assign entries_barrier_6_io_x_ppn = _GEN_580[34:15]; // @[package.scala 266:18]
  assign entries_barrier_6_io_x_u = _GEN_580[14]; // @[package.scala 266:18]
  assign entries_barrier_6_io_x_ae = _GEN_580[12]; // @[package.scala 266:18]
  assign entries_barrier_6_io_x_sw = _GEN_580[11]; // @[package.scala 266:18]
  assign entries_barrier_6_io_x_sx = _GEN_580[10]; // @[package.scala 266:18]
  assign entries_barrier_6_io_x_sr = _GEN_580[9]; // @[package.scala 266:18]
  assign entries_barrier_6_io_x_pw = _GEN_580[8]; // @[package.scala 266:18]
  assign entries_barrier_6_io_x_px = _GEN_580[7]; // @[package.scala 266:18]
  assign entries_barrier_6_io_x_pr = _GEN_580[6]; // @[package.scala 266:18]
  assign entries_barrier_6_io_x_ppp = _GEN_580[5]; // @[package.scala 266:18]
  assign entries_barrier_6_io_x_pal = _GEN_580[4]; // @[package.scala 266:18]
  assign entries_barrier_6_io_x_paa = _GEN_580[3]; // @[package.scala 266:18]
  assign entries_barrier_6_io_x_eff = _GEN_580[2]; // @[package.scala 266:18]
  assign entries_barrier_6_io_x_c = _GEN_580[1]; // @[package.scala 266:18]
  assign entries_barrier_7_io_x_ppn = _GEN_584[34:15]; // @[package.scala 266:18]
  assign entries_barrier_7_io_x_u = _GEN_584[14]; // @[package.scala 266:18]
  assign entries_barrier_7_io_x_ae = _GEN_584[12]; // @[package.scala 266:18]
  assign entries_barrier_7_io_x_sw = _GEN_584[11]; // @[package.scala 266:18]
  assign entries_barrier_7_io_x_sx = _GEN_584[10]; // @[package.scala 266:18]
  assign entries_barrier_7_io_x_sr = _GEN_584[9]; // @[package.scala 266:18]
  assign entries_barrier_7_io_x_pw = _GEN_584[8]; // @[package.scala 266:18]
  assign entries_barrier_7_io_x_px = _GEN_584[7]; // @[package.scala 266:18]
  assign entries_barrier_7_io_x_pr = _GEN_584[6]; // @[package.scala 266:18]
  assign entries_barrier_7_io_x_ppp = _GEN_584[5]; // @[package.scala 266:18]
  assign entries_barrier_7_io_x_pal = _GEN_584[4]; // @[package.scala 266:18]
  assign entries_barrier_7_io_x_paa = _GEN_584[3]; // @[package.scala 266:18]
  assign entries_barrier_7_io_x_eff = _GEN_584[2]; // @[package.scala 266:18]
  assign entries_barrier_7_io_x_c = _GEN_584[1]; // @[package.scala 266:18]
  assign entries_barrier_8_io_x_ppn = superpage_entries_0_data_0[34:15]; // @[package.scala 266:18]
  assign entries_barrier_8_io_x_u = superpage_entries_0_data_0[14]; // @[package.scala 266:18]
  assign entries_barrier_8_io_x_ae = superpage_entries_0_data_0[12]; // @[package.scala 266:18]
  assign entries_barrier_8_io_x_sw = superpage_entries_0_data_0[11]; // @[package.scala 266:18]
  assign entries_barrier_8_io_x_sx = superpage_entries_0_data_0[10]; // @[package.scala 266:18]
  assign entries_barrier_8_io_x_sr = superpage_entries_0_data_0[9]; // @[package.scala 266:18]
  assign entries_barrier_8_io_x_pw = superpage_entries_0_data_0[8]; // @[package.scala 266:18]
  assign entries_barrier_8_io_x_px = superpage_entries_0_data_0[7]; // @[package.scala 266:18]
  assign entries_barrier_8_io_x_pr = superpage_entries_0_data_0[6]; // @[package.scala 266:18]
  assign entries_barrier_8_io_x_ppp = superpage_entries_0_data_0[5]; // @[package.scala 266:18]
  assign entries_barrier_8_io_x_pal = superpage_entries_0_data_0[4]; // @[package.scala 266:18]
  assign entries_barrier_8_io_x_paa = superpage_entries_0_data_0[3]; // @[package.scala 266:18]
  assign entries_barrier_8_io_x_eff = superpage_entries_0_data_0[2]; // @[package.scala 266:18]
  assign entries_barrier_8_io_x_c = superpage_entries_0_data_0[1]; // @[package.scala 266:18]
  assign entries_barrier_9_io_x_ppn = superpage_entries_1_data_0[34:15]; // @[package.scala 266:18]
  assign entries_barrier_9_io_x_u = superpage_entries_1_data_0[14]; // @[package.scala 266:18]
  assign entries_barrier_9_io_x_ae = superpage_entries_1_data_0[12]; // @[package.scala 266:18]
  assign entries_barrier_9_io_x_sw = superpage_entries_1_data_0[11]; // @[package.scala 266:18]
  assign entries_barrier_9_io_x_sx = superpage_entries_1_data_0[10]; // @[package.scala 266:18]
  assign entries_barrier_9_io_x_sr = superpage_entries_1_data_0[9]; // @[package.scala 266:18]
  assign entries_barrier_9_io_x_pw = superpage_entries_1_data_0[8]; // @[package.scala 266:18]
  assign entries_barrier_9_io_x_px = superpage_entries_1_data_0[7]; // @[package.scala 266:18]
  assign entries_barrier_9_io_x_pr = superpage_entries_1_data_0[6]; // @[package.scala 266:18]
  assign entries_barrier_9_io_x_ppp = superpage_entries_1_data_0[5]; // @[package.scala 266:18]
  assign entries_barrier_9_io_x_pal = superpage_entries_1_data_0[4]; // @[package.scala 266:18]
  assign entries_barrier_9_io_x_paa = superpage_entries_1_data_0[3]; // @[package.scala 266:18]
  assign entries_barrier_9_io_x_eff = superpage_entries_1_data_0[2]; // @[package.scala 266:18]
  assign entries_barrier_9_io_x_c = superpage_entries_1_data_0[1]; // @[package.scala 266:18]
  assign entries_barrier_10_io_x_ppn = superpage_entries_2_data_0[34:15]; // @[package.scala 266:18]
  assign entries_barrier_10_io_x_u = superpage_entries_2_data_0[14]; // @[package.scala 266:18]
  assign entries_barrier_10_io_x_ae = superpage_entries_2_data_0[12]; // @[package.scala 266:18]
  assign entries_barrier_10_io_x_sw = superpage_entries_2_data_0[11]; // @[package.scala 266:18]
  assign entries_barrier_10_io_x_sx = superpage_entries_2_data_0[10]; // @[package.scala 266:18]
  assign entries_barrier_10_io_x_sr = superpage_entries_2_data_0[9]; // @[package.scala 266:18]
  assign entries_barrier_10_io_x_pw = superpage_entries_2_data_0[8]; // @[package.scala 266:18]
  assign entries_barrier_10_io_x_px = superpage_entries_2_data_0[7]; // @[package.scala 266:18]
  assign entries_barrier_10_io_x_pr = superpage_entries_2_data_0[6]; // @[package.scala 266:18]
  assign entries_barrier_10_io_x_ppp = superpage_entries_2_data_0[5]; // @[package.scala 266:18]
  assign entries_barrier_10_io_x_pal = superpage_entries_2_data_0[4]; // @[package.scala 266:18]
  assign entries_barrier_10_io_x_paa = superpage_entries_2_data_0[3]; // @[package.scala 266:18]
  assign entries_barrier_10_io_x_eff = superpage_entries_2_data_0[2]; // @[package.scala 266:18]
  assign entries_barrier_10_io_x_c = superpage_entries_2_data_0[1]; // @[package.scala 266:18]
  assign entries_barrier_11_io_x_ppn = superpage_entries_3_data_0[34:15]; // @[package.scala 266:18]
  assign entries_barrier_11_io_x_u = superpage_entries_3_data_0[14]; // @[package.scala 266:18]
  assign entries_barrier_11_io_x_ae = superpage_entries_3_data_0[12]; // @[package.scala 266:18]
  assign entries_barrier_11_io_x_sw = superpage_entries_3_data_0[11]; // @[package.scala 266:18]
  assign entries_barrier_11_io_x_sx = superpage_entries_3_data_0[10]; // @[package.scala 266:18]
  assign entries_barrier_11_io_x_sr = superpage_entries_3_data_0[9]; // @[package.scala 266:18]
  assign entries_barrier_11_io_x_pw = superpage_entries_3_data_0[8]; // @[package.scala 266:18]
  assign entries_barrier_11_io_x_px = superpage_entries_3_data_0[7]; // @[package.scala 266:18]
  assign entries_barrier_11_io_x_pr = superpage_entries_3_data_0[6]; // @[package.scala 266:18]
  assign entries_barrier_11_io_x_ppp = superpage_entries_3_data_0[5]; // @[package.scala 266:18]
  assign entries_barrier_11_io_x_pal = superpage_entries_3_data_0[4]; // @[package.scala 266:18]
  assign entries_barrier_11_io_x_paa = superpage_entries_3_data_0[3]; // @[package.scala 266:18]
  assign entries_barrier_11_io_x_eff = superpage_entries_3_data_0[2]; // @[package.scala 266:18]
  assign entries_barrier_11_io_x_c = superpage_entries_3_data_0[1]; // @[package.scala 266:18]
  assign entries_barrier_12_io_x_ppn = special_entry_data_0[34:15]; // @[package.scala 266:18]
  assign entries_barrier_12_io_x_u = special_entry_data_0[14]; // @[package.scala 266:18]
  assign entries_barrier_12_io_x_ae = special_entry_data_0[12]; // @[package.scala 266:18]
  assign entries_barrier_12_io_x_sw = special_entry_data_0[11]; // @[package.scala 266:18]
  assign entries_barrier_12_io_x_sx = special_entry_data_0[10]; // @[package.scala 266:18]
  assign entries_barrier_12_io_x_sr = special_entry_data_0[9]; // @[package.scala 266:18]
  assign entries_barrier_12_io_x_pw = special_entry_data_0[8]; // @[package.scala 266:18]
  assign entries_barrier_12_io_x_px = special_entry_data_0[7]; // @[package.scala 266:18]
  assign entries_barrier_12_io_x_pr = special_entry_data_0[6]; // @[package.scala 266:18]
  assign entries_barrier_12_io_x_ppp = special_entry_data_0[5]; // @[package.scala 266:18]
  assign entries_barrier_12_io_x_pal = special_entry_data_0[4]; // @[package.scala 266:18]
  assign entries_barrier_12_io_x_paa = special_entry_data_0[3]; // @[package.scala 266:18]
  assign entries_barrier_12_io_x_eff = special_entry_data_0[2]; // @[package.scala 266:18]
  assign entries_barrier_12_io_x_c = special_entry_data_0[1]; // @[package.scala 266:18]
  assign TLB_1_cov_read_addr = TLB_1_state;
  assign TLB_1_cov_read_data = TLB_1_cov[TLB_1_cov_read_addr]; // @[Coverage map for TLB_1]
  assign TLB_1_cov_write_data = 1'h1;
  assign TLB_1_cov_write_addr = TLB_1_state;
  assign TLB_1_cov_write_mask = 1'h1;
  assign TLB_1_cov_write_en = 1'h1;
  assign mux_cond_0 = sectored_entries_0_6_data_1[0];
  assign mux_cond_1 = sectored_entries_0_7_data_1[0];
  assign mux_cond_2 = ~sectored_entries_0_2_data_0[13];
  assign mux_cond_3 = ~sectored_entries_0_7_data_1[13];
  assign mux_cond_4 = sectored_entries_0_7_data_3[0];
  assign mux_cond_5 = sectored_entries_0_4_data_0[0];
  assign mux_cond_6 = sectored_entries_0_3_data_3[0];
  assign mux_cond_7 = sectored_entries_0_2_data_3[0];
  assign mux_cond_8 = sectored_entries_0_2_data_0[0];
  assign mux_cond_9 = ~sectored_entries_0_6_data_1[13];
  assign mux_cond_10 = ~sectored_entries_0_2_data_2[13];
  assign mux_cond_11 = ~superpage_entries_0_data_0[13];
  assign mux_cond_12 = sectored_entries_0_3_data_1[0];
  assign mux_cond_13 = sectored_entries_0_4_data_3[0];
  assign mux_cond_14 = ~sectored_entries_0_3_data_3[13];
  assign mux_cond_15 = sectored_entries_0_3_data_2[0];
  assign mux_cond_16 = ~sectored_entries_0_4_data_3[13];
  assign mux_cond_17 = ~sectored_entries_0_4_data_0[13];
  assign mux_cond_18 = ~sectored_entries_0_4_data_1[13];
  assign mux_cond_19 = sectored_entries_0_6_data_0[0];
  assign mux_cond_20 = sectored_entries_0_5_data_0[0];
  assign mux_cond_21 = sectored_entries_0_6_data_2[0];
  assign mux_cond_22 = sectored_entries_0_0_data_3[0];
  assign mux_cond_23 = ~sectored_entries_0_3_data_1[13];
  assign mux_cond_24 = ~sectored_entries_0_7_data_0[13];
  assign mux_cond_25 = sectored_entries_0_7_data_0[0];
  assign mux_cond_26 = ~sectored_entries_0_7_data_3[13];
  assign mux_cond_27 = ~sectored_entries_0_0_data_3[13];
  assign mux_cond_28 = ~superpage_entries_1_data_0[13];
  assign mux_cond_29 = ~sectored_entries_0_7_data_2[13];
  assign mux_cond_30 = ~sectored_entries_0_6_data_0[13];
  assign mux_cond_31 = ~sectored_entries_0_6_data_3[13];
  assign mux_cond_32 = sectored_entries_0_2_data_2[0];
  assign mux_cond_33 = sectored_entries_0_1_data_1[0];
  assign mux_cond_34 = ~sectored_entries_0_2_data_1[13];
  assign mux_cond_35 = ~sectored_entries_0_4_data_2[13];
  assign mux_cond_36 = ~sectored_entries_0_1_data_3[13];
  assign mux_cond_37 = ~sectored_entries_0_0_data_2[13];
  assign mux_cond_38 = ~sectored_entries_0_0_data_0[13];
  assign mux_cond_39 = ~sectored_entries_0_2_data_3[13];
  assign mux_cond_40 = sectored_entries_0_7_data_2[0];
  assign mux_cond_41 = sectored_entries_0_0_data_0[0];
  assign mux_cond_42 = ~sectored_entries_0_5_data_0[13];
  assign mux_cond_43 = sectored_entries_0_4_data_1[0];
  assign mux_cond_44 = sectored_entries_0_5_data_1[0];
  assign mux_cond_45 = ~sectored_entries_0_5_data_3[13];
  assign mux_cond_46 = sectored_entries_0_1_data_0[0];
  assign mux_cond_47 = sectored_entries_0_5_data_3[0];
  assign mux_cond_48 = ~sectored_entries_0_0_data_1[13];
  assign mux_cond_49 = ~special_entry_data_0[13];
  assign mux_cond_50 = ~superpage_entries_2_data_0[13];
  assign mux_cond_51 = sectored_entries_0_0_data_2[0];
  assign mux_cond_52 = sectored_entries_0_6_data_3[0];
  assign mux_cond_53 = ~sectored_entries_0_3_data_0[13];
  assign mux_cond_54 = ~sectored_entries_0_1_data_0[13];
  assign mux_cond_55 = sectored_entries_0_1_data_2[0];
  assign mux_cond_56 = ~sectored_entries_0_5_data_2[13];
  assign mux_cond_57 = ~sectored_entries_0_6_data_2[13];
  assign mux_cond_58 = sectored_entries_0_1_data_3[0];
  assign mux_cond_59 = ~sectored_entries_0_3_data_2[13];
  assign mux_cond_60 = ~sectored_entries_0_1_data_1[13];
  assign mux_cond_61 = ~sectored_entries_0_1_data_2[13];
  assign mux_cond_62 = sectored_entries_0_3_data_0[0];
  assign mux_cond_63 = sectored_entries_0_5_data_2[0];
  assign mux_cond_64 = sectored_entries_0_0_data_1[0];
  assign mux_cond_65 = sectored_entries_0_2_data_1[0];
  assign mux_cond_66 = ~sectored_entries_0_5_data_1[13];
  assign mux_cond_67 = ~superpage_entries_3_data_0[13];
  assign mux_cond_68 = sectored_entries_0_4_data_2[0];
  assign r_sectored_hit_shl = r_sectored_hit;
  assign r_sectored_hit_pad = {19'h0,r_sectored_hit_shl};
  assign r_sectored_repl_addr_shl = {r_sectored_repl_addr, 8'h0};
  assign r_sectored_repl_addr_pad = {9'h0,r_sectored_repl_addr_shl};
  assign r_superpage_repl_addr_shl = r_superpage_repl_addr;
  assign r_superpage_repl_addr_pad = {18'h0,r_superpage_repl_addr_shl};
  assign special_entry_valid_0_shl = {special_entry_valid_0, 13'h0};
  assign special_entry_valid_0_pad = {6'h0,special_entry_valid_0_shl};
  assign special_entry_level_shl = {special_entry_level, 12'h0};
  assign special_entry_level_pad = {6'h0,special_entry_level_shl};
  assign state_shl = {state, 12'h0};
  assign state_pad = {6'h0,state_shl};
  assign r_sectored_hit_addr_shl = {r_sectored_hit_addr, 1'h0};
  assign r_sectored_hit_addr_pad = {16'h0,r_sectored_hit_addr_shl};
  assign mux_cond_0_shl = {mux_cond_0, 16'h0};
  assign mux_cond_0_pad = {3'h0,mux_cond_0_shl};
  assign mux_cond_1_shl = {mux_cond_1, 10'h0};
  assign mux_cond_1_pad = {9'h0,mux_cond_1_shl};
  assign mux_cond_2_shl = {mux_cond_2, 2'h0};
  assign mux_cond_2_pad = {17'h0,mux_cond_2_shl};
  assign mux_cond_3_shl = {mux_cond_3, 15'h0};
  assign mux_cond_3_pad = {4'h0,mux_cond_3_shl};
  assign mux_cond_4_shl = {mux_cond_4, 4'h0};
  assign mux_cond_4_pad = {15'h0,mux_cond_4_shl};
  assign mux_cond_5_shl = {mux_cond_5, 13'h0};
  assign mux_cond_5_pad = {6'h0,mux_cond_5_shl};
  assign mux_cond_6_shl = {mux_cond_6, 9'h0};
  assign mux_cond_6_pad = {10'h0,mux_cond_6_shl};
  assign mux_cond_7_shl = {mux_cond_7, 8'h0};
  assign mux_cond_7_pad = {11'h0,mux_cond_7_shl};
  assign mux_cond_8_shl = {mux_cond_8, 12'h0};
  assign mux_cond_8_pad = {7'h0,mux_cond_8_shl};
  assign mux_cond_9_shl = {mux_cond_9, 19'h0};
  assign mux_cond_9_pad = mux_cond_9_shl;
  assign mux_cond_10_shl = {mux_cond_10, 18'h0};
  assign mux_cond_10_pad = {1'h0,mux_cond_10_shl};
  assign mux_cond_11_shl = {mux_cond_11, 9'h0};
  assign mux_cond_11_pad = {10'h0,mux_cond_11_shl};
  assign mux_cond_12_shl = {mux_cond_12, 19'h0};
  assign mux_cond_12_pad = mux_cond_12_shl;
  assign mux_cond_13_shl = {mux_cond_13, 7'h0};
  assign mux_cond_13_pad = {12'h0,mux_cond_13_shl};
  assign mux_cond_14_shl = {mux_cond_14, 11'h0};
  assign mux_cond_14_pad = {8'h0,mux_cond_14_shl};
  assign mux_cond_15_shl = mux_cond_15;
  assign mux_cond_15_pad = {19'h0,mux_cond_15_shl};
  assign mux_cond_16_shl = {mux_cond_16, 4'h0};
  assign mux_cond_16_pad = {15'h0,mux_cond_16_shl};
  assign mux_cond_17_shl = {mux_cond_17, 19'h0};
  assign mux_cond_17_pad = mux_cond_17_shl;
  assign mux_cond_18_shl = {mux_cond_18, 9'h0};
  assign mux_cond_18_pad = {10'h0,mux_cond_18_shl};
  assign mux_cond_19_shl = {mux_cond_19, 8'h0};
  assign mux_cond_19_pad = {11'h0,mux_cond_19_shl};
  assign mux_cond_20_shl = {mux_cond_20, 4'h0};
  assign mux_cond_20_pad = {15'h0,mux_cond_20_shl};
  assign mux_cond_21_shl = {mux_cond_21, 6'h0};
  assign mux_cond_21_pad = {13'h0,mux_cond_21_shl};
  assign mux_cond_22_shl = {mux_cond_22, 11'h0};
  assign mux_cond_22_pad = {8'h0,mux_cond_22_shl};
  assign mux_cond_23_shl = {mux_cond_23, 14'h0};
  assign mux_cond_23_pad = {5'h0,mux_cond_23_shl};
  assign mux_cond_24_shl = {mux_cond_24, 7'h0};
  assign mux_cond_24_pad = {12'h0,mux_cond_24_shl};
  assign mux_cond_25_shl = {mux_cond_25, 7'h0};
  assign mux_cond_25_pad = {12'h0,mux_cond_25_shl};
  assign mux_cond_26_shl = {mux_cond_26, 19'h0};
  assign mux_cond_26_pad = mux_cond_26_shl;
  assign mux_cond_27_shl = {mux_cond_27, 10'h0};
  assign mux_cond_27_pad = {9'h0,mux_cond_27_shl};
  assign mux_cond_28_shl = {mux_cond_28, 17'h0};
  assign mux_cond_28_pad = {2'h0,mux_cond_28_shl};
  assign mux_cond_29_shl = {mux_cond_29, 3'h0};
  assign mux_cond_29_pad = {16'h0,mux_cond_29_shl};
  assign mux_cond_30_shl = {mux_cond_30, 9'h0};
  assign mux_cond_30_pad = {10'h0,mux_cond_30_shl};
  assign mux_cond_31_shl = {mux_cond_31, 15'h0};
  assign mux_cond_31_pad = {4'h0,mux_cond_31_shl};
  assign mux_cond_32_shl = mux_cond_32;
  assign mux_cond_32_pad = {19'h0,mux_cond_32_shl};
  assign mux_cond_33_shl = {mux_cond_33, 12'h0};
  assign mux_cond_33_pad = {7'h0,mux_cond_33_shl};
  assign mux_cond_34_shl = {mux_cond_34, 17'h0};
  assign mux_cond_34_pad = {2'h0,mux_cond_34_shl};
  assign mux_cond_35_shl = {mux_cond_35, 9'h0};
  assign mux_cond_35_pad = {10'h0,mux_cond_35_shl};
  assign mux_cond_36_shl = {mux_cond_36, 12'h0};
  assign mux_cond_36_pad = {7'h0,mux_cond_36_shl};
  assign mux_cond_37_shl = mux_cond_37;
  assign mux_cond_37_pad = {19'h0,mux_cond_37_shl};
  assign mux_cond_38_shl = {mux_cond_38, 5'h0};
  assign mux_cond_38_pad = {14'h0,mux_cond_38_shl};
  assign mux_cond_39_shl = {mux_cond_39, 2'h0};
  assign mux_cond_39_pad = {17'h0,mux_cond_39_shl};
  assign mux_cond_40_shl = {mux_cond_40, 18'h0};
  assign mux_cond_40_pad = {1'h0,mux_cond_40_shl};
  assign mux_cond_41_shl = {mux_cond_41, 13'h0};
  assign mux_cond_41_pad = {6'h0,mux_cond_41_shl};
  assign mux_cond_42_shl = {mux_cond_42, 5'h0};
  assign mux_cond_42_pad = {14'h0,mux_cond_42_shl};
  assign mux_cond_43_shl = {mux_cond_43, 18'h0};
  assign mux_cond_43_pad = {1'h0,mux_cond_43_shl};
  assign mux_cond_44_shl = {mux_cond_44, 18'h0};
  assign mux_cond_44_pad = {1'h0,mux_cond_44_shl};
  assign mux_cond_45_shl = {mux_cond_45, 2'h0};
  assign mux_cond_45_pad = {17'h0,mux_cond_45_shl};
  assign mux_cond_46_shl = {mux_cond_46, 12'h0};
  assign mux_cond_46_pad = {7'h0,mux_cond_46_shl};
  assign mux_cond_47_shl = {mux_cond_47, 18'h0};
  assign mux_cond_47_pad = {1'h0,mux_cond_47_shl};
  assign mux_cond_48_shl = {mux_cond_48, 16'h0};
  assign mux_cond_48_pad = {3'h0,mux_cond_48_shl};
  assign mux_cond_49_shl = mux_cond_49;
  assign mux_cond_49_pad = {19'h0,mux_cond_49_shl};
  assign mux_cond_50_shl = {mux_cond_50, 4'h0};
  assign mux_cond_50_pad = {15'h0,mux_cond_50_shl};
  assign mux_cond_51_shl = {mux_cond_51, 9'h0};
  assign mux_cond_51_pad = {10'h0,mux_cond_51_shl};
  assign mux_cond_52_shl = {mux_cond_52, 13'h0};
  assign mux_cond_52_pad = {6'h0,mux_cond_52_shl};
  assign mux_cond_53_shl = {mux_cond_53, 4'h0};
  assign mux_cond_53_pad = {15'h0,mux_cond_53_shl};
  assign mux_cond_54_shl = {mux_cond_54, 5'h0};
  assign mux_cond_54_pad = {14'h0,mux_cond_54_shl};
  assign mux_cond_55_shl = {mux_cond_55, 10'h0};
  assign mux_cond_55_pad = {9'h0,mux_cond_55_shl};
  assign mux_cond_56_shl = {mux_cond_56, 12'h0};
  assign mux_cond_56_pad = {7'h0,mux_cond_56_shl};
  assign mux_cond_57_shl = {mux_cond_57, 4'h0};
  assign mux_cond_57_pad = {15'h0,mux_cond_57_shl};
  assign mux_cond_58_shl = {mux_cond_58, 19'h0};
  assign mux_cond_58_pad = mux_cond_58_shl;
  assign mux_cond_59_shl = {mux_cond_59, 8'h0};
  assign mux_cond_59_pad = {11'h0,mux_cond_59_shl};
  assign mux_cond_60_shl = {mux_cond_60, 12'h0};
  assign mux_cond_60_pad = {7'h0,mux_cond_60_shl};
  assign mux_cond_61_shl = {mux_cond_61, 13'h0};
  assign mux_cond_61_pad = {6'h0,mux_cond_61_shl};
  assign mux_cond_62_shl = {mux_cond_62, 19'h0};
  assign mux_cond_62_pad = mux_cond_62_shl;
  assign mux_cond_63_shl = {mux_cond_63, 7'h0};
  assign mux_cond_63_pad = {12'h0,mux_cond_63_shl};
  assign mux_cond_64_shl = {mux_cond_64, 1'h0};
  assign mux_cond_64_pad = {18'h0,mux_cond_64_shl};
  assign mux_cond_65_shl = {mux_cond_65, 3'h0};
  assign mux_cond_65_pad = {16'h0,mux_cond_65_shl};
  assign mux_cond_66_shl = {mux_cond_66, 1'h0};
  assign mux_cond_66_pad = {18'h0,mux_cond_66_shl};
  assign mux_cond_67_shl = {mux_cond_67, 15'h0};
  assign mux_cond_67_pad = {4'h0,mux_cond_67_shl};
  assign mux_cond_68_shl = {mux_cond_68, 15'h0};
  assign mux_cond_68_pad = {4'h0,mux_cond_68_shl};
  assign sectored_entries_0_0_valid_3_shl = {sectored_entries_0_0_valid_3, 5'h0};
  assign sectored_entries_0_0_valid_3_pad = {14'h0,sectored_entries_0_0_valid_3_shl};
  assign sectored_entries_0_0_valid_2_shl = {sectored_entries_0_0_valid_2, 4'h0};
  assign sectored_entries_0_0_valid_2_pad = {15'h0,sectored_entries_0_0_valid_2_shl};
  assign sectored_entries_0_2_valid_0_shl = {sectored_entries_0_2_valid_0, 5'h0};
  assign sectored_entries_0_2_valid_0_pad = {14'h0,sectored_entries_0_2_valid_0_shl};
  assign sectored_entries_0_3_valid_0_shl = {sectored_entries_0_3_valid_0, 5'h0};
  assign sectored_entries_0_3_valid_0_pad = {14'h0,sectored_entries_0_3_valid_0_shl};
  assign superpage_entries_2_level_shl = {superpage_entries_2_level, 13'h0};
  assign superpage_entries_2_level_pad = {5'h0,superpage_entries_2_level_shl};
  assign sectored_entries_0_7_valid_1_shl = {sectored_entries_0_7_valid_1, 4'h0};
  assign sectored_entries_0_7_valid_1_pad = {15'h0,sectored_entries_0_7_valid_1_shl};
  assign sectored_entries_0_4_valid_0_shl = {sectored_entries_0_4_valid_0, 5'h0};
  assign sectored_entries_0_4_valid_0_pad = {14'h0,sectored_entries_0_4_valid_0_shl};
  assign sectored_entries_0_1_valid_3_shl = {sectored_entries_0_1_valid_3, 5'h0};
  assign sectored_entries_0_1_valid_3_pad = {14'h0,sectored_entries_0_1_valid_3_shl};
  assign sectored_entries_0_1_valid_1_shl = {sectored_entries_0_1_valid_1, 4'h0};
  assign sectored_entries_0_1_valid_1_pad = {15'h0,sectored_entries_0_1_valid_1_shl};
  assign sectored_entries_0_2_valid_3_shl = {sectored_entries_0_2_valid_3, 5'h0};
  assign sectored_entries_0_2_valid_3_pad = {14'h0,sectored_entries_0_2_valid_3_shl};
  assign sectored_entries_0_2_valid_1_shl = {sectored_entries_0_2_valid_1, 4'h0};
  assign sectored_entries_0_2_valid_1_pad = {15'h0,sectored_entries_0_2_valid_1_shl};
  assign superpage_entries_1_valid_0_shl = {superpage_entries_1_valid_0, 1'h0};
  assign superpage_entries_1_valid_0_pad = {18'h0,superpage_entries_1_valid_0_shl};
  assign sectored_entries_0_7_valid_0_shl = {sectored_entries_0_7_valid_0, 5'h0};
  assign sectored_entries_0_7_valid_0_pad = {14'h0,sectored_entries_0_7_valid_0_shl};
  assign superpage_entries_3_valid_0_shl = {superpage_entries_3_valid_0, 1'h0};
  assign superpage_entries_3_valid_0_pad = {18'h0,superpage_entries_3_valid_0_shl};
  assign sectored_entries_0_5_valid_3_shl = {sectored_entries_0_5_valid_3, 5'h0};
  assign sectored_entries_0_5_valid_3_pad = {14'h0,sectored_entries_0_5_valid_3_shl};
  assign sectored_entries_0_5_valid_1_shl = {sectored_entries_0_5_valid_1, 4'h0};
  assign sectored_entries_0_5_valid_1_pad = {15'h0,sectored_entries_0_5_valid_1_shl};
  assign sectored_entries_0_4_valid_3_shl = {sectored_entries_0_4_valid_3, 5'h0};
  assign sectored_entries_0_4_valid_3_pad = {14'h0,sectored_entries_0_4_valid_3_shl};
  assign sectored_entries_0_5_valid_2_shl = {sectored_entries_0_5_valid_2, 4'h0};
  assign sectored_entries_0_5_valid_2_pad = {15'h0,sectored_entries_0_5_valid_2_shl};
  assign sectored_entries_0_1_valid_2_shl = {sectored_entries_0_1_valid_2, 4'h0};
  assign sectored_entries_0_1_valid_2_pad = {15'h0,sectored_entries_0_1_valid_2_shl};
  assign sectored_entries_0_3_valid_1_shl = {sectored_entries_0_3_valid_1, 4'h0};
  assign sectored_entries_0_3_valid_1_pad = {15'h0,sectored_entries_0_3_valid_1_shl};
  assign sectored_entries_0_1_valid_0_shl = {sectored_entries_0_1_valid_0, 5'h0};
  assign sectored_entries_0_1_valid_0_pad = {14'h0,sectored_entries_0_1_valid_0_shl};
  assign sectored_entries_0_4_valid_2_shl = {sectored_entries_0_4_valid_2, 4'h0};
  assign sectored_entries_0_4_valid_2_pad = {15'h0,sectored_entries_0_4_valid_2_shl};
  assign sectored_entries_0_4_valid_1_shl = {sectored_entries_0_4_valid_1, 4'h0};
  assign sectored_entries_0_4_valid_1_pad = {15'h0,sectored_entries_0_4_valid_1_shl};
  assign superpage_entries_3_level_shl = {superpage_entries_3_level, 13'h0};
  assign superpage_entries_3_level_pad = {5'h0,superpage_entries_3_level_shl};
  assign sectored_entries_0_0_valid_1_shl = {sectored_entries_0_0_valid_1, 4'h0};
  assign sectored_entries_0_0_valid_1_pad = {15'h0,sectored_entries_0_0_valid_1_shl};
  assign sectored_entries_0_3_valid_2_shl = {sectored_entries_0_3_valid_2, 4'h0};
  assign sectored_entries_0_3_valid_2_pad = {15'h0,sectored_entries_0_3_valid_2_shl};
  assign sectored_entries_0_6_valid_1_shl = {sectored_entries_0_6_valid_1, 4'h0};
  assign sectored_entries_0_6_valid_1_pad = {15'h0,sectored_entries_0_6_valid_1_shl};
  assign sectored_entries_0_7_valid_3_shl = {sectored_entries_0_7_valid_3, 5'h0};
  assign sectored_entries_0_7_valid_3_pad = {14'h0,sectored_entries_0_7_valid_3_shl};
  assign sectored_entries_0_3_valid_3_shl = {sectored_entries_0_3_valid_3, 5'h0};
  assign sectored_entries_0_3_valid_3_pad = {14'h0,sectored_entries_0_3_valid_3_shl};
  assign sectored_entries_0_0_valid_0_shl = {sectored_entries_0_0_valid_0, 5'h0};
  assign sectored_entries_0_0_valid_0_pad = {14'h0,sectored_entries_0_0_valid_0_shl};
  assign superpage_entries_0_valid_0_shl = {superpage_entries_0_valid_0, 1'h0};
  assign superpage_entries_0_valid_0_pad = {18'h0,superpage_entries_0_valid_0_shl};
  assign sectored_entries_0_2_valid_2_shl = {sectored_entries_0_2_valid_2, 4'h0};
  assign sectored_entries_0_2_valid_2_pad = {15'h0,sectored_entries_0_2_valid_2_shl};
  assign sectored_entries_0_6_valid_2_shl = {sectored_entries_0_6_valid_2, 4'h0};
  assign sectored_entries_0_6_valid_2_pad = {15'h0,sectored_entries_0_6_valid_2_shl};
  assign superpage_entries_2_valid_0_shl = {superpage_entries_2_valid_0, 1'h0};
  assign superpage_entries_2_valid_0_pad = {18'h0,superpage_entries_2_valid_0_shl};
  assign sectored_entries_0_6_valid_3_shl = {sectored_entries_0_6_valid_3, 5'h0};
  assign sectored_entries_0_6_valid_3_pad = {14'h0,sectored_entries_0_6_valid_3_shl};
  assign sectored_entries_0_6_valid_0_shl = {sectored_entries_0_6_valid_0, 5'h0};
  assign sectored_entries_0_6_valid_0_pad = {14'h0,sectored_entries_0_6_valid_0_shl};
  assign sectored_entries_0_7_valid_2_shl = {sectored_entries_0_7_valid_2, 4'h0};
  assign sectored_entries_0_7_valid_2_pad = {15'h0,sectored_entries_0_7_valid_2_shl};
  assign superpage_entries_0_level_shl = {superpage_entries_0_level, 13'h0};
  assign superpage_entries_0_level_pad = {5'h0,superpage_entries_0_level_shl};
  assign superpage_entries_1_level_shl = {superpage_entries_1_level, 13'h0};
  assign superpage_entries_1_level_pad = {5'h0,superpage_entries_1_level_shl};
  assign sectored_entries_0_5_valid_0_shl = {sectored_entries_0_5_valid_0, 5'h0};
  assign sectored_entries_0_5_valid_0_pad = {14'h0,sectored_entries_0_5_valid_0_shl};
  assign TLB_1_xor64 = r_sectored_repl_addr_pad ^ r_superpage_repl_addr_pad;
  assign TLB_1_xor31 = r_sectored_hit_pad ^ TLB_1_xor64;
  assign TLB_1_xor65 = special_entry_valid_0_pad ^ special_entry_level_pad;
  assign TLB_1_xor66 = state_pad ^ r_sectored_hit_addr_pad;
  assign TLB_1_xor32 = TLB_1_xor65 ^ TLB_1_xor66;
  assign TLB_1_xor15 = TLB_1_xor31 ^ TLB_1_xor32;
  assign TLB_1_xor68 = mux_cond_1_pad ^ mux_cond_2_pad;
  assign TLB_1_xor33 = mux_cond_0_pad ^ TLB_1_xor68;
  assign TLB_1_xor69 = mux_cond_3_pad ^ mux_cond_4_pad;
  assign TLB_1_xor70 = mux_cond_5_pad ^ mux_cond_6_pad;
  assign TLB_1_xor34 = TLB_1_xor69 ^ TLB_1_xor70;
  assign TLB_1_xor16 = TLB_1_xor33 ^ TLB_1_xor34;
  assign TLB_1_xor7 = TLB_1_xor15 ^ TLB_1_xor16;
  assign TLB_1_xor72 = mux_cond_8_pad ^ mux_cond_9_pad;
  assign TLB_1_xor35 = mux_cond_7_pad ^ TLB_1_xor72;
  assign TLB_1_xor73 = mux_cond_10_pad ^ mux_cond_11_pad;
  assign TLB_1_xor74 = mux_cond_12_pad ^ mux_cond_13_pad;
  assign TLB_1_xor36 = TLB_1_xor73 ^ TLB_1_xor74;
  assign TLB_1_xor17 = TLB_1_xor35 ^ TLB_1_xor36;
  assign TLB_1_xor75 = mux_cond_14_pad ^ mux_cond_15_pad;
  assign TLB_1_xor76 = mux_cond_16_pad ^ mux_cond_17_pad;
  assign TLB_1_xor37 = TLB_1_xor75 ^ TLB_1_xor76;
  assign TLB_1_xor77 = mux_cond_18_pad ^ mux_cond_19_pad;
  assign TLB_1_xor78 = mux_cond_20_pad ^ mux_cond_21_pad;
  assign TLB_1_xor38 = TLB_1_xor77 ^ TLB_1_xor78;
  assign TLB_1_xor18 = TLB_1_xor37 ^ TLB_1_xor38;
  assign TLB_1_xor8 = TLB_1_xor17 ^ TLB_1_xor18;
  assign TLB_1_xor3 = TLB_1_xor7 ^ TLB_1_xor8;
  assign TLB_1_xor80 = mux_cond_23_pad ^ mux_cond_24_pad;
  assign TLB_1_xor39 = mux_cond_22_pad ^ TLB_1_xor80;
  assign TLB_1_xor81 = mux_cond_25_pad ^ mux_cond_26_pad;
  assign TLB_1_xor82 = mux_cond_27_pad ^ mux_cond_28_pad;
  assign TLB_1_xor40 = TLB_1_xor81 ^ TLB_1_xor82;
  assign TLB_1_xor19 = TLB_1_xor39 ^ TLB_1_xor40;
  assign TLB_1_xor84 = mux_cond_30_pad ^ mux_cond_31_pad;
  assign TLB_1_xor41 = mux_cond_29_pad ^ TLB_1_xor84;
  assign TLB_1_xor85 = mux_cond_32_pad ^ mux_cond_33_pad;
  assign TLB_1_xor86 = mux_cond_34_pad ^ mux_cond_35_pad;
  assign TLB_1_xor42 = TLB_1_xor85 ^ TLB_1_xor86;
  assign TLB_1_xor20 = TLB_1_xor41 ^ TLB_1_xor42;
  assign TLB_1_xor9 = TLB_1_xor19 ^ TLB_1_xor20;
  assign TLB_1_xor88 = mux_cond_37_pad ^ mux_cond_38_pad;
  assign TLB_1_xor43 = mux_cond_36_pad ^ TLB_1_xor88;
  assign TLB_1_xor89 = mux_cond_39_pad ^ mux_cond_40_pad;
  assign TLB_1_xor90 = mux_cond_41_pad ^ mux_cond_42_pad;
  assign TLB_1_xor44 = TLB_1_xor89 ^ TLB_1_xor90;
  assign TLB_1_xor21 = TLB_1_xor43 ^ TLB_1_xor44;
  assign TLB_1_xor91 = mux_cond_43_pad ^ mux_cond_44_pad;
  assign TLB_1_xor92 = mux_cond_45_pad ^ mux_cond_46_pad;
  assign TLB_1_xor45 = TLB_1_xor91 ^ TLB_1_xor92;
  assign TLB_1_xor93 = mux_cond_47_pad ^ mux_cond_48_pad;
  assign TLB_1_xor94 = mux_cond_49_pad ^ mux_cond_50_pad;
  assign TLB_1_xor46 = TLB_1_xor93 ^ TLB_1_xor94;
  assign TLB_1_xor22 = TLB_1_xor45 ^ TLB_1_xor46;
  assign TLB_1_xor10 = TLB_1_xor21 ^ TLB_1_xor22;
  assign TLB_1_xor4 = TLB_1_xor9 ^ TLB_1_xor10;
  assign TLB_1_xor1 = TLB_1_xor3 ^ TLB_1_xor4;
  assign TLB_1_xor96 = mux_cond_52_pad ^ mux_cond_53_pad;
  assign TLB_1_xor47 = mux_cond_51_pad ^ TLB_1_xor96;
  assign TLB_1_xor97 = mux_cond_54_pad ^ mux_cond_55_pad;
  assign TLB_1_xor98 = mux_cond_56_pad ^ mux_cond_57_pad;
  assign TLB_1_xor48 = TLB_1_xor97 ^ TLB_1_xor98;
  assign TLB_1_xor23 = TLB_1_xor47 ^ TLB_1_xor48;
  assign TLB_1_xor100 = mux_cond_59_pad ^ mux_cond_60_pad;
  assign TLB_1_xor49 = mux_cond_58_pad ^ TLB_1_xor100;
  assign TLB_1_xor101 = mux_cond_61_pad ^ mux_cond_62_pad;
  assign TLB_1_xor102 = mux_cond_63_pad ^ mux_cond_64_pad;
  assign TLB_1_xor50 = TLB_1_xor101 ^ TLB_1_xor102;
  assign TLB_1_xor24 = TLB_1_xor49 ^ TLB_1_xor50;
  assign TLB_1_xor11 = TLB_1_xor23 ^ TLB_1_xor24;
  assign TLB_1_xor104 = mux_cond_66_pad ^ mux_cond_67_pad;
  assign TLB_1_xor51 = mux_cond_65_pad ^ TLB_1_xor104;
  assign TLB_1_xor105 = mux_cond_68_pad ^ sectored_entries_0_0_valid_3_pad;
  assign TLB_1_xor106 = sectored_entries_0_0_valid_2_pad ^ sectored_entries_0_2_valid_0_pad;
  assign TLB_1_xor52 = TLB_1_xor105 ^ TLB_1_xor106;
  assign TLB_1_xor25 = TLB_1_xor51 ^ TLB_1_xor52;
  assign TLB_1_xor107 = sectored_entries_0_3_valid_0_pad ^ superpage_entries_2_level_pad;
  assign TLB_1_xor108 = sectored_entries_0_7_valid_1_pad ^ sectored_entries_0_4_valid_0_pad;
  assign TLB_1_xor53 = TLB_1_xor107 ^ TLB_1_xor108;
  assign TLB_1_xor109 = sectored_entries_0_1_valid_3_pad ^ sectored_entries_0_1_valid_1_pad;
  assign TLB_1_xor110 = sectored_entries_0_2_valid_3_pad ^ sectored_entries_0_2_valid_1_pad;
  assign TLB_1_xor54 = TLB_1_xor109 ^ TLB_1_xor110;
  assign TLB_1_xor26 = TLB_1_xor53 ^ TLB_1_xor54;
  assign TLB_1_xor12 = TLB_1_xor25 ^ TLB_1_xor26;
  assign TLB_1_xor5 = TLB_1_xor11 ^ TLB_1_xor12;
  assign TLB_1_xor112 = sectored_entries_0_7_valid_0_pad ^ superpage_entries_3_valid_0_pad;
  assign TLB_1_xor55 = superpage_entries_1_valid_0_pad ^ TLB_1_xor112;
  assign TLB_1_xor113 = sectored_entries_0_5_valid_3_pad ^ sectored_entries_0_5_valid_1_pad;
  assign TLB_1_xor114 = sectored_entries_0_4_valid_3_pad ^ sectored_entries_0_5_valid_2_pad;
  assign TLB_1_xor56 = TLB_1_xor113 ^ TLB_1_xor114;
  assign TLB_1_xor27 = TLB_1_xor55 ^ TLB_1_xor56;
  assign TLB_1_xor116 = sectored_entries_0_3_valid_1_pad ^ sectored_entries_0_1_valid_0_pad;
  assign TLB_1_xor57 = sectored_entries_0_1_valid_2_pad ^ TLB_1_xor116;
  assign TLB_1_xor117 = sectored_entries_0_4_valid_2_pad ^ sectored_entries_0_4_valid_1_pad;
  assign TLB_1_xor118 = superpage_entries_3_level_pad ^ sectored_entries_0_0_valid_1_pad;
  assign TLB_1_xor58 = TLB_1_xor117 ^ TLB_1_xor118;
  assign TLB_1_xor28 = TLB_1_xor57 ^ TLB_1_xor58;
  assign TLB_1_xor13 = TLB_1_xor27 ^ TLB_1_xor28;
  assign TLB_1_xor120 = sectored_entries_0_6_valid_1_pad ^ sectored_entries_0_7_valid_3_pad;
  assign TLB_1_xor59 = sectored_entries_0_3_valid_2_pad ^ TLB_1_xor120;
  assign TLB_1_xor121 = sectored_entries_0_3_valid_3_pad ^ sectored_entries_0_0_valid_0_pad;
  assign TLB_1_xor122 = superpage_entries_0_valid_0_pad ^ sectored_entries_0_2_valid_2_pad;
  assign TLB_1_xor60 = TLB_1_xor121 ^ TLB_1_xor122;
  assign TLB_1_xor29 = TLB_1_xor59 ^ TLB_1_xor60;
  assign TLB_1_xor123 = sectored_entries_0_6_valid_2_pad ^ superpage_entries_2_valid_0_pad;
  assign TLB_1_xor124 = sectored_entries_0_6_valid_3_pad ^ sectored_entries_0_6_valid_0_pad;
  assign TLB_1_xor61 = TLB_1_xor123 ^ TLB_1_xor124;
  assign TLB_1_xor125 = sectored_entries_0_7_valid_2_pad ^ superpage_entries_0_level_pad;
  assign TLB_1_xor126 = superpage_entries_1_level_pad ^ sectored_entries_0_5_valid_0_pad;
  assign TLB_1_xor62 = TLB_1_xor125 ^ TLB_1_xor126;
  assign TLB_1_xor30 = TLB_1_xor61 ^ TLB_1_xor62;
  assign TLB_1_xor14 = TLB_1_xor29 ^ TLB_1_xor30;
  assign TLB_1_xor6 = TLB_1_xor13 ^ TLB_1_xor14;
  assign TLB_1_xor2 = TLB_1_xor5 ^ TLB_1_xor6;
  assign TLB_1_xor0 = TLB_1_xor1 ^ TLB_1_xor2;
  assign mpu_ppn_barrier_sum = TLB_1_covSum + mpu_ppn_barrier_io_covSum;
  assign entries_barrier_10_sum = mpu_ppn_barrier_sum + entries_barrier_10_io_covSum;
  assign entries_barrier_9_sum = entries_barrier_10_sum + entries_barrier_9_io_covSum;
  assign entries_barrier_7_sum = entries_barrier_9_sum + entries_barrier_7_io_covSum;
  assign entries_barrier_sum = entries_barrier_7_sum + entries_barrier_io_covSum;
  assign pmp_sum = entries_barrier_sum + pmp_io_covSum;
  assign entries_barrier_6_sum = pmp_sum + entries_barrier_6_io_covSum;
  assign entries_barrier_12_sum = entries_barrier_6_sum + entries_barrier_12_io_covSum;
  assign entries_barrier_1_sum = entries_barrier_12_sum + entries_barrier_1_io_covSum;
  assign entries_barrier_11_sum = entries_barrier_1_sum + entries_barrier_11_io_covSum;
  assign entries_barrier_8_sum = entries_barrier_11_sum + entries_barrier_8_io_covSum;
  assign entries_barrier_2_sum = entries_barrier_8_sum + entries_barrier_2_io_covSum;
  assign entries_barrier_4_sum = entries_barrier_2_sum + entries_barrier_4_io_covSum;
  assign entries_barrier_5_sum = entries_barrier_4_sum + entries_barrier_5_io_covSum;
  assign entries_barrier_3_sum = entries_barrier_5_sum + entries_barrier_3_io_covSum;
  assign io_covSum = entries_barrier_3_sum;
  assign stopEn0 = io_sfence_valid & ~_T_51;
  assign entries_barrier_12_metaAssert_wire = entries_barrier_12_metaAssert;
  assign entries_barrier_metaAssert_wire = entries_barrier_metaAssert;
  assign entries_barrier_10_metaAssert_wire = entries_barrier_10_metaAssert;
  assign entries_barrier_5_metaAssert_wire = entries_barrier_5_metaAssert;
  assign entries_barrier_11_metaAssert_wire = entries_barrier_11_metaAssert;
  assign entries_barrier_9_metaAssert_wire = entries_barrier_9_metaAssert;
  assign entries_barrier_8_metaAssert_wire = entries_barrier_8_metaAssert;
  assign entries_barrier_1_metaAssert_wire = entries_barrier_1_metaAssert;
  assign mpu_ppn_barrier_metaAssert_wire = mpu_ppn_barrier_metaAssert;
  assign entries_barrier_4_metaAssert_wire = entries_barrier_4_metaAssert;
  assign entries_barrier_6_metaAssert_wire = entries_barrier_6_metaAssert;
  assign entries_barrier_3_metaAssert_wire = entries_barrier_3_metaAssert;
  assign pmp_metaAssert_wire = pmp_metaAssert;
  assign entries_barrier_7_metaAssert_wire = entries_barrier_7_metaAssert;
  assign entries_barrier_2_metaAssert_wire = entries_barrier_2_metaAssert;
  assign TLB_1_or7 = stopEn0 | entries_barrier_6_metaAssert_wire;
  assign TLB_1_or8 = entries_barrier_10_metaAssert_wire | entries_barrier_7_metaAssert_wire;
  assign TLB_1_or3 = TLB_1_or7 | TLB_1_or8;
  assign TLB_1_or9 = entries_barrier_4_metaAssert_wire | entries_barrier_11_metaAssert_wire;
  assign TLB_1_or10 = entries_barrier_8_metaAssert_wire | entries_barrier_9_metaAssert_wire;
  assign TLB_1_or4 = TLB_1_or9 | TLB_1_or10;
  assign TLB_1_or1 = TLB_1_or3 | TLB_1_or4;
  assign TLB_1_or11 = entries_barrier_metaAssert_wire | entries_barrier_3_metaAssert_wire;
  assign TLB_1_or12 = pmp_metaAssert_wire | mpu_ppn_barrier_metaAssert_wire;
  assign TLB_1_or5 = TLB_1_or11 | TLB_1_or12;
  assign TLB_1_or13 = entries_barrier_12_metaAssert_wire | entries_barrier_5_metaAssert_wire;
  assign TLB_1_or14 = entries_barrier_2_metaAssert_wire | entries_barrier_1_metaAssert_wire;
  assign TLB_1_or6 = TLB_1_or13 | TLB_1_or14;
  assign TLB_1_or2 = TLB_1_or5 | TLB_1_or6;
  assign TLB_1_or0 = TLB_1_or1 | TLB_1_or2;
  assign metaAssert = TLB_1_metaAssert;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sectored_entries_0_0_tag = _RAND_0[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {2{`RANDOM}};
  sectored_entries_0_0_data_0 = _RAND_1[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {2{`RANDOM}};
  sectored_entries_0_0_data_1 = _RAND_2[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {2{`RANDOM}};
  sectored_entries_0_0_data_2 = _RAND_3[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {2{`RANDOM}};
  sectored_entries_0_0_data_3 = _RAND_4[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  sectored_entries_0_0_valid_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  sectored_entries_0_0_valid_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  sectored_entries_0_0_valid_2 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  sectored_entries_0_0_valid_3 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  sectored_entries_0_1_tag = _RAND_9[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {2{`RANDOM}};
  sectored_entries_0_1_data_0 = _RAND_10[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {2{`RANDOM}};
  sectored_entries_0_1_data_1 = _RAND_11[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {2{`RANDOM}};
  sectored_entries_0_1_data_2 = _RAND_12[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {2{`RANDOM}};
  sectored_entries_0_1_data_3 = _RAND_13[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  sectored_entries_0_1_valid_0 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  sectored_entries_0_1_valid_1 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  sectored_entries_0_1_valid_2 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  sectored_entries_0_1_valid_3 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  sectored_entries_0_2_tag = _RAND_18[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {2{`RANDOM}};
  sectored_entries_0_2_data_0 = _RAND_19[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {2{`RANDOM}};
  sectored_entries_0_2_data_1 = _RAND_20[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {2{`RANDOM}};
  sectored_entries_0_2_data_2 = _RAND_21[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {2{`RANDOM}};
  sectored_entries_0_2_data_3 = _RAND_22[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  sectored_entries_0_2_valid_0 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  sectored_entries_0_2_valid_1 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  sectored_entries_0_2_valid_2 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  sectored_entries_0_2_valid_3 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  sectored_entries_0_3_tag = _RAND_27[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {2{`RANDOM}};
  sectored_entries_0_3_data_0 = _RAND_28[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {2{`RANDOM}};
  sectored_entries_0_3_data_1 = _RAND_29[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {2{`RANDOM}};
  sectored_entries_0_3_data_2 = _RAND_30[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {2{`RANDOM}};
  sectored_entries_0_3_data_3 = _RAND_31[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  sectored_entries_0_3_valid_0 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  sectored_entries_0_3_valid_1 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  sectored_entries_0_3_valid_2 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  sectored_entries_0_3_valid_3 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  sectored_entries_0_4_tag = _RAND_36[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {2{`RANDOM}};
  sectored_entries_0_4_data_0 = _RAND_37[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {2{`RANDOM}};
  sectored_entries_0_4_data_1 = _RAND_38[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {2{`RANDOM}};
  sectored_entries_0_4_data_2 = _RAND_39[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {2{`RANDOM}};
  sectored_entries_0_4_data_3 = _RAND_40[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  sectored_entries_0_4_valid_0 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  sectored_entries_0_4_valid_1 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  sectored_entries_0_4_valid_2 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  sectored_entries_0_4_valid_3 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  sectored_entries_0_5_tag = _RAND_45[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {2{`RANDOM}};
  sectored_entries_0_5_data_0 = _RAND_46[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {2{`RANDOM}};
  sectored_entries_0_5_data_1 = _RAND_47[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {2{`RANDOM}};
  sectored_entries_0_5_data_2 = _RAND_48[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {2{`RANDOM}};
  sectored_entries_0_5_data_3 = _RAND_49[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  sectored_entries_0_5_valid_0 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  sectored_entries_0_5_valid_1 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  sectored_entries_0_5_valid_2 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  sectored_entries_0_5_valid_3 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  sectored_entries_0_6_tag = _RAND_54[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {2{`RANDOM}};
  sectored_entries_0_6_data_0 = _RAND_55[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {2{`RANDOM}};
  sectored_entries_0_6_data_1 = _RAND_56[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {2{`RANDOM}};
  sectored_entries_0_6_data_2 = _RAND_57[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {2{`RANDOM}};
  sectored_entries_0_6_data_3 = _RAND_58[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  sectored_entries_0_6_valid_0 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  sectored_entries_0_6_valid_1 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  sectored_entries_0_6_valid_2 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  sectored_entries_0_6_valid_3 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  sectored_entries_0_7_tag = _RAND_63[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {2{`RANDOM}};
  sectored_entries_0_7_data_0 = _RAND_64[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {2{`RANDOM}};
  sectored_entries_0_7_data_1 = _RAND_65[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {2{`RANDOM}};
  sectored_entries_0_7_data_2 = _RAND_66[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {2{`RANDOM}};
  sectored_entries_0_7_data_3 = _RAND_67[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  sectored_entries_0_7_valid_0 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  sectored_entries_0_7_valid_1 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  sectored_entries_0_7_valid_2 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  sectored_entries_0_7_valid_3 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  superpage_entries_0_level = _RAND_72[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  superpage_entries_0_tag = _RAND_73[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {2{`RANDOM}};
  superpage_entries_0_data_0 = _RAND_74[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  superpage_entries_0_valid_0 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  superpage_entries_1_level = _RAND_76[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  superpage_entries_1_tag = _RAND_77[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {2{`RANDOM}};
  superpage_entries_1_data_0 = _RAND_78[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  superpage_entries_1_valid_0 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  superpage_entries_2_level = _RAND_80[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  superpage_entries_2_tag = _RAND_81[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {2{`RANDOM}};
  superpage_entries_2_data_0 = _RAND_82[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  superpage_entries_2_valid_0 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  superpage_entries_3_level = _RAND_84[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  superpage_entries_3_tag = _RAND_85[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {2{`RANDOM}};
  superpage_entries_3_data_0 = _RAND_86[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  superpage_entries_3_valid_0 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  special_entry_level = _RAND_88[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  special_entry_tag = _RAND_89[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {2{`RANDOM}};
  special_entry_data_0 = _RAND_90[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  special_entry_valid_0 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  state = _RAND_92[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  r_refill_tag = _RAND_93[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  r_superpage_repl_addr = _RAND_94[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  r_sectored_repl_addr = _RAND_95[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  r_sectored_hit_addr = _RAND_96[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  r_sectored_hit = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  state_vec_0 = _RAND_98[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  state_reg_1 = _RAND_99[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  TLB_1_state = _RAND_100[19:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1048576; initvar = initvar+1)
    TLB_1_cov[initvar] = _RAND_101[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  TLB_1_covSum = _RAND_102[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  TLB_1_metaAssert = _RAND_103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      sectored_entries_0_0_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_7) begin
            sectored_entries_0_0_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_0_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_7) begin
            if (2'h0 == idx) begin
              sectored_entries_0_0_data_0 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_0_data_1 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_7) begin
            if (2'h1 == idx) begin
              sectored_entries_0_0_data_1 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_0_data_2 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_7) begin
            if (2'h2 == idx) begin
              sectored_entries_0_0_data_2 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_0_data_3 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_7) begin
            if (2'h3 == idx) begin
              sectored_entries_0_0_data_3 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_0_valid_0 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_0_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_59) begin
          if (sectored_entries_0_0_data_0[0]) begin
            sectored_entries_0_0_valid_0 <= 1'h0;
          end else if (_sector_hits_T_5) begin
            if (2'h0 == hitsVec_idx) begin
              sectored_entries_0_0_valid_0 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_7) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_0_valid_0 <= 1'h0;
                    end else begin
                      sectored_entries_0_0_valid_0 <= _GEN_53;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_7) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_0_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_0_0_valid_0 <= _GEN_53;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_5) begin
          if (2'h0 == hitsVec_idx) begin
            sectored_entries_0_0_valid_0 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_7) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_0_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_0_0_valid_0 <= _GEN_53;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_7) begin
                if (invalidate_refill) begin
                  sectored_entries_0_0_valid_0 <= 1'h0;
                end else begin
                  sectored_entries_0_0_valid_0 <= _GEN_53;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_0_valid_0 <= _GEN_621;
      end
    end else begin
      sectored_entries_0_0_valid_0 <= _GEN_473;
    end
    if (metaReset) begin
      sectored_entries_0_0_valid_1 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_0_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_59) begin
          if (sectored_entries_0_0_data_1[0]) begin
            sectored_entries_0_0_valid_1 <= 1'h0;
          end else if (_sector_hits_T_5) begin
            if (2'h1 == hitsVec_idx) begin
              sectored_entries_0_0_valid_1 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_7) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_0_valid_1 <= 1'h0;
                    end else begin
                      sectored_entries_0_0_valid_1 <= _GEN_54;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_7) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_0_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_0_0_valid_1 <= _GEN_54;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_5) begin
          if (2'h1 == hitsVec_idx) begin
            sectored_entries_0_0_valid_1 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_7) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_0_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_0_0_valid_1 <= _GEN_54;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_7) begin
                if (invalidate_refill) begin
                  sectored_entries_0_0_valid_1 <= 1'h0;
                end else begin
                  sectored_entries_0_0_valid_1 <= _GEN_54;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_0_valid_1 <= _GEN_622;
      end
    end else begin
      sectored_entries_0_0_valid_1 <= _GEN_474;
    end
    if (metaReset) begin
      sectored_entries_0_0_valid_2 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_0_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_59) begin
          if (sectored_entries_0_0_data_2[0]) begin
            sectored_entries_0_0_valid_2 <= 1'h0;
          end else if (_sector_hits_T_5) begin
            if (2'h2 == hitsVec_idx) begin
              sectored_entries_0_0_valid_2 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_7) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_0_valid_2 <= 1'h0;
                    end else begin
                      sectored_entries_0_0_valid_2 <= _GEN_55;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_7) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_0_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_0_0_valid_2 <= _GEN_55;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_5) begin
          if (2'h2 == hitsVec_idx) begin
            sectored_entries_0_0_valid_2 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_7) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_0_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_0_0_valid_2 <= _GEN_55;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_7) begin
                if (invalidate_refill) begin
                  sectored_entries_0_0_valid_2 <= 1'h0;
                end else begin
                  sectored_entries_0_0_valid_2 <= _GEN_55;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_0_valid_2 <= _GEN_623;
      end
    end else begin
      sectored_entries_0_0_valid_2 <= _GEN_475;
    end
    if (metaReset) begin
      sectored_entries_0_0_valid_3 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_0_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_59) begin
          if (sectored_entries_0_0_data_3[0]) begin
            sectored_entries_0_0_valid_3 <= 1'h0;
          end else if (_sector_hits_T_5) begin
            if (2'h3 == hitsVec_idx) begin
              sectored_entries_0_0_valid_3 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_7) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_0_valid_3 <= 1'h0;
                    end else begin
                      sectored_entries_0_0_valid_3 <= _GEN_56;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_7) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_0_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_0_0_valid_3 <= _GEN_56;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_5) begin
          if (2'h3 == hitsVec_idx) begin
            sectored_entries_0_0_valid_3 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_7) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_0_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_0_0_valid_3 <= _GEN_56;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_7) begin
                if (invalidate_refill) begin
                  sectored_entries_0_0_valid_3 <= 1'h0;
                end else begin
                  sectored_entries_0_0_valid_3 <= _GEN_56;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_0_valid_3 <= _GEN_624;
      end
    end else begin
      sectored_entries_0_0_valid_3 <= _GEN_476;
    end
    if (metaReset) begin
      sectored_entries_0_1_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_9) begin
            sectored_entries_0_1_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_1_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_9) begin
            if (2'h0 == idx) begin
              sectored_entries_0_1_data_0 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_1_data_1 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_9) begin
            if (2'h1 == idx) begin
              sectored_entries_0_1_data_1 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_1_data_2 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_9) begin
            if (2'h2 == idx) begin
              sectored_entries_0_1_data_2 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_1_data_3 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_9) begin
            if (2'h3 == idx) begin
              sectored_entries_0_1_data_3 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_1_valid_0 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_1_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_198) begin
          if (sectored_entries_0_1_data_0[0]) begin
            sectored_entries_0_1_valid_0 <= 1'h0;
          end else if (_sector_hits_T_11) begin
            if (2'h0 == hitsVec_idx) begin
              sectored_entries_0_1_valid_0 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_9) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_1_valid_0 <= 1'h0;
                    end else begin
                      sectored_entries_0_1_valid_0 <= _GEN_79;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_9) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_1_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_0_1_valid_0 <= _GEN_79;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_11) begin
          if (2'h0 == hitsVec_idx) begin
            sectored_entries_0_1_valid_0 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_9) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_1_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_0_1_valid_0 <= _GEN_79;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_9) begin
                if (invalidate_refill) begin
                  sectored_entries_0_1_valid_0 <= 1'h0;
                end else begin
                  sectored_entries_0_1_valid_0 <= _GEN_79;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_1_valid_0 <= _GEN_649;
      end
    end else begin
      sectored_entries_0_1_valid_0 <= _GEN_483;
    end
    if (metaReset) begin
      sectored_entries_0_1_valid_1 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_1_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_198) begin
          if (sectored_entries_0_1_data_1[0]) begin
            sectored_entries_0_1_valid_1 <= 1'h0;
          end else if (_sector_hits_T_11) begin
            if (2'h1 == hitsVec_idx) begin
              sectored_entries_0_1_valid_1 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_9) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_1_valid_1 <= 1'h0;
                    end else begin
                      sectored_entries_0_1_valid_1 <= _GEN_80;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_9) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_1_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_0_1_valid_1 <= _GEN_80;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_11) begin
          if (2'h1 == hitsVec_idx) begin
            sectored_entries_0_1_valid_1 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_9) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_1_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_0_1_valid_1 <= _GEN_80;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_9) begin
                if (invalidate_refill) begin
                  sectored_entries_0_1_valid_1 <= 1'h0;
                end else begin
                  sectored_entries_0_1_valid_1 <= _GEN_80;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_1_valid_1 <= _GEN_650;
      end
    end else begin
      sectored_entries_0_1_valid_1 <= _GEN_484;
    end
    if (metaReset) begin
      sectored_entries_0_1_valid_2 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_1_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_198) begin
          if (sectored_entries_0_1_data_2[0]) begin
            sectored_entries_0_1_valid_2 <= 1'h0;
          end else if (_sector_hits_T_11) begin
            if (2'h2 == hitsVec_idx) begin
              sectored_entries_0_1_valid_2 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_9) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_1_valid_2 <= 1'h0;
                    end else begin
                      sectored_entries_0_1_valid_2 <= _GEN_81;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_9) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_1_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_0_1_valid_2 <= _GEN_81;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_11) begin
          if (2'h2 == hitsVec_idx) begin
            sectored_entries_0_1_valid_2 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_9) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_1_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_0_1_valid_2 <= _GEN_81;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_9) begin
                if (invalidate_refill) begin
                  sectored_entries_0_1_valid_2 <= 1'h0;
                end else begin
                  sectored_entries_0_1_valid_2 <= _GEN_81;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_1_valid_2 <= _GEN_651;
      end
    end else begin
      sectored_entries_0_1_valid_2 <= _GEN_485;
    end
    if (metaReset) begin
      sectored_entries_0_1_valid_3 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_1_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_198) begin
          if (sectored_entries_0_1_data_3[0]) begin
            sectored_entries_0_1_valid_3 <= 1'h0;
          end else if (_sector_hits_T_11) begin
            if (2'h3 == hitsVec_idx) begin
              sectored_entries_0_1_valid_3 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_9) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_1_valid_3 <= 1'h0;
                    end else begin
                      sectored_entries_0_1_valid_3 <= _GEN_82;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_9) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_1_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_0_1_valid_3 <= _GEN_82;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_11) begin
          if (2'h3 == hitsVec_idx) begin
            sectored_entries_0_1_valid_3 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_9) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_1_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_0_1_valid_3 <= _GEN_82;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_9) begin
                if (invalidate_refill) begin
                  sectored_entries_0_1_valid_3 <= 1'h0;
                end else begin
                  sectored_entries_0_1_valid_3 <= _GEN_82;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_1_valid_3 <= _GEN_652;
      end
    end else begin
      sectored_entries_0_1_valid_3 <= _GEN_486;
    end
    if (metaReset) begin
      sectored_entries_0_2_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_11) begin
            sectored_entries_0_2_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_2_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_11) begin
            if (2'h0 == idx) begin
              sectored_entries_0_2_data_0 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_2_data_1 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_11) begin
            if (2'h1 == idx) begin
              sectored_entries_0_2_data_1 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_2_data_2 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_11) begin
            if (2'h2 == idx) begin
              sectored_entries_0_2_data_2 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_2_data_3 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_11) begin
            if (2'h3 == idx) begin
              sectored_entries_0_2_data_3 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_2_valid_0 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_2_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_337) begin
          if (sectored_entries_0_2_data_0[0]) begin
            sectored_entries_0_2_valid_0 <= 1'h0;
          end else if (_sector_hits_T_17) begin
            if (2'h0 == hitsVec_idx) begin
              sectored_entries_0_2_valid_0 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_11) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_2_valid_0 <= 1'h0;
                    end else begin
                      sectored_entries_0_2_valid_0 <= _GEN_105;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_11) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_2_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_0_2_valid_0 <= _GEN_105;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_17) begin
          if (2'h0 == hitsVec_idx) begin
            sectored_entries_0_2_valid_0 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_11) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_2_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_0_2_valid_0 <= _GEN_105;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_11) begin
                if (invalidate_refill) begin
                  sectored_entries_0_2_valid_0 <= 1'h0;
                end else begin
                  sectored_entries_0_2_valid_0 <= _GEN_105;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_2_valid_0 <= _GEN_677;
      end
    end else begin
      sectored_entries_0_2_valid_0 <= _GEN_493;
    end
    if (metaReset) begin
      sectored_entries_0_2_valid_1 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_2_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_337) begin
          if (sectored_entries_0_2_data_1[0]) begin
            sectored_entries_0_2_valid_1 <= 1'h0;
          end else if (_sector_hits_T_17) begin
            if (2'h1 == hitsVec_idx) begin
              sectored_entries_0_2_valid_1 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_11) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_2_valid_1 <= 1'h0;
                    end else begin
                      sectored_entries_0_2_valid_1 <= _GEN_106;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_11) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_2_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_0_2_valid_1 <= _GEN_106;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_17) begin
          if (2'h1 == hitsVec_idx) begin
            sectored_entries_0_2_valid_1 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_11) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_2_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_0_2_valid_1 <= _GEN_106;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_11) begin
                if (invalidate_refill) begin
                  sectored_entries_0_2_valid_1 <= 1'h0;
                end else begin
                  sectored_entries_0_2_valid_1 <= _GEN_106;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_2_valid_1 <= _GEN_678;
      end
    end else begin
      sectored_entries_0_2_valid_1 <= _GEN_494;
    end
    if (metaReset) begin
      sectored_entries_0_2_valid_2 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_2_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_337) begin
          if (sectored_entries_0_2_data_2[0]) begin
            sectored_entries_0_2_valid_2 <= 1'h0;
          end else if (_sector_hits_T_17) begin
            if (2'h2 == hitsVec_idx) begin
              sectored_entries_0_2_valid_2 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_11) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_2_valid_2 <= 1'h0;
                    end else begin
                      sectored_entries_0_2_valid_2 <= _GEN_107;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_11) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_2_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_0_2_valid_2 <= _GEN_107;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_17) begin
          if (2'h2 == hitsVec_idx) begin
            sectored_entries_0_2_valid_2 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_11) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_2_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_0_2_valid_2 <= _GEN_107;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_11) begin
                if (invalidate_refill) begin
                  sectored_entries_0_2_valid_2 <= 1'h0;
                end else begin
                  sectored_entries_0_2_valid_2 <= _GEN_107;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_2_valid_2 <= _GEN_679;
      end
    end else begin
      sectored_entries_0_2_valid_2 <= _GEN_495;
    end
    if (metaReset) begin
      sectored_entries_0_2_valid_3 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_2_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_337) begin
          if (sectored_entries_0_2_data_3[0]) begin
            sectored_entries_0_2_valid_3 <= 1'h0;
          end else if (_sector_hits_T_17) begin
            if (2'h3 == hitsVec_idx) begin
              sectored_entries_0_2_valid_3 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_11) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_2_valid_3 <= 1'h0;
                    end else begin
                      sectored_entries_0_2_valid_3 <= _GEN_108;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_11) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_2_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_0_2_valid_3 <= _GEN_108;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_17) begin
          if (2'h3 == hitsVec_idx) begin
            sectored_entries_0_2_valid_3 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_11) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_2_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_0_2_valid_3 <= _GEN_108;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_11) begin
                if (invalidate_refill) begin
                  sectored_entries_0_2_valid_3 <= 1'h0;
                end else begin
                  sectored_entries_0_2_valid_3 <= _GEN_108;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_2_valid_3 <= _GEN_680;
      end
    end else begin
      sectored_entries_0_2_valid_3 <= _GEN_496;
    end
    if (metaReset) begin
      sectored_entries_0_3_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_13) begin
            sectored_entries_0_3_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_3_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_13) begin
            if (2'h0 == idx) begin
              sectored_entries_0_3_data_0 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_3_data_1 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_13) begin
            if (2'h1 == idx) begin
              sectored_entries_0_3_data_1 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_3_data_2 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_13) begin
            if (2'h2 == idx) begin
              sectored_entries_0_3_data_2 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_3_data_3 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_13) begin
            if (2'h3 == idx) begin
              sectored_entries_0_3_data_3 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_3_valid_0 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_3_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_476) begin
          if (sectored_entries_0_3_data_0[0]) begin
            sectored_entries_0_3_valid_0 <= 1'h0;
          end else if (_sector_hits_T_23) begin
            if (2'h0 == hitsVec_idx) begin
              sectored_entries_0_3_valid_0 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_13) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_3_valid_0 <= 1'h0;
                    end else begin
                      sectored_entries_0_3_valid_0 <= _GEN_131;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_13) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_3_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_0_3_valid_0 <= _GEN_131;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_23) begin
          if (2'h0 == hitsVec_idx) begin
            sectored_entries_0_3_valid_0 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_13) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_3_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_0_3_valid_0 <= _GEN_131;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_13) begin
                if (invalidate_refill) begin
                  sectored_entries_0_3_valid_0 <= 1'h0;
                end else begin
                  sectored_entries_0_3_valid_0 <= _GEN_131;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_3_valid_0 <= _GEN_705;
      end
    end else begin
      sectored_entries_0_3_valid_0 <= _GEN_503;
    end
    if (metaReset) begin
      sectored_entries_0_3_valid_1 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_3_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_476) begin
          if (sectored_entries_0_3_data_1[0]) begin
            sectored_entries_0_3_valid_1 <= 1'h0;
          end else if (_sector_hits_T_23) begin
            if (2'h1 == hitsVec_idx) begin
              sectored_entries_0_3_valid_1 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_13) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_3_valid_1 <= 1'h0;
                    end else begin
                      sectored_entries_0_3_valid_1 <= _GEN_132;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_13) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_3_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_0_3_valid_1 <= _GEN_132;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_23) begin
          if (2'h1 == hitsVec_idx) begin
            sectored_entries_0_3_valid_1 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_13) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_3_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_0_3_valid_1 <= _GEN_132;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_13) begin
                if (invalidate_refill) begin
                  sectored_entries_0_3_valid_1 <= 1'h0;
                end else begin
                  sectored_entries_0_3_valid_1 <= _GEN_132;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_3_valid_1 <= _GEN_706;
      end
    end else begin
      sectored_entries_0_3_valid_1 <= _GEN_504;
    end
    if (metaReset) begin
      sectored_entries_0_3_valid_2 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_3_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_476) begin
          if (sectored_entries_0_3_data_2[0]) begin
            sectored_entries_0_3_valid_2 <= 1'h0;
          end else if (_sector_hits_T_23) begin
            if (2'h2 == hitsVec_idx) begin
              sectored_entries_0_3_valid_2 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_13) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_3_valid_2 <= 1'h0;
                    end else begin
                      sectored_entries_0_3_valid_2 <= _GEN_133;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_13) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_3_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_0_3_valid_2 <= _GEN_133;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_23) begin
          if (2'h2 == hitsVec_idx) begin
            sectored_entries_0_3_valid_2 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_13) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_3_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_0_3_valid_2 <= _GEN_133;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_13) begin
                if (invalidate_refill) begin
                  sectored_entries_0_3_valid_2 <= 1'h0;
                end else begin
                  sectored_entries_0_3_valid_2 <= _GEN_133;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_3_valid_2 <= _GEN_707;
      end
    end else begin
      sectored_entries_0_3_valid_2 <= _GEN_505;
    end
    if (metaReset) begin
      sectored_entries_0_3_valid_3 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_3_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_476) begin
          if (sectored_entries_0_3_data_3[0]) begin
            sectored_entries_0_3_valid_3 <= 1'h0;
          end else if (_sector_hits_T_23) begin
            if (2'h3 == hitsVec_idx) begin
              sectored_entries_0_3_valid_3 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_13) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_3_valid_3 <= 1'h0;
                    end else begin
                      sectored_entries_0_3_valid_3 <= _GEN_134;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_13) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_3_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_0_3_valid_3 <= _GEN_134;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_23) begin
          if (2'h3 == hitsVec_idx) begin
            sectored_entries_0_3_valid_3 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_13) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_3_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_0_3_valid_3 <= _GEN_134;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_13) begin
                if (invalidate_refill) begin
                  sectored_entries_0_3_valid_3 <= 1'h0;
                end else begin
                  sectored_entries_0_3_valid_3 <= _GEN_134;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_3_valid_3 <= _GEN_708;
      end
    end else begin
      sectored_entries_0_3_valid_3 <= _GEN_506;
    end
    if (metaReset) begin
      sectored_entries_0_4_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_15) begin
            sectored_entries_0_4_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_4_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_15) begin
            if (2'h0 == idx) begin
              sectored_entries_0_4_data_0 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_4_data_1 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_15) begin
            if (2'h1 == idx) begin
              sectored_entries_0_4_data_1 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_4_data_2 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_15) begin
            if (2'h2 == idx) begin
              sectored_entries_0_4_data_2 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_4_data_3 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_15) begin
            if (2'h3 == idx) begin
              sectored_entries_0_4_data_3 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_4_valid_0 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_4_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_615) begin
          if (sectored_entries_0_4_data_0[0]) begin
            sectored_entries_0_4_valid_0 <= 1'h0;
          end else if (_sector_hits_T_29) begin
            if (2'h0 == hitsVec_idx) begin
              sectored_entries_0_4_valid_0 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_15) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_4_valid_0 <= 1'h0;
                    end else begin
                      sectored_entries_0_4_valid_0 <= _GEN_157;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_15) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_4_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_0_4_valid_0 <= _GEN_157;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_29) begin
          if (2'h0 == hitsVec_idx) begin
            sectored_entries_0_4_valid_0 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_15) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_4_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_0_4_valid_0 <= _GEN_157;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_15) begin
                if (invalidate_refill) begin
                  sectored_entries_0_4_valid_0 <= 1'h0;
                end else begin
                  sectored_entries_0_4_valid_0 <= _GEN_157;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_4_valid_0 <= _GEN_733;
      end
    end else begin
      sectored_entries_0_4_valid_0 <= _GEN_513;
    end
    if (metaReset) begin
      sectored_entries_0_4_valid_1 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_4_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_615) begin
          if (sectored_entries_0_4_data_1[0]) begin
            sectored_entries_0_4_valid_1 <= 1'h0;
          end else if (_sector_hits_T_29) begin
            if (2'h1 == hitsVec_idx) begin
              sectored_entries_0_4_valid_1 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_15) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_4_valid_1 <= 1'h0;
                    end else begin
                      sectored_entries_0_4_valid_1 <= _GEN_158;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_15) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_4_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_0_4_valid_1 <= _GEN_158;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_29) begin
          if (2'h1 == hitsVec_idx) begin
            sectored_entries_0_4_valid_1 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_15) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_4_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_0_4_valid_1 <= _GEN_158;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_15) begin
                if (invalidate_refill) begin
                  sectored_entries_0_4_valid_1 <= 1'h0;
                end else begin
                  sectored_entries_0_4_valid_1 <= _GEN_158;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_4_valid_1 <= _GEN_734;
      end
    end else begin
      sectored_entries_0_4_valid_1 <= _GEN_514;
    end
    if (metaReset) begin
      sectored_entries_0_4_valid_2 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_4_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_615) begin
          if (sectored_entries_0_4_data_2[0]) begin
            sectored_entries_0_4_valid_2 <= 1'h0;
          end else if (_sector_hits_T_29) begin
            if (2'h2 == hitsVec_idx) begin
              sectored_entries_0_4_valid_2 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_15) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_4_valid_2 <= 1'h0;
                    end else begin
                      sectored_entries_0_4_valid_2 <= _GEN_159;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_15) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_4_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_0_4_valid_2 <= _GEN_159;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_29) begin
          if (2'h2 == hitsVec_idx) begin
            sectored_entries_0_4_valid_2 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_15) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_4_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_0_4_valid_2 <= _GEN_159;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_15) begin
                if (invalidate_refill) begin
                  sectored_entries_0_4_valid_2 <= 1'h0;
                end else begin
                  sectored_entries_0_4_valid_2 <= _GEN_159;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_4_valid_2 <= _GEN_735;
      end
    end else begin
      sectored_entries_0_4_valid_2 <= _GEN_515;
    end
    if (metaReset) begin
      sectored_entries_0_4_valid_3 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_4_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_615) begin
          if (sectored_entries_0_4_data_3[0]) begin
            sectored_entries_0_4_valid_3 <= 1'h0;
          end else if (_sector_hits_T_29) begin
            if (2'h3 == hitsVec_idx) begin
              sectored_entries_0_4_valid_3 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_15) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_4_valid_3 <= 1'h0;
                    end else begin
                      sectored_entries_0_4_valid_3 <= _GEN_160;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_15) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_4_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_0_4_valid_3 <= _GEN_160;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_29) begin
          if (2'h3 == hitsVec_idx) begin
            sectored_entries_0_4_valid_3 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_15) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_4_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_0_4_valid_3 <= _GEN_160;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_15) begin
                if (invalidate_refill) begin
                  sectored_entries_0_4_valid_3 <= 1'h0;
                end else begin
                  sectored_entries_0_4_valid_3 <= _GEN_160;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_4_valid_3 <= _GEN_736;
      end
    end else begin
      sectored_entries_0_4_valid_3 <= _GEN_516;
    end
    if (metaReset) begin
      sectored_entries_0_5_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_17) begin
            sectored_entries_0_5_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_5_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_17) begin
            if (2'h0 == idx) begin
              sectored_entries_0_5_data_0 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_5_data_1 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_17) begin
            if (2'h1 == idx) begin
              sectored_entries_0_5_data_1 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_5_data_2 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_17) begin
            if (2'h2 == idx) begin
              sectored_entries_0_5_data_2 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_5_data_3 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_17) begin
            if (2'h3 == idx) begin
              sectored_entries_0_5_data_3 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_5_valid_0 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_5_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_754) begin
          if (sectored_entries_0_5_data_0[0]) begin
            sectored_entries_0_5_valid_0 <= 1'h0;
          end else if (_sector_hits_T_35) begin
            if (2'h0 == hitsVec_idx) begin
              sectored_entries_0_5_valid_0 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_17) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_5_valid_0 <= 1'h0;
                    end else begin
                      sectored_entries_0_5_valid_0 <= _GEN_183;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_17) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_5_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_0_5_valid_0 <= _GEN_183;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_35) begin
          if (2'h0 == hitsVec_idx) begin
            sectored_entries_0_5_valid_0 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_17) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_5_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_0_5_valid_0 <= _GEN_183;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_17) begin
                if (invalidate_refill) begin
                  sectored_entries_0_5_valid_0 <= 1'h0;
                end else begin
                  sectored_entries_0_5_valid_0 <= _GEN_183;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_5_valid_0 <= _GEN_761;
      end
    end else begin
      sectored_entries_0_5_valid_0 <= _GEN_523;
    end
    if (metaReset) begin
      sectored_entries_0_5_valid_1 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_5_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_754) begin
          if (sectored_entries_0_5_data_1[0]) begin
            sectored_entries_0_5_valid_1 <= 1'h0;
          end else if (_sector_hits_T_35) begin
            if (2'h1 == hitsVec_idx) begin
              sectored_entries_0_5_valid_1 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_17) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_5_valid_1 <= 1'h0;
                    end else begin
                      sectored_entries_0_5_valid_1 <= _GEN_184;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_17) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_5_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_0_5_valid_1 <= _GEN_184;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_35) begin
          if (2'h1 == hitsVec_idx) begin
            sectored_entries_0_5_valid_1 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_17) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_5_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_0_5_valid_1 <= _GEN_184;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_17) begin
                if (invalidate_refill) begin
                  sectored_entries_0_5_valid_1 <= 1'h0;
                end else begin
                  sectored_entries_0_5_valid_1 <= _GEN_184;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_5_valid_1 <= _GEN_762;
      end
    end else begin
      sectored_entries_0_5_valid_1 <= _GEN_524;
    end
    if (metaReset) begin
      sectored_entries_0_5_valid_2 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_5_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_754) begin
          if (sectored_entries_0_5_data_2[0]) begin
            sectored_entries_0_5_valid_2 <= 1'h0;
          end else if (_sector_hits_T_35) begin
            if (2'h2 == hitsVec_idx) begin
              sectored_entries_0_5_valid_2 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_17) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_5_valid_2 <= 1'h0;
                    end else begin
                      sectored_entries_0_5_valid_2 <= _GEN_185;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_17) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_5_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_0_5_valid_2 <= _GEN_185;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_35) begin
          if (2'h2 == hitsVec_idx) begin
            sectored_entries_0_5_valid_2 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_17) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_5_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_0_5_valid_2 <= _GEN_185;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_17) begin
                if (invalidate_refill) begin
                  sectored_entries_0_5_valid_2 <= 1'h0;
                end else begin
                  sectored_entries_0_5_valid_2 <= _GEN_185;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_5_valid_2 <= _GEN_763;
      end
    end else begin
      sectored_entries_0_5_valid_2 <= _GEN_525;
    end
    if (metaReset) begin
      sectored_entries_0_5_valid_3 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_5_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_754) begin
          if (sectored_entries_0_5_data_3[0]) begin
            sectored_entries_0_5_valid_3 <= 1'h0;
          end else if (_sector_hits_T_35) begin
            if (2'h3 == hitsVec_idx) begin
              sectored_entries_0_5_valid_3 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_17) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_5_valid_3 <= 1'h0;
                    end else begin
                      sectored_entries_0_5_valid_3 <= _GEN_186;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_17) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_5_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_0_5_valid_3 <= _GEN_186;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_35) begin
          if (2'h3 == hitsVec_idx) begin
            sectored_entries_0_5_valid_3 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_17) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_5_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_0_5_valid_3 <= _GEN_186;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_17) begin
                if (invalidate_refill) begin
                  sectored_entries_0_5_valid_3 <= 1'h0;
                end else begin
                  sectored_entries_0_5_valid_3 <= _GEN_186;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_5_valid_3 <= _GEN_764;
      end
    end else begin
      sectored_entries_0_5_valid_3 <= _GEN_526;
    end
    if (metaReset) begin
      sectored_entries_0_6_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_19) begin
            sectored_entries_0_6_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_6_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_19) begin
            if (2'h0 == idx) begin
              sectored_entries_0_6_data_0 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_6_data_1 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_19) begin
            if (2'h1 == idx) begin
              sectored_entries_0_6_data_1 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_6_data_2 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_19) begin
            if (2'h2 == idx) begin
              sectored_entries_0_6_data_2 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_6_data_3 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_19) begin
            if (2'h3 == idx) begin
              sectored_entries_0_6_data_3 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_6_valid_0 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_6_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_893) begin
          if (sectored_entries_0_6_data_0[0]) begin
            sectored_entries_0_6_valid_0 <= 1'h0;
          end else if (_sector_hits_T_41) begin
            if (2'h0 == hitsVec_idx) begin
              sectored_entries_0_6_valid_0 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_19) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_6_valid_0 <= 1'h0;
                    end else begin
                      sectored_entries_0_6_valid_0 <= _GEN_209;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_19) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_6_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_0_6_valid_0 <= _GEN_209;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_41) begin
          if (2'h0 == hitsVec_idx) begin
            sectored_entries_0_6_valid_0 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_19) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_6_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_0_6_valid_0 <= _GEN_209;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_19) begin
                if (invalidate_refill) begin
                  sectored_entries_0_6_valid_0 <= 1'h0;
                end else begin
                  sectored_entries_0_6_valid_0 <= _GEN_209;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_6_valid_0 <= _GEN_789;
      end
    end else begin
      sectored_entries_0_6_valid_0 <= _GEN_533;
    end
    if (metaReset) begin
      sectored_entries_0_6_valid_1 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_6_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_893) begin
          if (sectored_entries_0_6_data_1[0]) begin
            sectored_entries_0_6_valid_1 <= 1'h0;
          end else if (_sector_hits_T_41) begin
            if (2'h1 == hitsVec_idx) begin
              sectored_entries_0_6_valid_1 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_19) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_6_valid_1 <= 1'h0;
                    end else begin
                      sectored_entries_0_6_valid_1 <= _GEN_210;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_19) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_6_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_0_6_valid_1 <= _GEN_210;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_41) begin
          if (2'h1 == hitsVec_idx) begin
            sectored_entries_0_6_valid_1 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_19) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_6_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_0_6_valid_1 <= _GEN_210;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_19) begin
                if (invalidate_refill) begin
                  sectored_entries_0_6_valid_1 <= 1'h0;
                end else begin
                  sectored_entries_0_6_valid_1 <= _GEN_210;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_6_valid_1 <= _GEN_790;
      end
    end else begin
      sectored_entries_0_6_valid_1 <= _GEN_534;
    end
    if (metaReset) begin
      sectored_entries_0_6_valid_2 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_6_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_893) begin
          if (sectored_entries_0_6_data_2[0]) begin
            sectored_entries_0_6_valid_2 <= 1'h0;
          end else if (_sector_hits_T_41) begin
            if (2'h2 == hitsVec_idx) begin
              sectored_entries_0_6_valid_2 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_19) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_6_valid_2 <= 1'h0;
                    end else begin
                      sectored_entries_0_6_valid_2 <= _GEN_211;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_19) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_6_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_0_6_valid_2 <= _GEN_211;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_41) begin
          if (2'h2 == hitsVec_idx) begin
            sectored_entries_0_6_valid_2 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_19) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_6_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_0_6_valid_2 <= _GEN_211;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_19) begin
                if (invalidate_refill) begin
                  sectored_entries_0_6_valid_2 <= 1'h0;
                end else begin
                  sectored_entries_0_6_valid_2 <= _GEN_211;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_6_valid_2 <= _GEN_791;
      end
    end else begin
      sectored_entries_0_6_valid_2 <= _GEN_535;
    end
    if (metaReset) begin
      sectored_entries_0_6_valid_3 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_6_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_893) begin
          if (sectored_entries_0_6_data_3[0]) begin
            sectored_entries_0_6_valid_3 <= 1'h0;
          end else if (_sector_hits_T_41) begin
            if (2'h3 == hitsVec_idx) begin
              sectored_entries_0_6_valid_3 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_19) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_6_valid_3 <= 1'h0;
                    end else begin
                      sectored_entries_0_6_valid_3 <= _GEN_212;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_19) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_6_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_0_6_valid_3 <= _GEN_212;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_41) begin
          if (2'h3 == hitsVec_idx) begin
            sectored_entries_0_6_valid_3 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_19) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_6_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_0_6_valid_3 <= _GEN_212;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_19) begin
                if (invalidate_refill) begin
                  sectored_entries_0_6_valid_3 <= 1'h0;
                end else begin
                  sectored_entries_0_6_valid_3 <= _GEN_212;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_6_valid_3 <= _GEN_792;
      end
    end else begin
      sectored_entries_0_6_valid_3 <= _GEN_536;
    end
    if (metaReset) begin
      sectored_entries_0_7_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_21) begin
            sectored_entries_0_7_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_7_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_21) begin
            if (2'h0 == idx) begin
              sectored_entries_0_7_data_0 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_7_data_1 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_21) begin
            if (2'h1 == idx) begin
              sectored_entries_0_7_data_1 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_7_data_2 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_21) begin
            if (2'h2 == idx) begin
              sectored_entries_0_7_data_2 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_7_data_3 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (!(_T_2)) begin
          if (_T_21) begin
            if (2'h3 == idx) begin
              sectored_entries_0_7_data_3 <= _special_entry_data_0_T;
            end
          end
        end
      end
    end
    if (metaReset) begin
      sectored_entries_0_7_valid_0 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_7_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_1032) begin
          if (sectored_entries_0_7_data_0[0]) begin
            sectored_entries_0_7_valid_0 <= 1'h0;
          end else if (_sector_hits_T_47) begin
            if (2'h0 == hitsVec_idx) begin
              sectored_entries_0_7_valid_0 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_21) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_7_valid_0 <= 1'h0;
                    end else begin
                      sectored_entries_0_7_valid_0 <= _GEN_235;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_21) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_7_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_0_7_valid_0 <= _GEN_235;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_47) begin
          if (2'h0 == hitsVec_idx) begin
            sectored_entries_0_7_valid_0 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_21) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_7_valid_0 <= 1'h0;
                  end else begin
                    sectored_entries_0_7_valid_0 <= _GEN_235;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_21) begin
                if (invalidate_refill) begin
                  sectored_entries_0_7_valid_0 <= 1'h0;
                end else begin
                  sectored_entries_0_7_valid_0 <= _GEN_235;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_7_valid_0 <= _GEN_817;
      end
    end else begin
      sectored_entries_0_7_valid_0 <= _GEN_543;
    end
    if (metaReset) begin
      sectored_entries_0_7_valid_1 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_7_valid_1 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_1032) begin
          if (sectored_entries_0_7_data_1[0]) begin
            sectored_entries_0_7_valid_1 <= 1'h0;
          end else if (_sector_hits_T_47) begin
            if (2'h1 == hitsVec_idx) begin
              sectored_entries_0_7_valid_1 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_21) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_7_valid_1 <= 1'h0;
                    end else begin
                      sectored_entries_0_7_valid_1 <= _GEN_236;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_21) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_7_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_0_7_valid_1 <= _GEN_236;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_47) begin
          if (2'h1 == hitsVec_idx) begin
            sectored_entries_0_7_valid_1 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_21) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_7_valid_1 <= 1'h0;
                  end else begin
                    sectored_entries_0_7_valid_1 <= _GEN_236;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_21) begin
                if (invalidate_refill) begin
                  sectored_entries_0_7_valid_1 <= 1'h0;
                end else begin
                  sectored_entries_0_7_valid_1 <= _GEN_236;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_7_valid_1 <= _GEN_818;
      end
    end else begin
      sectored_entries_0_7_valid_1 <= _GEN_544;
    end
    if (metaReset) begin
      sectored_entries_0_7_valid_2 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_7_valid_2 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_1032) begin
          if (sectored_entries_0_7_data_2[0]) begin
            sectored_entries_0_7_valid_2 <= 1'h0;
          end else if (_sector_hits_T_47) begin
            if (2'h2 == hitsVec_idx) begin
              sectored_entries_0_7_valid_2 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_21) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_7_valid_2 <= 1'h0;
                    end else begin
                      sectored_entries_0_7_valid_2 <= _GEN_237;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_21) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_7_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_0_7_valid_2 <= _GEN_237;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_47) begin
          if (2'h2 == hitsVec_idx) begin
            sectored_entries_0_7_valid_2 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_21) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_7_valid_2 <= 1'h0;
                  end else begin
                    sectored_entries_0_7_valid_2 <= _GEN_237;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_21) begin
                if (invalidate_refill) begin
                  sectored_entries_0_7_valid_2 <= 1'h0;
                end else begin
                  sectored_entries_0_7_valid_2 <= _GEN_237;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_7_valid_2 <= _GEN_819;
      end
    end else begin
      sectored_entries_0_7_valid_2 <= _GEN_545;
    end
    if (metaReset) begin
      sectored_entries_0_7_valid_3 <= 1'h0;
    end else if (_T_1326) begin
      sectored_entries_0_7_valid_3 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_T_1032) begin
          if (sectored_entries_0_7_data_3[0]) begin
            sectored_entries_0_7_valid_3 <= 1'h0;
          end else if (_sector_hits_T_47) begin
            if (2'h3 == hitsVec_idx) begin
              sectored_entries_0_7_valid_3 <= 1'h0;
            end else if (io_ptw_resp_valid) begin
              if (!(~io_ptw_resp_bits_homogeneous)) begin
                if (!(_T_2)) begin
                  if (_T_21) begin
                    if (invalidate_refill) begin
                      sectored_entries_0_7_valid_3 <= 1'h0;
                    end else begin
                      sectored_entries_0_7_valid_3 <= _GEN_238;
                    end
                  end
                end
              end
            end
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_21) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_7_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_0_7_valid_3 <= _GEN_238;
                  end
                end
              end
            end
          end
        end else if (_sector_hits_T_47) begin
          if (2'h3 == hitsVec_idx) begin
            sectored_entries_0_7_valid_3 <= 1'h0;
          end else if (io_ptw_resp_valid) begin
            if (!(~io_ptw_resp_bits_homogeneous)) begin
              if (!(_T_2)) begin
                if (_T_21) begin
                  if (invalidate_refill) begin
                    sectored_entries_0_7_valid_3 <= 1'h0;
                  end else begin
                    sectored_entries_0_7_valid_3 <= _GEN_238;
                  end
                end
              end
            end
          end
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (!(_T_2)) begin
              if (_T_21) begin
                if (invalidate_refill) begin
                  sectored_entries_0_7_valid_3 <= 1'h0;
                end else begin
                  sectored_entries_0_7_valid_3 <= _GEN_238;
                end
              end
            end
          end
        end
      end else begin
        sectored_entries_0_7_valid_3 <= _GEN_820;
      end
    end else begin
      sectored_entries_0_7_valid_3 <= _GEN_546;
    end
    if (metaReset) begin
      superpage_entries_0_level <= 2'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_2) begin
          if (_T_3) begin
            superpage_entries_0_level <= {{1'd0}, io_ptw_resp_bits_level[0]};
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_0_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_2) begin
          if (_T_3) begin
            superpage_entries_0_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_0_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_2) begin
          if (_T_3) begin
            superpage_entries_0_data_0 <= _special_entry_data_0_T;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_0_valid_0 <= 1'h0;
    end else if (_T_1326) begin
      superpage_entries_0_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (superpage_hits_0) begin
          superpage_entries_0_valid_0 <= 1'h0;
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (_T_2) begin
              if (_T_3) begin
                if (invalidate_refill) begin
                  superpage_entries_0_valid_0 <= 1'h0;
                end else begin
                  superpage_entries_0_valid_0 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        superpage_entries_0_valid_0 <= _GEN_827;
      end
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_2) begin
          if (_T_3) begin
            if (invalidate_refill) begin
              superpage_entries_0_valid_0 <= 1'h0;
            end else begin
              superpage_entries_0_valid_0 <= 1'h1;
            end
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_1_level <= 2'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_2) begin
          if (_T_4) begin
            superpage_entries_1_level <= {{1'd0}, io_ptw_resp_bits_level[0]};
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_1_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_2) begin
          if (_T_4) begin
            superpage_entries_1_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_1_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_2) begin
          if (_T_4) begin
            superpage_entries_1_data_0 <= _special_entry_data_0_T;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_1_valid_0 <= 1'h0;
    end else if (_T_1326) begin
      superpage_entries_1_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (superpage_hits_1) begin
          superpage_entries_1_valid_0 <= 1'h0;
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (_T_2) begin
              if (_T_4) begin
                if (invalidate_refill) begin
                  superpage_entries_1_valid_0 <= 1'h0;
                end else begin
                  superpage_entries_1_valid_0 <= 1'h1;
                end
              end
            end
          end
        end
      end else begin
        superpage_entries_1_valid_0 <= _GEN_831;
      end
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_2) begin
          if (_T_4) begin
            if (invalidate_refill) begin
              superpage_entries_1_valid_0 <= 1'h0;
            end else begin
              superpage_entries_1_valid_0 <= 1'h1;
            end
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_2_level <= 2'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_2) begin
          if (_T_5) begin
            superpage_entries_2_level <= {{1'd0}, io_ptw_resp_bits_level[0]};
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_2_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_2) begin
          if (_T_5) begin
            superpage_entries_2_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_2_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_2) begin
          if (_T_5) begin
            superpage_entries_2_data_0 <= _special_entry_data_0_T;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_2_valid_0 <= 1'h0;
    end else if (_T_1326) begin
      superpage_entries_2_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (superpage_hits_2) begin
          superpage_entries_2_valid_0 <= 1'h0;
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (_T_2) begin
              if (_T_5) begin
                superpage_entries_2_valid_0 <= _GEN_32;
              end
            end
          end
        end
      end else begin
        superpage_entries_2_valid_0 <= _GEN_835;
      end
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_2) begin
          if (_T_5) begin
            superpage_entries_2_valid_0 <= _GEN_32;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_3_level <= 2'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_2) begin
          if (_T_6) begin
            superpage_entries_3_level <= {{1'd0}, io_ptw_resp_bits_level[0]};
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_3_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_2) begin
          if (_T_6) begin
            superpage_entries_3_tag <= r_refill_tag;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_3_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_2) begin
          if (_T_6) begin
            superpage_entries_3_data_0 <= _special_entry_data_0_T;
          end
        end
      end
    end
    if (metaReset) begin
      superpage_entries_3_valid_0 <= 1'h0;
    end else if (_T_1326) begin
      superpage_entries_3_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (superpage_hits_3) begin
          superpage_entries_3_valid_0 <= 1'h0;
        end else if (io_ptw_resp_valid) begin
          if (!(~io_ptw_resp_bits_homogeneous)) begin
            if (_T_2) begin
              if (_T_6) begin
                superpage_entries_3_valid_0 <= _GEN_32;
              end
            end
          end
        end
      end else begin
        superpage_entries_3_valid_0 <= _GEN_839;
      end
    end else if (io_ptw_resp_valid) begin
      if (!(~io_ptw_resp_bits_homogeneous)) begin
        if (_T_2) begin
          if (_T_6) begin
            superpage_entries_3_valid_0 <= _GEN_32;
          end
        end
      end
    end
    if (metaReset) begin
      special_entry_level <= 2'h0;
    end else if (io_ptw_resp_valid) begin
      if (~io_ptw_resp_bits_homogeneous) begin
        special_entry_level <= io_ptw_resp_bits_level;
      end
    end
    if (metaReset) begin
      special_entry_tag <= 27'h0;
    end else if (io_ptw_resp_valid) begin
      if (~io_ptw_resp_bits_homogeneous) begin
        special_entry_tag <= r_refill_tag;
      end
    end
    if (metaReset) begin
      special_entry_data_0 <= 35'h0;
    end else if (io_ptw_resp_valid) begin
      if (~io_ptw_resp_bits_homogeneous) begin
        special_entry_data_0 <= _special_entry_data_0_T;
      end
    end
    if (metaReset) begin
      special_entry_valid_0 <= 1'h0;
    end else if (_T_1326) begin
      special_entry_valid_0 <= 1'h0;
    end else if (io_sfence_valid) begin
      if (io_sfence_bits_rs1) begin
        if (_hitsVec_T_106) begin
          special_entry_valid_0 <= 1'h0;
        end else if (io_ptw_resp_valid) begin
          if (~io_ptw_resp_bits_homogeneous) begin
            special_entry_valid_0 <= _GEN_32;
          end
        end
      end else begin
        special_entry_valid_0 <= _GEN_843;
      end
    end else if (io_ptw_resp_valid) begin
      if (~io_ptw_resp_bits_homogeneous) begin
        special_entry_valid_0 <= _GEN_32;
      end
    end
    if (metaReset) begin
      state <= 2'h0;
    end else if (reset) begin
      state <= 2'h0;
    end else if (io_ptw_resp_valid) begin
      state <= 2'h0;
    end else if (_T_45) begin
      state <= 2'h3;
    end else if (_invalidate_refill_T) begin
      if (io_kill) begin
        state <= 2'h0;
      end else if (io_ptw_req_ready) begin
        if (io_sfence_valid) begin
          state <= 2'h3;
        end else begin
          state <= 2'h2;
        end
      end else if (io_sfence_valid) begin
        state <= 2'h0;
      end else if (_T_42) begin
        state <= 2'h1;
      end
    end else if (_T_42) begin
      state <= 2'h1;
    end
    if (metaReset) begin
      r_refill_tag <= 27'h0;
    end else if (_T_42) begin
      r_refill_tag <= vpn;
    end
    if (metaReset) begin
      r_superpage_repl_addr <= 2'h0;
    end else if (_T_42) begin
      if (_r_superpage_repl_addr_T_3) begin
        r_superpage_repl_addr <= _r_superpage_repl_addr_T_2;
      end else if (_r_superpage_repl_addr_T_5) begin
        r_superpage_repl_addr <= 2'h0;
      end else if (_r_superpage_repl_addr_T_6) begin
        r_superpage_repl_addr <= 2'h1;
      end else if (_r_superpage_repl_addr_T_7) begin
        r_superpage_repl_addr <= 2'h2;
      end else begin
        r_superpage_repl_addr <= 2'h3;
      end
    end
    if (metaReset) begin
      r_sectored_repl_addr <= 3'h0;
    end else if (_T_42) begin
      if (_r_sectored_repl_addr_T_7) begin
        r_sectored_repl_addr <= _r_sectored_repl_addr_T_6;
      end else if (_r_sectored_repl_addr_T_9) begin
        r_sectored_repl_addr <= 3'h0;
      end else if (_r_sectored_repl_addr_T_10) begin
        r_sectored_repl_addr <= 3'h1;
      end else if (_r_sectored_repl_addr_T_11) begin
        r_sectored_repl_addr <= 3'h2;
      end else if (_r_sectored_repl_addr_T_12) begin
        r_sectored_repl_addr <= 3'h3;
      end else if (_r_sectored_repl_addr_T_13) begin
        r_sectored_repl_addr <= 3'h4;
      end else if (_r_sectored_repl_addr_T_14) begin
        r_sectored_repl_addr <= 3'h5;
      end else if (_r_sectored_repl_addr_T_15) begin
        r_sectored_repl_addr <= 3'h6;
      end else begin
        r_sectored_repl_addr <= 3'h7;
      end
    end
    if (metaReset) begin
      r_sectored_hit_addr <= 3'h0;
    end else if (_T_42) begin
      r_sectored_hit_addr <= state_vec_0_touch_way_sized;
    end
    if (metaReset) begin
      r_sectored_hit <= 1'h0;
    end else if (_T_42) begin
      r_sectored_hit <= _T_30;
    end
    if (metaReset) begin
      state_vec_0 <= 7'h0;
    end else if (reset) begin
      state_vec_0 <= 7'h0;
    end else if (_T_23) begin
      if (_T_30) begin
        state_vec_0 <= _state_vec_0_T_16;
      end
    end
    if (metaReset) begin
      state_reg_1 <= 3'h0;
    end else if (reset) begin
      state_reg_1 <= 3'h0;
    end else if (_T_23) begin
      if (_T_37) begin
        state_reg_1 <= _state_reg_T_6;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_sfence_valid & ~_T_51) begin
          $fwrite(32'h80000002,"Assertion failed\n    at TLB.scala:385 assert(!io.sfence.bits.rs1 || (io.sfence.bits.addr >> pgIdxBits) === vpn)\n"); // @[TLB.scala 385:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_sfence_valid & ~_T_51) begin
          $fatal; // @[TLB.scala 385:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    TLB_1_state <= TLB_1_xor0;
    if (!(TLB_1_cov_read_data)) begin
      TLB_1_covSum <= TLB_1_covSum + 1'h1;
    end
    if (metaReset) begin
      TLB_1_metaAssert <= 1'h0;
    end else begin
      TLB_1_metaAssert <= TLB_1_metaAssert | TLB_1_or0;
    end
  end
  always @(posedge clock) begin
    if(TLB_1_cov_write_en & TLB_1_cov_write_mask) begin
      TLB_1_cov[TLB_1_cov_write_addr] <= TLB_1_cov_write_data; // @[Coverage map for TLB_1]
    end
  end
endmodule
module BTB(
  input         clock,
  input         reset,
  input  [38:0] io_req_bits_addr,
  output        io_resp_valid,
  output        io_resp_bits_taken,
  output        io_resp_bits_bridx,
  output [38:0] io_resp_bits_target,
  output [4:0]  io_resp_bits_entry,
  output [7:0]  io_resp_bits_bht_history,
  output        io_resp_bits_bht_value,
  input         io_btb_update_valid,
  input  [4:0]  io_btb_update_bits_prediction_entry,
  input  [38:0] io_btb_update_bits_pc,
  input         io_btb_update_bits_isValid,
  input  [38:0] io_btb_update_bits_br_pc,
  input  [1:0]  io_btb_update_bits_cfiType,
  input         io_bht_update_valid,
  input  [7:0]  io_bht_update_bits_prediction_history,
  input  [38:0] io_bht_update_bits_pc,
  input         io_bht_update_bits_branch,
  input         io_bht_update_bits_taken,
  input         io_bht_update_bits_mispredict,
  input         io_bht_advance_valid,
  input         io_bht_advance_bits_bht_value,
  input         io_ras_update_valid,
  input  [1:0]  io_ras_update_bits_cfiType,
  input  [38:0] io_ras_update_bits_returnAddr,
  output        io_ras_head_valid,
  output [38:0] io_ras_head_bits,
  input         io_flush,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  reg  table_ [0:511]; // @[BTB.scala 118:26]
  reg [31:0] _RAND_0;
  wire  table__res_res_value_MPORT_data; // @[BTB.scala 118:26]
  wire [8:0] table__res_res_value_MPORT_addr; // @[BTB.scala 118:26]
  wire  table__MPORT_data; // @[BTB.scala 118:26]
  wire [8:0] table__MPORT_addr; // @[BTB.scala 118:26]
  wire  table__MPORT_mask; // @[BTB.scala 118:26]
  wire  table__MPORT_en; // @[BTB.scala 118:26]
  reg [12:0] idxs_0; // @[BTB.scala 201:17]
  reg [31:0] _RAND_1;
  reg [12:0] idxs_1; // @[BTB.scala 201:17]
  reg [31:0] _RAND_2;
  reg [12:0] idxs_2; // @[BTB.scala 201:17]
  reg [31:0] _RAND_3;
  reg [12:0] idxs_3; // @[BTB.scala 201:17]
  reg [31:0] _RAND_4;
  reg [12:0] idxs_4; // @[BTB.scala 201:17]
  reg [31:0] _RAND_5;
  reg [12:0] idxs_5; // @[BTB.scala 201:17]
  reg [31:0] _RAND_6;
  reg [12:0] idxs_6; // @[BTB.scala 201:17]
  reg [31:0] _RAND_7;
  reg [12:0] idxs_7; // @[BTB.scala 201:17]
  reg [31:0] _RAND_8;
  reg [12:0] idxs_8; // @[BTB.scala 201:17]
  reg [31:0] _RAND_9;
  reg [12:0] idxs_9; // @[BTB.scala 201:17]
  reg [31:0] _RAND_10;
  reg [12:0] idxs_10; // @[BTB.scala 201:17]
  reg [31:0] _RAND_11;
  reg [12:0] idxs_11; // @[BTB.scala 201:17]
  reg [31:0] _RAND_12;
  reg [12:0] idxs_12; // @[BTB.scala 201:17]
  reg [31:0] _RAND_13;
  reg [12:0] idxs_13; // @[BTB.scala 201:17]
  reg [31:0] _RAND_14;
  reg [12:0] idxs_14; // @[BTB.scala 201:17]
  reg [31:0] _RAND_15;
  reg [12:0] idxs_15; // @[BTB.scala 201:17]
  reg [31:0] _RAND_16;
  reg [12:0] idxs_16; // @[BTB.scala 201:17]
  reg [31:0] _RAND_17;
  reg [12:0] idxs_17; // @[BTB.scala 201:17]
  reg [31:0] _RAND_18;
  reg [12:0] idxs_18; // @[BTB.scala 201:17]
  reg [31:0] _RAND_19;
  reg [12:0] idxs_19; // @[BTB.scala 201:17]
  reg [31:0] _RAND_20;
  reg [12:0] idxs_20; // @[BTB.scala 201:17]
  reg [31:0] _RAND_21;
  reg [12:0] idxs_21; // @[BTB.scala 201:17]
  reg [31:0] _RAND_22;
  reg [12:0] idxs_22; // @[BTB.scala 201:17]
  reg [31:0] _RAND_23;
  reg [12:0] idxs_23; // @[BTB.scala 201:17]
  reg [31:0] _RAND_24;
  reg [12:0] idxs_24; // @[BTB.scala 201:17]
  reg [31:0] _RAND_25;
  reg [12:0] idxs_25; // @[BTB.scala 201:17]
  reg [31:0] _RAND_26;
  reg [12:0] idxs_26; // @[BTB.scala 201:17]
  reg [31:0] _RAND_27;
  reg [12:0] idxs_27; // @[BTB.scala 201:17]
  reg [31:0] _RAND_28;
  reg [2:0] idxPages_0; // @[BTB.scala 202:21]
  reg [31:0] _RAND_29;
  reg [2:0] idxPages_1; // @[BTB.scala 202:21]
  reg [31:0] _RAND_30;
  reg [2:0] idxPages_2; // @[BTB.scala 202:21]
  reg [31:0] _RAND_31;
  reg [2:0] idxPages_3; // @[BTB.scala 202:21]
  reg [31:0] _RAND_32;
  reg [2:0] idxPages_4; // @[BTB.scala 202:21]
  reg [31:0] _RAND_33;
  reg [2:0] idxPages_5; // @[BTB.scala 202:21]
  reg [31:0] _RAND_34;
  reg [2:0] idxPages_6; // @[BTB.scala 202:21]
  reg [31:0] _RAND_35;
  reg [2:0] idxPages_7; // @[BTB.scala 202:21]
  reg [31:0] _RAND_36;
  reg [2:0] idxPages_8; // @[BTB.scala 202:21]
  reg [31:0] _RAND_37;
  reg [2:0] idxPages_9; // @[BTB.scala 202:21]
  reg [31:0] _RAND_38;
  reg [2:0] idxPages_10; // @[BTB.scala 202:21]
  reg [31:0] _RAND_39;
  reg [2:0] idxPages_11; // @[BTB.scala 202:21]
  reg [31:0] _RAND_40;
  reg [2:0] idxPages_12; // @[BTB.scala 202:21]
  reg [31:0] _RAND_41;
  reg [2:0] idxPages_13; // @[BTB.scala 202:21]
  reg [31:0] _RAND_42;
  reg [2:0] idxPages_14; // @[BTB.scala 202:21]
  reg [31:0] _RAND_43;
  reg [2:0] idxPages_15; // @[BTB.scala 202:21]
  reg [31:0] _RAND_44;
  reg [2:0] idxPages_16; // @[BTB.scala 202:21]
  reg [31:0] _RAND_45;
  reg [2:0] idxPages_17; // @[BTB.scala 202:21]
  reg [31:0] _RAND_46;
  reg [2:0] idxPages_18; // @[BTB.scala 202:21]
  reg [31:0] _RAND_47;
  reg [2:0] idxPages_19; // @[BTB.scala 202:21]
  reg [31:0] _RAND_48;
  reg [2:0] idxPages_20; // @[BTB.scala 202:21]
  reg [31:0] _RAND_49;
  reg [2:0] idxPages_21; // @[BTB.scala 202:21]
  reg [31:0] _RAND_50;
  reg [2:0] idxPages_22; // @[BTB.scala 202:21]
  reg [31:0] _RAND_51;
  reg [2:0] idxPages_23; // @[BTB.scala 202:21]
  reg [31:0] _RAND_52;
  reg [2:0] idxPages_24; // @[BTB.scala 202:21]
  reg [31:0] _RAND_53;
  reg [2:0] idxPages_25; // @[BTB.scala 202:21]
  reg [31:0] _RAND_54;
  reg [2:0] idxPages_26; // @[BTB.scala 202:21]
  reg [31:0] _RAND_55;
  reg [2:0] idxPages_27; // @[BTB.scala 202:21]
  reg [31:0] _RAND_56;
  reg [12:0] tgts_0; // @[BTB.scala 203:17]
  reg [31:0] _RAND_57;
  reg [12:0] tgts_1; // @[BTB.scala 203:17]
  reg [31:0] _RAND_58;
  reg [12:0] tgts_2; // @[BTB.scala 203:17]
  reg [31:0] _RAND_59;
  reg [12:0] tgts_3; // @[BTB.scala 203:17]
  reg [31:0] _RAND_60;
  reg [12:0] tgts_4; // @[BTB.scala 203:17]
  reg [31:0] _RAND_61;
  reg [12:0] tgts_5; // @[BTB.scala 203:17]
  reg [31:0] _RAND_62;
  reg [12:0] tgts_6; // @[BTB.scala 203:17]
  reg [31:0] _RAND_63;
  reg [12:0] tgts_7; // @[BTB.scala 203:17]
  reg [31:0] _RAND_64;
  reg [12:0] tgts_8; // @[BTB.scala 203:17]
  reg [31:0] _RAND_65;
  reg [12:0] tgts_9; // @[BTB.scala 203:17]
  reg [31:0] _RAND_66;
  reg [12:0] tgts_10; // @[BTB.scala 203:17]
  reg [31:0] _RAND_67;
  reg [12:0] tgts_11; // @[BTB.scala 203:17]
  reg [31:0] _RAND_68;
  reg [12:0] tgts_12; // @[BTB.scala 203:17]
  reg [31:0] _RAND_69;
  reg [12:0] tgts_13; // @[BTB.scala 203:17]
  reg [31:0] _RAND_70;
  reg [12:0] tgts_14; // @[BTB.scala 203:17]
  reg [31:0] _RAND_71;
  reg [12:0] tgts_15; // @[BTB.scala 203:17]
  reg [31:0] _RAND_72;
  reg [12:0] tgts_16; // @[BTB.scala 203:17]
  reg [31:0] _RAND_73;
  reg [12:0] tgts_17; // @[BTB.scala 203:17]
  reg [31:0] _RAND_74;
  reg [12:0] tgts_18; // @[BTB.scala 203:17]
  reg [31:0] _RAND_75;
  reg [12:0] tgts_19; // @[BTB.scala 203:17]
  reg [31:0] _RAND_76;
  reg [12:0] tgts_20; // @[BTB.scala 203:17]
  reg [31:0] _RAND_77;
  reg [12:0] tgts_21; // @[BTB.scala 203:17]
  reg [31:0] _RAND_78;
  reg [12:0] tgts_22; // @[BTB.scala 203:17]
  reg [31:0] _RAND_79;
  reg [12:0] tgts_23; // @[BTB.scala 203:17]
  reg [31:0] _RAND_80;
  reg [12:0] tgts_24; // @[BTB.scala 203:17]
  reg [31:0] _RAND_81;
  reg [12:0] tgts_25; // @[BTB.scala 203:17]
  reg [31:0] _RAND_82;
  reg [12:0] tgts_26; // @[BTB.scala 203:17]
  reg [31:0] _RAND_83;
  reg [12:0] tgts_27; // @[BTB.scala 203:17]
  reg [31:0] _RAND_84;
  reg [2:0] tgtPages_0; // @[BTB.scala 204:21]
  reg [31:0] _RAND_85;
  reg [2:0] tgtPages_1; // @[BTB.scala 204:21]
  reg [31:0] _RAND_86;
  reg [2:0] tgtPages_2; // @[BTB.scala 204:21]
  reg [31:0] _RAND_87;
  reg [2:0] tgtPages_3; // @[BTB.scala 204:21]
  reg [31:0] _RAND_88;
  reg [2:0] tgtPages_4; // @[BTB.scala 204:21]
  reg [31:0] _RAND_89;
  reg [2:0] tgtPages_5; // @[BTB.scala 204:21]
  reg [31:0] _RAND_90;
  reg [2:0] tgtPages_6; // @[BTB.scala 204:21]
  reg [31:0] _RAND_91;
  reg [2:0] tgtPages_7; // @[BTB.scala 204:21]
  reg [31:0] _RAND_92;
  reg [2:0] tgtPages_8; // @[BTB.scala 204:21]
  reg [31:0] _RAND_93;
  reg [2:0] tgtPages_9; // @[BTB.scala 204:21]
  reg [31:0] _RAND_94;
  reg [2:0] tgtPages_10; // @[BTB.scala 204:21]
  reg [31:0] _RAND_95;
  reg [2:0] tgtPages_11; // @[BTB.scala 204:21]
  reg [31:0] _RAND_96;
  reg [2:0] tgtPages_12; // @[BTB.scala 204:21]
  reg [31:0] _RAND_97;
  reg [2:0] tgtPages_13; // @[BTB.scala 204:21]
  reg [31:0] _RAND_98;
  reg [2:0] tgtPages_14; // @[BTB.scala 204:21]
  reg [31:0] _RAND_99;
  reg [2:0] tgtPages_15; // @[BTB.scala 204:21]
  reg [31:0] _RAND_100;
  reg [2:0] tgtPages_16; // @[BTB.scala 204:21]
  reg [31:0] _RAND_101;
  reg [2:0] tgtPages_17; // @[BTB.scala 204:21]
  reg [31:0] _RAND_102;
  reg [2:0] tgtPages_18; // @[BTB.scala 204:21]
  reg [31:0] _RAND_103;
  reg [2:0] tgtPages_19; // @[BTB.scala 204:21]
  reg [31:0] _RAND_104;
  reg [2:0] tgtPages_20; // @[BTB.scala 204:21]
  reg [31:0] _RAND_105;
  reg [2:0] tgtPages_21; // @[BTB.scala 204:21]
  reg [31:0] _RAND_106;
  reg [2:0] tgtPages_22; // @[BTB.scala 204:21]
  reg [31:0] _RAND_107;
  reg [2:0] tgtPages_23; // @[BTB.scala 204:21]
  reg [31:0] _RAND_108;
  reg [2:0] tgtPages_24; // @[BTB.scala 204:21]
  reg [31:0] _RAND_109;
  reg [2:0] tgtPages_25; // @[BTB.scala 204:21]
  reg [31:0] _RAND_110;
  reg [2:0] tgtPages_26; // @[BTB.scala 204:21]
  reg [31:0] _RAND_111;
  reg [2:0] tgtPages_27; // @[BTB.scala 204:21]
  reg [31:0] _RAND_112;
  reg [24:0] pages_0; // @[BTB.scala 205:18]
  reg [31:0] _RAND_113;
  reg [24:0] pages_1; // @[BTB.scala 205:18]
  reg [31:0] _RAND_114;
  reg [24:0] pages_2; // @[BTB.scala 205:18]
  reg [31:0] _RAND_115;
  reg [24:0] pages_3; // @[BTB.scala 205:18]
  reg [31:0] _RAND_116;
  reg [24:0] pages_4; // @[BTB.scala 205:18]
  reg [31:0] _RAND_117;
  reg [24:0] pages_5; // @[BTB.scala 205:18]
  reg [31:0] _RAND_118;
  reg [5:0] pageValid; // @[BTB.scala 206:22]
  reg [31:0] _RAND_119;
  wire [24:0] pagesMasked_0; // @[BTB.scala 207:75]
  wire [24:0] pagesMasked_1; // @[BTB.scala 207:75]
  wire [24:0] pagesMasked_2; // @[BTB.scala 207:75]
  wire [24:0] pagesMasked_3; // @[BTB.scala 207:75]
  wire [24:0] pagesMasked_4; // @[BTB.scala 207:75]
  wire [24:0] pagesMasked_5; // @[BTB.scala 207:75]
  reg [27:0] isValid; // @[BTB.scala 209:20]
  reg [31:0] _RAND_120;
  reg [1:0] cfiType_0; // @[BTB.scala 210:20]
  reg [31:0] _RAND_121;
  reg [1:0] cfiType_1; // @[BTB.scala 210:20]
  reg [31:0] _RAND_122;
  reg [1:0] cfiType_2; // @[BTB.scala 210:20]
  reg [31:0] _RAND_123;
  reg [1:0] cfiType_3; // @[BTB.scala 210:20]
  reg [31:0] _RAND_124;
  reg [1:0] cfiType_4; // @[BTB.scala 210:20]
  reg [31:0] _RAND_125;
  reg [1:0] cfiType_5; // @[BTB.scala 210:20]
  reg [31:0] _RAND_126;
  reg [1:0] cfiType_6; // @[BTB.scala 210:20]
  reg [31:0] _RAND_127;
  reg [1:0] cfiType_7; // @[BTB.scala 210:20]
  reg [31:0] _RAND_128;
  reg [1:0] cfiType_8; // @[BTB.scala 210:20]
  reg [31:0] _RAND_129;
  reg [1:0] cfiType_9; // @[BTB.scala 210:20]
  reg [31:0] _RAND_130;
  reg [1:0] cfiType_10; // @[BTB.scala 210:20]
  reg [31:0] _RAND_131;
  reg [1:0] cfiType_11; // @[BTB.scala 210:20]
  reg [31:0] _RAND_132;
  reg [1:0] cfiType_12; // @[BTB.scala 210:20]
  reg [31:0] _RAND_133;
  reg [1:0] cfiType_13; // @[BTB.scala 210:20]
  reg [31:0] _RAND_134;
  reg [1:0] cfiType_14; // @[BTB.scala 210:20]
  reg [31:0] _RAND_135;
  reg [1:0] cfiType_15; // @[BTB.scala 210:20]
  reg [31:0] _RAND_136;
  reg [1:0] cfiType_16; // @[BTB.scala 210:20]
  reg [31:0] _RAND_137;
  reg [1:0] cfiType_17; // @[BTB.scala 210:20]
  reg [31:0] _RAND_138;
  reg [1:0] cfiType_18; // @[BTB.scala 210:20]
  reg [31:0] _RAND_139;
  reg [1:0] cfiType_19; // @[BTB.scala 210:20]
  reg [31:0] _RAND_140;
  reg [1:0] cfiType_20; // @[BTB.scala 210:20]
  reg [31:0] _RAND_141;
  reg [1:0] cfiType_21; // @[BTB.scala 210:20]
  reg [31:0] _RAND_142;
  reg [1:0] cfiType_22; // @[BTB.scala 210:20]
  reg [31:0] _RAND_143;
  reg [1:0] cfiType_23; // @[BTB.scala 210:20]
  reg [31:0] _RAND_144;
  reg [1:0] cfiType_24; // @[BTB.scala 210:20]
  reg [31:0] _RAND_145;
  reg [1:0] cfiType_25; // @[BTB.scala 210:20]
  reg [31:0] _RAND_146;
  reg [1:0] cfiType_26; // @[BTB.scala 210:20]
  reg [31:0] _RAND_147;
  reg [1:0] cfiType_27; // @[BTB.scala 210:20]
  reg [31:0] _RAND_148;
  reg  brIdx_0; // @[BTB.scala 211:18]
  reg [31:0] _RAND_149;
  reg  brIdx_1; // @[BTB.scala 211:18]
  reg [31:0] _RAND_150;
  reg  brIdx_2; // @[BTB.scala 211:18]
  reg [31:0] _RAND_151;
  reg  brIdx_3; // @[BTB.scala 211:18]
  reg [31:0] _RAND_152;
  reg  brIdx_4; // @[BTB.scala 211:18]
  reg [31:0] _RAND_153;
  reg  brIdx_5; // @[BTB.scala 211:18]
  reg [31:0] _RAND_154;
  reg  brIdx_6; // @[BTB.scala 211:18]
  reg [31:0] _RAND_155;
  reg  brIdx_7; // @[BTB.scala 211:18]
  reg [31:0] _RAND_156;
  reg  brIdx_8; // @[BTB.scala 211:18]
  reg [31:0] _RAND_157;
  reg  brIdx_9; // @[BTB.scala 211:18]
  reg [31:0] _RAND_158;
  reg  brIdx_10; // @[BTB.scala 211:18]
  reg [31:0] _RAND_159;
  reg  brIdx_11; // @[BTB.scala 211:18]
  reg [31:0] _RAND_160;
  reg  brIdx_12; // @[BTB.scala 211:18]
  reg [31:0] _RAND_161;
  reg  brIdx_13; // @[BTB.scala 211:18]
  reg [31:0] _RAND_162;
  reg  brIdx_14; // @[BTB.scala 211:18]
  reg [31:0] _RAND_163;
  reg  brIdx_15; // @[BTB.scala 211:18]
  reg [31:0] _RAND_164;
  reg  brIdx_16; // @[BTB.scala 211:18]
  reg [31:0] _RAND_165;
  reg  brIdx_17; // @[BTB.scala 211:18]
  reg [31:0] _RAND_166;
  reg  brIdx_18; // @[BTB.scala 211:18]
  reg [31:0] _RAND_167;
  reg  brIdx_19; // @[BTB.scala 211:18]
  reg [31:0] _RAND_168;
  reg  brIdx_20; // @[BTB.scala 211:18]
  reg [31:0] _RAND_169;
  reg  brIdx_21; // @[BTB.scala 211:18]
  reg [31:0] _RAND_170;
  reg  brIdx_22; // @[BTB.scala 211:18]
  reg [31:0] _RAND_171;
  reg  brIdx_23; // @[BTB.scala 211:18]
  reg [31:0] _RAND_172;
  reg  brIdx_24; // @[BTB.scala 211:18]
  reg [31:0] _RAND_173;
  reg  brIdx_25; // @[BTB.scala 211:18]
  reg [31:0] _RAND_174;
  reg  brIdx_26; // @[BTB.scala 211:18]
  reg [31:0] _RAND_175;
  reg  brIdx_27; // @[BTB.scala 211:18]
  reg [31:0] _RAND_176;
  reg  r_btb_updatePipe_valid; // @[Valid.scala 117:22]
  reg [31:0] _RAND_177;
  reg [4:0] r_btb_updatePipe_bits_prediction_entry; // @[Reg.scala 15:16]
  reg [31:0] _RAND_178;
  reg [38:0] r_btb_updatePipe_bits_pc; // @[Reg.scala 15:16]
  reg [63:0] _RAND_179;
  reg  r_btb_updatePipe_bits_isValid; // @[Reg.scala 15:16]
  reg [31:0] _RAND_180;
  reg [38:0] r_btb_updatePipe_bits_br_pc; // @[Reg.scala 15:16]
  reg [63:0] _RAND_181;
  reg [1:0] r_btb_updatePipe_bits_cfiType; // @[Reg.scala 15:16]
  reg [31:0] _RAND_182;
  wire [24:0] pageHit_p; // @[BTB.scala 213:39]
  wire  pageHit_lo_lo; // @[BTB.scala 216:29]
  wire  pageHit_lo_hi_lo; // @[BTB.scala 216:29]
  wire  pageHit_lo_hi_hi; // @[BTB.scala 216:29]
  wire  pageHit_hi_lo; // @[BTB.scala 216:29]
  wire  pageHit_hi_hi_lo; // @[BTB.scala 216:29]
  wire  pageHit_hi_hi_hi; // @[BTB.scala 216:29]
  wire [5:0] _pageHit_T; // @[Cat.scala 30:58]
  wire [5:0] pageHit; // @[BTB.scala 216:15]
  wire [12:0] idxHit_idx; // @[BTB.scala 219:19]
  wire  idxHit_lo_lo_lo_lo; // @[BTB.scala 220:16]
  wire  idxHit_lo_lo_lo_hi_lo; // @[BTB.scala 220:16]
  wire  idxHit_lo_lo_lo_hi_hi; // @[BTB.scala 220:16]
  wire  idxHit_lo_lo_hi_lo_lo; // @[BTB.scala 220:16]
  wire  idxHit_lo_lo_hi_lo_hi; // @[BTB.scala 220:16]
  wire  idxHit_lo_lo_hi_hi_lo; // @[BTB.scala 220:16]
  wire  idxHit_lo_lo_hi_hi_hi; // @[BTB.scala 220:16]
  wire  idxHit_lo_hi_lo_lo; // @[BTB.scala 220:16]
  wire  idxHit_lo_hi_lo_hi_lo; // @[BTB.scala 220:16]
  wire  idxHit_lo_hi_lo_hi_hi; // @[BTB.scala 220:16]
  wire  idxHit_lo_hi_hi_lo_lo; // @[BTB.scala 220:16]
  wire  idxHit_lo_hi_hi_lo_hi; // @[BTB.scala 220:16]
  wire  idxHit_lo_hi_hi_hi_lo; // @[BTB.scala 220:16]
  wire  idxHit_lo_hi_hi_hi_hi; // @[BTB.scala 220:16]
  wire  idxHit_hi_lo_lo_lo; // @[BTB.scala 220:16]
  wire  idxHit_hi_lo_lo_hi_lo; // @[BTB.scala 220:16]
  wire  idxHit_hi_lo_lo_hi_hi; // @[BTB.scala 220:16]
  wire  idxHit_hi_lo_hi_lo_lo; // @[BTB.scala 220:16]
  wire  idxHit_hi_lo_hi_lo_hi; // @[BTB.scala 220:16]
  wire  idxHit_hi_lo_hi_hi_lo; // @[BTB.scala 220:16]
  wire  idxHit_hi_lo_hi_hi_hi; // @[BTB.scala 220:16]
  wire  idxHit_hi_hi_lo_lo; // @[BTB.scala 220:16]
  wire  idxHit_hi_hi_lo_hi_lo; // @[BTB.scala 220:16]
  wire  idxHit_hi_hi_lo_hi_hi; // @[BTB.scala 220:16]
  wire  idxHit_hi_hi_hi_lo_lo; // @[BTB.scala 220:16]
  wire  idxHit_hi_hi_hi_lo_hi; // @[BTB.scala 220:16]
  wire  idxHit_hi_hi_hi_hi_lo; // @[BTB.scala 220:16]
  wire  idxHit_hi_hi_hi_hi_hi; // @[BTB.scala 220:16]
  wire [6:0] idxHit_lo_lo; // @[Cat.scala 30:58]
  wire [13:0] idxHit_lo; // @[Cat.scala 30:58]
  wire [6:0] idxHit_hi_lo; // @[Cat.scala 30:58]
  wire [27:0] _idxHit_T; // @[Cat.scala 30:58]
  wire [27:0] idxHit; // @[BTB.scala 220:32]
  wire [24:0] updatePageHit_p; // @[BTB.scala 213:39]
  wire  updatePageHit_lo_lo; // @[BTB.scala 216:29]
  wire  updatePageHit_lo_hi_lo; // @[BTB.scala 216:29]
  wire  updatePageHit_lo_hi_hi; // @[BTB.scala 216:29]
  wire  updatePageHit_hi_lo; // @[BTB.scala 216:29]
  wire  updatePageHit_hi_hi_lo; // @[BTB.scala 216:29]
  wire  updatePageHit_hi_hi_hi; // @[BTB.scala 216:29]
  wire [5:0] _updatePageHit_T; // @[Cat.scala 30:58]
  wire [5:0] updatePageHit; // @[BTB.scala 216:15]
  wire  updateHit; // @[BTB.scala 234:48]
  wire  useUpdatePageHit; // @[BTB.scala 236:40]
  wire  usePageHit; // @[BTB.scala 237:28]
  wire  doIdxPageRepl; // @[BTB.scala 238:23]
  reg [2:0] nextPageRepl; // @[BTB.scala 239:29]
  reg [31:0] _RAND_183;
  wire [4:0] idxPageRepl_hi; // @[BTB.scala 240:32]
  wire  idxPageRepl_lo; // @[BTB.scala 240:53]
  wire [5:0] _idxPageRepl_T; // @[Cat.scala 30:58]
  wire [7:0] _idxPageRepl_T_1; // @[OneHot.scala 58:35]
  wire [7:0] _idxPageRepl_T_2; // @[BTB.scala 240:70]
  wire [7:0] _GEN_430; // @[BTB.scala 240:65]
  wire [7:0] idxPageRepl; // @[BTB.scala 240:65]
  wire [7:0] idxPageUpdateOH; // @[BTB.scala 241:28]
  wire [3:0] idxPageUpdate_hi; // @[OneHot.scala 30:18]
  wire [3:0] idxPageUpdate_lo; // @[OneHot.scala 31:18]
  wire  idxPageUpdate_hi_1; // @[OneHot.scala 32:14]
  wire [3:0] _idxPageUpdate_T; // @[OneHot.scala 32:28]
  wire [1:0] idxPageUpdate_hi_2; // @[OneHot.scala 30:18]
  wire [1:0] idxPageUpdate_lo_1; // @[OneHot.scala 31:18]
  wire  idxPageUpdate_hi_3; // @[OneHot.scala 32:14]
  wire [1:0] _idxPageUpdate_T_1; // @[OneHot.scala 32:28]
  wire  idxPageUpdate_lo_2; // @[CircuitMath.scala 30:8]
  wire [2:0] idxPageUpdate; // @[Cat.scala 30:58]
  wire [7:0] idxPageReplEn; // @[BTB.scala 243:26]
  wire  samePage; // @[BTB.scala 245:45]
  wire  doTgtPageRepl; // @[BTB.scala 246:33]
  wire [4:0] tgtPageRepl_hi; // @[BTB.scala 247:71]
  wire  tgtPageRepl_lo; // @[BTB.scala 247:100]
  wire [5:0] _tgtPageRepl_T; // @[Cat.scala 30:58]
  wire [7:0] tgtPageRepl; // @[BTB.scala 247:24]
  wire [7:0] _tgtPageUpdate_T; // @[BTB.scala 248:45]
  wire [7:0] _GEN_431; // @[BTB.scala 248:40]
  wire [7:0] _tgtPageUpdate_T_1; // @[BTB.scala 248:40]
  wire [3:0] tgtPageUpdate_hi; // @[OneHot.scala 30:18]
  wire [3:0] tgtPageUpdate_lo; // @[OneHot.scala 31:18]
  wire  tgtPageUpdate_hi_1; // @[OneHot.scala 32:14]
  wire [3:0] _tgtPageUpdate_T_2; // @[OneHot.scala 32:28]
  wire [1:0] tgtPageUpdate_hi_2; // @[OneHot.scala 30:18]
  wire [1:0] tgtPageUpdate_lo_1; // @[OneHot.scala 31:18]
  wire  tgtPageUpdate_hi_3; // @[OneHot.scala 32:14]
  wire [1:0] _tgtPageUpdate_T_3; // @[OneHot.scala 32:28]
  wire  tgtPageUpdate_lo_2; // @[CircuitMath.scala 30:8]
  wire [2:0] tgtPageUpdate; // @[Cat.scala 30:58]
  wire [7:0] tgtPageReplEn; // @[BTB.scala 249:26]
  wire  _T; // @[BTB.scala 251:46]
  wire  _T_1; // @[BTB.scala 251:28]
  wire  both; // @[BTB.scala 252:30]
  wire [1:0] _next_T; // @[BTB.scala 253:40]
  wire [2:0] _GEN_432; // @[BTB.scala 253:29]
  wire [2:0] next; // @[BTB.scala 253:29]
  wire  _nextPageRepl_T; // @[BTB.scala 254:30]
  reg [26:0] state_reg; // @[Replacement.scala 168:70]
  reg [31:0] _RAND_184;
  wire  waddr_hi; // @[Replacement.scala 243:38]
  wire [10:0] waddr_left_subtree_state; // @[package.scala 154:13]
  wire [14:0] waddr_right_subtree_state; // @[Replacement.scala 245:38]
  wire  waddr_hi_1; // @[Replacement.scala 243:38]
  wire [2:0] waddr_left_subtree_state_1; // @[package.scala 154:13]
  wire [6:0] waddr_right_subtree_state_1; // @[Replacement.scala 245:38]
  wire  waddr_hi_2; // @[Replacement.scala 243:38]
  wire  waddr_left_subtree_state_2; // @[package.scala 154:13]
  wire  waddr_right_subtree_state_2; // @[Replacement.scala 245:38]
  wire  waddr_lo; // @[Replacement.scala 250:16]
  wire [1:0] _waddr_T_2; // @[Cat.scala 30:58]
  wire  waddr_hi_3; // @[Replacement.scala 243:38]
  wire [2:0] waddr_left_subtree_state_3; // @[package.scala 154:13]
  wire [2:0] waddr_right_subtree_state_3; // @[Replacement.scala 245:38]
  wire  waddr_hi_4; // @[Replacement.scala 243:38]
  wire  waddr_left_subtree_state_4; // @[package.scala 154:13]
  wire  waddr_right_subtree_state_4; // @[Replacement.scala 245:38]
  wire  waddr_lo_1; // @[Replacement.scala 250:16]
  wire [1:0] _waddr_T_5; // @[Cat.scala 30:58]
  wire  waddr_hi_5; // @[Replacement.scala 243:38]
  wire  waddr_left_subtree_state_5; // @[package.scala 154:13]
  wire  waddr_right_subtree_state_5; // @[Replacement.scala 245:38]
  wire  waddr_lo_2; // @[Replacement.scala 250:16]
  wire [1:0] _waddr_T_8; // @[Cat.scala 30:58]
  wire [1:0] waddr_lo_3; // @[Replacement.scala 250:16]
  wire [2:0] _waddr_T_9; // @[Cat.scala 30:58]
  wire [2:0] waddr_lo_4; // @[Replacement.scala 250:16]
  wire [3:0] _waddr_T_10; // @[Cat.scala 30:58]
  wire  waddr_hi_6; // @[Replacement.scala 243:38]
  wire [6:0] waddr_left_subtree_state_6; // @[package.scala 154:13]
  wire [6:0] waddr_right_subtree_state_6; // @[Replacement.scala 245:38]
  wire  waddr_hi_7; // @[Replacement.scala 243:38]
  wire [2:0] waddr_left_subtree_state_7; // @[package.scala 154:13]
  wire [2:0] waddr_right_subtree_state_7; // @[Replacement.scala 245:38]
  wire  waddr_hi_8; // @[Replacement.scala 243:38]
  wire  waddr_left_subtree_state_8; // @[package.scala 154:13]
  wire  waddr_right_subtree_state_8; // @[Replacement.scala 245:38]
  wire  waddr_lo_5; // @[Replacement.scala 250:16]
  wire [1:0] _waddr_T_13; // @[Cat.scala 30:58]
  wire  waddr_hi_9; // @[Replacement.scala 243:38]
  wire  waddr_left_subtree_state_9; // @[package.scala 154:13]
  wire  waddr_right_subtree_state_9; // @[Replacement.scala 245:38]
  wire  waddr_lo_6; // @[Replacement.scala 250:16]
  wire [1:0] _waddr_T_16; // @[Cat.scala 30:58]
  wire [1:0] waddr_lo_7; // @[Replacement.scala 250:16]
  wire [2:0] _waddr_T_17; // @[Cat.scala 30:58]
  wire  waddr_hi_10; // @[Replacement.scala 243:38]
  wire [2:0] waddr_left_subtree_state_10; // @[package.scala 154:13]
  wire [2:0] waddr_right_subtree_state_10; // @[Replacement.scala 245:38]
  wire  waddr_hi_11; // @[Replacement.scala 243:38]
  wire  waddr_left_subtree_state_11; // @[package.scala 154:13]
  wire  waddr_right_subtree_state_11; // @[Replacement.scala 245:38]
  wire  waddr_lo_8; // @[Replacement.scala 250:16]
  wire [1:0] _waddr_T_20; // @[Cat.scala 30:58]
  wire  waddr_hi_12; // @[Replacement.scala 243:38]
  wire  waddr_left_subtree_state_12; // @[package.scala 154:13]
  wire  waddr_right_subtree_state_12; // @[Replacement.scala 245:38]
  wire  waddr_lo_9; // @[Replacement.scala 250:16]
  wire [1:0] _waddr_T_23; // @[Cat.scala 30:58]
  wire [1:0] waddr_lo_10; // @[Replacement.scala 250:16]
  wire [2:0] _waddr_T_24; // @[Cat.scala 30:58]
  wire [2:0] waddr_lo_11; // @[Replacement.scala 250:16]
  wire [3:0] _waddr_T_25; // @[Cat.scala 30:58]
  wire [3:0] waddr_lo_12; // @[Replacement.scala 250:16]
  wire [4:0] _waddr_T_26; // @[Cat.scala 30:58]
  wire [4:0] waddr; // @[BTB.scala 258:18]
  reg  r_respPipe_valid; // @[Valid.scala 117:22]
  reg [31:0] _RAND_185;
  reg  r_respPipe_bits_taken; // @[Reg.scala 15:16]
  reg [31:0] _RAND_186;
  reg [4:0] r_respPipe_bits_entry; // @[Reg.scala 15:16]
  reg [31:0] _RAND_187;
  wire  _T_2; // @[BTB.scala 260:22]
  wire  _T_3; // @[BTB.scala 260:43]
  wire [4:0] state_reg_touch_way_sized; // @[BTB.scala 261:20]
  wire  state_reg_hi_hi; // @[Replacement.scala 196:33]
  wire  state_reg_hi_hi_1; // @[Replacement.scala 196:33]
  wire  state_reg_hi_hi_2; // @[Replacement.scala 196:33]
  wire  state_reg_hi_lo; // @[Replacement.scala 203:16]
  wire  state_reg_lo; // @[Replacement.scala 206:16]
  wire [2:0] _state_reg_T_8; // @[Cat.scala 30:58]
  wire [2:0] state_reg_hi_lo_1; // @[Replacement.scala 203:16]
  wire  state_reg_hi_hi_3; // @[Replacement.scala 196:33]
  wire  state_reg_hi_hi_4; // @[Replacement.scala 196:33]
  wire  state_reg_hi_lo_2; // @[Replacement.scala 203:16]
  wire  state_reg_lo_1; // @[Replacement.scala 206:16]
  wire [2:0] _state_reg_T_17; // @[Cat.scala 30:58]
  wire [2:0] state_reg_hi_lo_3; // @[Replacement.scala 203:16]
  wire  state_reg_hi_lo_4; // @[Replacement.scala 203:16]
  wire  state_reg_lo_2; // @[Replacement.scala 206:16]
  wire [2:0] _state_reg_T_25; // @[Cat.scala 30:58]
  wire [2:0] state_reg_lo_3; // @[Replacement.scala 206:16]
  wire [6:0] _state_reg_T_26; // @[Cat.scala 30:58]
  wire [6:0] state_reg_lo_4; // @[Replacement.scala 206:16]
  wire [10:0] _state_reg_T_27; // @[Cat.scala 30:58]
  wire [10:0] state_reg_hi_lo_5; // @[Replacement.scala 203:16]
  wire  state_reg_hi_lo_6; // @[Replacement.scala 203:16]
  wire  state_reg_lo_5; // @[Replacement.scala 206:16]
  wire [2:0] _state_reg_T_37; // @[Cat.scala 30:58]
  wire [2:0] state_reg_hi_lo_7; // @[Replacement.scala 203:16]
  wire  state_reg_hi_lo_8; // @[Replacement.scala 203:16]
  wire  state_reg_lo_6; // @[Replacement.scala 206:16]
  wire [2:0] _state_reg_T_45; // @[Cat.scala 30:58]
  wire [2:0] state_reg_lo_7; // @[Replacement.scala 206:16]
  wire [6:0] _state_reg_T_46; // @[Cat.scala 30:58]
  wire [6:0] state_reg_hi_lo_9; // @[Replacement.scala 203:16]
  wire  state_reg_hi_lo_10; // @[Replacement.scala 203:16]
  wire  state_reg_lo_8; // @[Replacement.scala 206:16]
  wire [2:0] _state_reg_T_55; // @[Cat.scala 30:58]
  wire [2:0] state_reg_hi_lo_11; // @[Replacement.scala 203:16]
  wire  state_reg_hi_lo_12; // @[Replacement.scala 203:16]
  wire  state_reg_lo_9; // @[Replacement.scala 206:16]
  wire [2:0] _state_reg_T_63; // @[Cat.scala 30:58]
  wire [2:0] state_reg_lo_10; // @[Replacement.scala 206:16]
  wire [6:0] _state_reg_T_64; // @[Cat.scala 30:58]
  wire [6:0] state_reg_lo_11; // @[Replacement.scala 206:16]
  wire [14:0] _state_reg_T_65; // @[Cat.scala 30:58]
  wire [14:0] state_reg_lo_12; // @[Replacement.scala 206:16]
  wire [26:0] _state_reg_T_66; // @[Cat.scala 30:58]
  wire [31:0] mask; // @[OneHot.scala 58:35]
  wire [3:0] _idxPages_T; // @[BTB.scala 268:38]
  wire [31:0] _GEN_433; // @[BTB.scala 271:55]
  wire [31:0] _isValid_T; // @[BTB.scala 271:55]
  wire [31:0] _isValid_T_2; // @[BTB.scala 271:71]
  wire [31:0] _isValid_T_3; // @[BTB.scala 271:19]
  wire  idxWritesEven; // @[BTB.scala 276:25]
  wire [7:0] _T_5; // @[BTB.scala 282:24]
  wire [7:0] _T_12; // @[BTB.scala 284:24]
  wire [7:0] _GEN_435; // @[BTB.scala 286:28]
  wire [7:0] _pageValid_T; // @[BTB.scala 286:28]
  wire [7:0] _pageValid_T_1; // @[BTB.scala 286:44]
  wire [31:0] _GEN_338; // @[BTB.scala 264:29]
  wire [7:0] _GEN_373; // @[BTB.scala 264:29]
  wire [6:0] _io_resp_valid_T; // @[BTB.scala 289:29]
  wire [2:0] _io_resp_valid_T_29; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_30; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_31; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_32; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_33; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_34; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_35; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_36; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_37; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_38; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_39; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_40; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_41; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_42; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_43; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_44; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_45; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_46; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_47; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_48; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_49; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_50; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_51; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_52; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_53; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_54; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_55; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_56; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_57; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_58; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_59; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_60; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_61; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_62; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_63; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_64; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_65; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_66; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_67; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_68; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_69; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_70; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_71; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_72; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_73; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_74; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_75; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_76; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_77; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_78; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_79; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_80; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_81; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_82; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_valid_T_83; // @[Mux.scala 27:72]
  wire [6:0] _io_resp_valid_T_84; // @[BTB.scala 289:34]
  wire [2:0] _io_resp_bits_target_T_28; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_29; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_30; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_31; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_32; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_33; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_34; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_35; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_36; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_37; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_38; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_39; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_40; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_41; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_42; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_43; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_44; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_45; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_46; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_47; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_48; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_49; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_50; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_51; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_52; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_53; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_54; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_55; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_56; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_57; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_58; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_59; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_60; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_61; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_62; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_63; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_64; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_65; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_66; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_67; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_68; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_69; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_70; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_71; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_72; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_73; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_74; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_75; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_76; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_77; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_78; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_79; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_80; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_81; // @[Mux.scala 27:72]
  wire [2:0] _io_resp_bits_target_T_82; // @[Mux.scala 27:72]
  wire  _io_resp_bits_target_T_83; // @[package.scala 32:86]
  wire [24:0] _io_resp_bits_target_T_84; // @[package.scala 32:76]
  wire  _io_resp_bits_target_T_85; // @[package.scala 32:86]
  wire [24:0] _io_resp_bits_target_T_86; // @[package.scala 32:76]
  wire  _io_resp_bits_target_T_87; // @[package.scala 32:86]
  wire [24:0] _io_resp_bits_target_T_88; // @[package.scala 32:76]
  wire  _io_resp_bits_target_T_89; // @[package.scala 32:86]
  wire [24:0] _io_resp_bits_target_T_90; // @[package.scala 32:76]
  wire  _io_resp_bits_target_T_91; // @[package.scala 32:86]
  wire [24:0] _io_resp_bits_target_T_92; // @[package.scala 32:76]
  wire  _io_resp_bits_target_T_93; // @[package.scala 32:86]
  wire [24:0] _io_resp_bits_target_T_94; // @[package.scala 32:76]
  wire  _io_resp_bits_target_T_95; // @[package.scala 32:86]
  wire [24:0] io_resp_bits_target_hi; // @[package.scala 32:76]
  wire [12:0] _io_resp_bits_target_T_124; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_125; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_126; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_127; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_128; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_129; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_130; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_131; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_132; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_133; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_134; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_135; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_136; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_137; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_138; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_139; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_140; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_141; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_142; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_143; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_144; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_145; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_146; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_147; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_148; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_149; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_150; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_151; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_152; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_153; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_154; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_155; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_156; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_157; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_158; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_159; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_160; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_161; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_162; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_163; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_164; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_165; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_166; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_167; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_168; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_169; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_170; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_171; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_172; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_173; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_174; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_175; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_176; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_177; // @[Mux.scala 27:72]
  wire [12:0] _io_resp_bits_target_T_178; // @[Mux.scala 27:72]
  wire [13:0] io_resp_bits_target_lo; // @[BTB.scala 291:88]
  wire [38:0] _io_resp_bits_target_T_179; // @[Cat.scala 30:58]
  wire [11:0] io_resp_bits_entry_hi; // @[OneHot.scala 30:18]
  wire [15:0] io_resp_bits_entry_lo; // @[OneHot.scala 31:18]
  wire  io_resp_bits_entry_hi_1; // @[OneHot.scala 32:14]
  wire [15:0] _GEN_436; // @[OneHot.scala 32:28]
  wire [15:0] _io_resp_bits_entry_T; // @[OneHot.scala 32:28]
  wire [7:0] io_resp_bits_entry_hi_2; // @[OneHot.scala 30:18]
  wire [7:0] io_resp_bits_entry_lo_1; // @[OneHot.scala 31:18]
  wire  io_resp_bits_entry_hi_3; // @[OneHot.scala 32:14]
  wire [7:0] _io_resp_bits_entry_T_1; // @[OneHot.scala 32:28]
  wire [3:0] io_resp_bits_entry_hi_4; // @[OneHot.scala 30:18]
  wire [3:0] io_resp_bits_entry_lo_2; // @[OneHot.scala 31:18]
  wire  io_resp_bits_entry_hi_5; // @[OneHot.scala 32:14]
  wire [3:0] _io_resp_bits_entry_T_2; // @[OneHot.scala 32:28]
  wire [1:0] io_resp_bits_entry_hi_6; // @[OneHot.scala 30:18]
  wire [1:0] io_resp_bits_entry_lo_3; // @[OneHot.scala 31:18]
  wire  io_resp_bits_entry_hi_7; // @[OneHot.scala 32:14]
  wire [1:0] _io_resp_bits_entry_T_3; // @[OneHot.scala 32:28]
  wire  io_resp_bits_entry_lo_4; // @[CircuitMath.scala 30:8]
  wire [3:0] io_resp_bits_entry_lo_7; // @[Cat.scala 30:58]
  wire  _io_resp_bits_bridx_T_28; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_29; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_30; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_31; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_32; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_33; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_34; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_35; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_36; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_37; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_38; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_39; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_40; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_41; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_42; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_43; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_44; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_45; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_46; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_47; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_48; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_49; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_50; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_51; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_52; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_53; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_54; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_55; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_56; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_57; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_58; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_59; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_60; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_61; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_62; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_63; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_64; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_65; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_66; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_67; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_68; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_69; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_70; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_71; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_72; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_73; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_74; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_75; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_76; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_77; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_78; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_79; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_80; // @[Mux.scala 27:72]
  wire  _io_resp_bits_bridx_T_81; // @[Mux.scala 27:72]
  wire  leftOne; // @[Misc.scala 180:37]
  wire  leftOne_1; // @[Misc.scala 180:37]
  wire  rightOne; // @[Misc.scala 181:39]
  wire  rightOne_1; // @[Misc.scala 182:16]
  wire  rightTwo; // @[Misc.scala 182:61]
  wire  leftOne_2; // @[Misc.scala 182:16]
  wire  _T_29; // @[Misc.scala 182:61]
  wire  leftTwo; // @[Misc.scala 182:49]
  wire  leftOne_3; // @[Misc.scala 180:37]
  wire  rightOne_2; // @[Misc.scala 181:39]
  wire  leftOne_4; // @[Misc.scala 182:16]
  wire  leftTwo_1; // @[Misc.scala 182:61]
  wire  leftOne_5; // @[Misc.scala 180:37]
  wire  rightOne_3; // @[Misc.scala 181:39]
  wire  rightOne_4; // @[Misc.scala 182:16]
  wire  rightTwo_1; // @[Misc.scala 182:61]
  wire  rightOne_5; // @[Misc.scala 182:16]
  wire  _T_41; // @[Misc.scala 182:37]
  wire  _T_42; // @[Misc.scala 182:61]
  wire  rightTwo_2; // @[Misc.scala 182:49]
  wire  leftOne_6; // @[Misc.scala 182:16]
  wire  _T_43; // @[Misc.scala 182:37]
  wire  _T_44; // @[Misc.scala 182:61]
  wire  leftTwo_2; // @[Misc.scala 182:49]
  wire  leftOne_7; // @[Misc.scala 180:37]
  wire  leftOne_8; // @[Misc.scala 180:37]
  wire  rightOne_6; // @[Misc.scala 181:39]
  wire  rightOne_7; // @[Misc.scala 182:16]
  wire  rightTwo_3; // @[Misc.scala 182:61]
  wire  leftOne_9; // @[Misc.scala 182:16]
  wire  _T_54; // @[Misc.scala 182:61]
  wire  leftTwo_3; // @[Misc.scala 182:49]
  wire  leftOne_10; // @[Misc.scala 180:37]
  wire  rightOne_8; // @[Misc.scala 181:39]
  wire  leftOne_11; // @[Misc.scala 182:16]
  wire  leftTwo_4; // @[Misc.scala 182:61]
  wire  leftOne_12; // @[Misc.scala 180:37]
  wire  rightOne_9; // @[Misc.scala 181:39]
  wire  rightOne_10; // @[Misc.scala 182:16]
  wire  rightTwo_4; // @[Misc.scala 182:61]
  wire  rightOne_11; // @[Misc.scala 182:16]
  wire  _T_66; // @[Misc.scala 182:37]
  wire  _T_67; // @[Misc.scala 182:61]
  wire  rightTwo_5; // @[Misc.scala 182:49]
  wire  rightOne_12; // @[Misc.scala 182:16]
  wire  _T_68; // @[Misc.scala 182:37]
  wire  _T_69; // @[Misc.scala 182:61]
  wire  rightTwo_6; // @[Misc.scala 182:49]
  wire  leftOne_13; // @[Misc.scala 182:16]
  wire  _T_70; // @[Misc.scala 182:37]
  wire  _T_71; // @[Misc.scala 182:61]
  wire  leftTwo_5; // @[Misc.scala 182:49]
  wire  leftOne_14; // @[Misc.scala 180:37]
  wire  leftOne_15; // @[Misc.scala 180:37]
  wire  rightOne_13; // @[Misc.scala 181:39]
  wire  rightOne_14; // @[Misc.scala 182:16]
  wire  rightTwo_7; // @[Misc.scala 182:61]
  wire  leftOne_16; // @[Misc.scala 182:16]
  wire  _T_82; // @[Misc.scala 182:61]
  wire  leftTwo_6; // @[Misc.scala 182:49]
  wire  leftOne_17; // @[Misc.scala 180:37]
  wire  rightOne_15; // @[Misc.scala 181:39]
  wire  leftOne_18; // @[Misc.scala 182:16]
  wire  leftTwo_7; // @[Misc.scala 182:61]
  wire  leftOne_19; // @[Misc.scala 180:37]
  wire  rightOne_16; // @[Misc.scala 181:39]
  wire  rightOne_17; // @[Misc.scala 182:16]
  wire  rightTwo_8; // @[Misc.scala 182:61]
  wire  rightOne_18; // @[Misc.scala 182:16]
  wire  _T_94; // @[Misc.scala 182:37]
  wire  _T_95; // @[Misc.scala 182:61]
  wire  rightTwo_9; // @[Misc.scala 182:49]
  wire  leftOne_20; // @[Misc.scala 182:16]
  wire  _T_96; // @[Misc.scala 182:37]
  wire  _T_97; // @[Misc.scala 182:61]
  wire  leftTwo_8; // @[Misc.scala 182:49]
  wire  leftOne_21; // @[Misc.scala 180:37]
  wire  leftOne_22; // @[Misc.scala 180:37]
  wire  rightOne_19; // @[Misc.scala 181:39]
  wire  rightOne_20; // @[Misc.scala 182:16]
  wire  rightTwo_10; // @[Misc.scala 182:61]
  wire  leftOne_23; // @[Misc.scala 182:16]
  wire  _T_107; // @[Misc.scala 182:61]
  wire  leftTwo_9; // @[Misc.scala 182:49]
  wire  leftOne_24; // @[Misc.scala 180:37]
  wire  rightOne_21; // @[Misc.scala 181:39]
  wire  leftOne_25; // @[Misc.scala 182:16]
  wire  leftTwo_10; // @[Misc.scala 182:61]
  wire  leftOne_26; // @[Misc.scala 180:37]
  wire  rightOne_22; // @[Misc.scala 181:39]
  wire  rightOne_23; // @[Misc.scala 182:16]
  wire  rightTwo_11; // @[Misc.scala 182:61]
  wire  rightOne_24; // @[Misc.scala 182:16]
  wire  _T_119; // @[Misc.scala 182:37]
  wire  _T_120; // @[Misc.scala 182:61]
  wire  rightTwo_12; // @[Misc.scala 182:49]
  wire  rightOne_25; // @[Misc.scala 182:16]
  wire  _T_121; // @[Misc.scala 182:37]
  wire  _T_122; // @[Misc.scala 182:61]
  wire  rightTwo_13; // @[Misc.scala 182:49]
  wire  rightOne_26; // @[Misc.scala 182:16]
  wire  _T_123; // @[Misc.scala 182:37]
  wire  _T_124; // @[Misc.scala 182:61]
  wire  rightTwo_14; // @[Misc.scala 182:49]
  wire  _T_126; // @[Misc.scala 182:37]
  wire  _T_127; // @[Misc.scala 182:61]
  wire  _T_128; // @[Misc.scala 182:49]
  wire [27:0] _isValid_T_5; // @[BTB.scala 299:24]
  wire [31:0] _GEN_374; // @[BTB.scala 298:37]
  wire [31:0] _GEN_375; // @[BTB.scala 301:19]
  reg [7:0] history; // @[BTB.scala 119:24]
  reg [31:0] _RAND_188;
  reg [9:0] reset_waddr; // @[BTB.scala 121:36]
  reg [31:0] _RAND_189;
  wire  resetting; // @[BTB.scala 122:27]
  wire [9:0] _reset_waddr_T_1; // @[BTB.scala 126:49]
  wire [36:0] waddr_hi_13; // @[BTB.scala 87:21]
  wire [8:0] _GEN_437; // @[BTB.scala 88:42]
  wire [8:0] _waddr_T_30; // @[BTB.scala 88:42]
  wire [15:0] _waddr_T_31; // @[BTB.scala 84:12]
  wire [8:0] _waddr_T_33; // @[BTB.scala 90:44]
  wire [8:0] _waddr_T_34; // @[BTB.scala 90:20]
  wire [9:0] _GEN_383; // @[BTB.scala 100:23]
  wire [9:0] _GEN_388; // @[BTB.scala 313:40]
  wire [9:0] waddr_1; // @[BTB.scala 312:32]
  wire  _GEN_387; // @[BTB.scala 313:40]
  wire  _GEN_384; // @[BTB.scala 100:23]
  wire  _GEN_389; // @[BTB.scala 313:40]
  wire  isBranch_lo_lo_lo_lo; // @[BTB.scala 307:44]
  wire  isBranch_lo_lo_lo_hi_lo; // @[BTB.scala 307:44]
  wire  isBranch_lo_lo_lo_hi_hi; // @[BTB.scala 307:44]
  wire  isBranch_lo_lo_hi_lo_lo; // @[BTB.scala 307:44]
  wire  isBranch_lo_lo_hi_lo_hi; // @[BTB.scala 307:44]
  wire  isBranch_lo_lo_hi_hi_lo; // @[BTB.scala 307:44]
  wire  isBranch_lo_lo_hi_hi_hi; // @[BTB.scala 307:44]
  wire  isBranch_lo_hi_lo_lo; // @[BTB.scala 307:44]
  wire  isBranch_lo_hi_lo_hi_lo; // @[BTB.scala 307:44]
  wire  isBranch_lo_hi_lo_hi_hi; // @[BTB.scala 307:44]
  wire  isBranch_lo_hi_hi_lo_lo; // @[BTB.scala 307:44]
  wire  isBranch_lo_hi_hi_lo_hi; // @[BTB.scala 307:44]
  wire  isBranch_lo_hi_hi_hi_lo; // @[BTB.scala 307:44]
  wire  isBranch_lo_hi_hi_hi_hi; // @[BTB.scala 307:44]
  wire  isBranch_hi_lo_lo_lo; // @[BTB.scala 307:44]
  wire  isBranch_hi_lo_lo_hi_lo; // @[BTB.scala 307:44]
  wire  isBranch_hi_lo_lo_hi_hi; // @[BTB.scala 307:44]
  wire  isBranch_hi_lo_hi_lo_lo; // @[BTB.scala 307:44]
  wire  isBranch_hi_lo_hi_lo_hi; // @[BTB.scala 307:44]
  wire  isBranch_hi_lo_hi_hi_lo; // @[BTB.scala 307:44]
  wire  isBranch_hi_lo_hi_hi_hi; // @[BTB.scala 307:44]
  wire  isBranch_hi_hi_lo_lo; // @[BTB.scala 307:44]
  wire  isBranch_hi_hi_lo_hi_lo; // @[BTB.scala 307:44]
  wire  isBranch_hi_hi_lo_hi_hi; // @[BTB.scala 307:44]
  wire  isBranch_hi_hi_hi_lo_lo; // @[BTB.scala 307:44]
  wire  isBranch_hi_hi_hi_lo_hi; // @[BTB.scala 307:44]
  wire  isBranch_hi_hi_hi_hi_lo; // @[BTB.scala 307:44]
  wire  isBranch_hi_hi_hi_hi_hi; // @[BTB.scala 307:44]
  wire [6:0] isBranch_lo_lo; // @[Cat.scala 30:58]
  wire [13:0] isBranch_lo; // @[Cat.scala 30:58]
  wire [6:0] isBranch_hi_lo; // @[Cat.scala 30:58]
  wire [27:0] _isBranch_T; // @[Cat.scala 30:58]
  wire [27:0] _isBranch_T_1; // @[BTB.scala 307:28]
  wire  isBranch; // @[BTB.scala 307:72]
  wire [36:0] res_res_value_hi; // @[BTB.scala 87:21]
  wire [8:0] _GEN_438; // @[BTB.scala 88:42]
  wire [8:0] _res_res_value_T_3; // @[BTB.scala 88:42]
  wire [15:0] _res_res_value_T_4; // @[BTB.scala 84:12]
  wire [8:0] _res_res_value_T_6; // @[BTB.scala 90:44]
  wire  res_value; // @[BTB.scala 94:21]
  wire [6:0] history_lo; // @[BTB.scala 115:35]
  wire [7:0] _history_T; // @[Cat.scala 30:58]
  wire [6:0] history_lo_1; // @[BTB.scala 112:37]
  wire [7:0] _history_T_1; // @[Cat.scala 30:58]
  wire  _T_134; // @[BTB.scala 322:22]
  reg [2:0] count; // @[BTB.scala 58:30]
  reg [31:0] _RAND_190;
  reg [2:0] pos; // @[BTB.scala 59:28]
  reg [31:0] _RAND_191;
  reg [38:0] stack_0; // @[BTB.scala 60:26]
  reg [63:0] _RAND_192;
  reg [38:0] stack_1; // @[BTB.scala 60:26]
  reg [63:0] _RAND_193;
  reg [38:0] stack_2; // @[BTB.scala 60:26]
  reg [63:0] _RAND_194;
  reg [38:0] stack_3; // @[BTB.scala 60:26]
  reg [63:0] _RAND_195;
  reg [38:0] stack_4; // @[BTB.scala 60:26]
  reg [63:0] _RAND_196;
  reg [38:0] stack_5; // @[BTB.scala 60:26]
  reg [63:0] _RAND_197;
  wire  doPeek_lo_lo_lo_lo; // @[BTB.scala 328:42]
  wire  doPeek_lo_lo_lo_hi_lo; // @[BTB.scala 328:42]
  wire  doPeek_lo_lo_lo_hi_hi; // @[BTB.scala 328:42]
  wire  doPeek_lo_lo_hi_lo_lo; // @[BTB.scala 328:42]
  wire  doPeek_lo_lo_hi_lo_hi; // @[BTB.scala 328:42]
  wire  doPeek_lo_lo_hi_hi_lo; // @[BTB.scala 328:42]
  wire  doPeek_lo_lo_hi_hi_hi; // @[BTB.scala 328:42]
  wire  doPeek_lo_hi_lo_lo; // @[BTB.scala 328:42]
  wire  doPeek_lo_hi_lo_hi_lo; // @[BTB.scala 328:42]
  wire  doPeek_lo_hi_lo_hi_hi; // @[BTB.scala 328:42]
  wire  doPeek_lo_hi_hi_lo_lo; // @[BTB.scala 328:42]
  wire  doPeek_lo_hi_hi_lo_hi; // @[BTB.scala 328:42]
  wire  doPeek_lo_hi_hi_hi_lo; // @[BTB.scala 328:42]
  wire  doPeek_lo_hi_hi_hi_hi; // @[BTB.scala 328:42]
  wire  doPeek_hi_lo_lo_lo; // @[BTB.scala 328:42]
  wire  doPeek_hi_lo_lo_hi_lo; // @[BTB.scala 328:42]
  wire  doPeek_hi_lo_lo_hi_hi; // @[BTB.scala 328:42]
  wire  doPeek_hi_lo_hi_lo_lo; // @[BTB.scala 328:42]
  wire  doPeek_hi_lo_hi_lo_hi; // @[BTB.scala 328:42]
  wire  doPeek_hi_lo_hi_hi_lo; // @[BTB.scala 328:42]
  wire  doPeek_hi_lo_hi_hi_hi; // @[BTB.scala 328:42]
  wire  doPeek_hi_hi_lo_lo; // @[BTB.scala 328:42]
  wire  doPeek_hi_hi_lo_hi_lo; // @[BTB.scala 328:42]
  wire  doPeek_hi_hi_lo_hi_hi; // @[BTB.scala 328:42]
  wire  doPeek_hi_hi_hi_lo_lo; // @[BTB.scala 328:42]
  wire  doPeek_hi_hi_hi_lo_hi; // @[BTB.scala 328:42]
  wire  doPeek_hi_hi_hi_hi_lo; // @[BTB.scala 328:42]
  wire  doPeek_hi_hi_hi_hi_hi; // @[BTB.scala 328:42]
  wire [6:0] doPeek_lo_lo; // @[Cat.scala 30:58]
  wire [13:0] doPeek_lo; // @[Cat.scala 30:58]
  wire [6:0] doPeek_hi_lo; // @[Cat.scala 30:58]
  wire [27:0] _doPeek_T; // @[Cat.scala 30:58]
  wire [27:0] _doPeek_T_1; // @[BTB.scala 328:26]
  wire  doPeek; // @[BTB.scala 328:67]
  wire  _io_ras_head_valid_T; // @[BTB.scala 56:29]
  wire [38:0] _GEN_397; // @[BTB.scala 330:22]
  wire [38:0] _GEN_398; // @[BTB.scala 330:22]
  wire [38:0] _GEN_399; // @[BTB.scala 330:22]
  wire [38:0] _GEN_400; // @[BTB.scala 330:22]
  wire [38:0] _GEN_401; // @[BTB.scala 330:22]
  wire  _T_137; // @[BTB.scala 331:24]
  wire  _T_138; // @[BTB.scala 335:40]
  wire  _T_139; // @[BTB.scala 45:17]
  wire [2:0] _count_T_1; // @[BTB.scala 45:42]
  wire  _nextPos_T; // @[BTB.scala 46:49]
  wire [2:0] _nextPos_T_3; // @[BTB.scala 46:62]
  wire [2:0] nextPos; // @[BTB.scala 46:22]
  wire  _T_140; // @[BTB.scala 337:46]
  wire [2:0] _count_T_3; // @[BTB.scala 52:20]
  wire  _pos_T; // @[BTB.scala 53:42]
  wire [2:0] _pos_T_3; // @[BTB.scala 53:50]
  reg [19:0] BTB_state; // @[Register tracking BTB state]
  reg [31:0] _RAND_198;
  reg  BTB_cov [0:1048575]; // @[Coverage map for BTB]
  reg [31:0] _RAND_199;
  wire  BTB_cov_read_data; // @[Coverage map for BTB]
  wire [19:0] BTB_cov_read_addr; // @[Coverage map for BTB]
  wire  BTB_cov_write_data; // @[Coverage map for BTB]
  wire [19:0] BTB_cov_write_addr; // @[Coverage map for BTB]
  wire  BTB_cov_write_mask; // @[Coverage map for BTB]
  wire  BTB_cov_write_en; // @[Coverage map for BTB]
  reg [29:0] BTB_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_200;
  wire  mux_cond_0;
  wire  mux_cond_1;
  wire  mux_cond_2;
  wire  mux_cond_3;
  wire  mux_cond_4;
  wire  mux_cond_5;
  wire  mux_cond_6;
  wire  mux_cond_7;
  wire  mux_cond_8;
  wire  mux_cond_9;
  wire  mux_cond_10;
  wire  mux_cond_11;
  wire  mux_cond_12;
  wire  mux_cond_13;
  wire  mux_cond_14;
  wire  mux_cond_15;
  wire  mux_cond_16;
  wire  mux_cond_17;
  wire  mux_cond_18;
  wire  mux_cond_19;
  wire  mux_cond_20;
  wire  mux_cond_21;
  wire  mux_cond_22;
  wire  mux_cond_23;
  wire  mux_cond_24;
  wire  mux_cond_25;
  wire  mux_cond_26;
  wire  mux_cond_27;
  wire  mux_cond_28;
  wire [9:0] nextPageRepl_shl;
  wire [19:0] nextPageRepl_pad;
  wire [3:0] r_respPipe_bits_taken_shl;
  wire [19:0] r_respPipe_bits_taken_pad;
  wire [16:0] r_btb_updatePipe_valid_shl;
  wire [19:0] r_btb_updatePipe_valid_pad;
  wire [14:0] count_shl;
  wire [19:0] count_pad;
  wire [13:0] r_respPipe_valid_shl;
  wire [19:0] r_respPipe_valid_pad;
  wire [3:0] pos_shl;
  wire [19:0] pos_pad;
  wire [13:0] pageValid_shl;
  wire [19:0] pageValid_pad;
  wire [17:0] r_btb_updatePipe_bits_isValid_shl;
  wire [19:0] r_btb_updatePipe_bits_isValid_pad;
  wire [14:0] mux_cond_0_shl;
  wire [19:0] mux_cond_0_pad;
  wire [17:0] mux_cond_1_shl;
  wire [19:0] mux_cond_1_pad;
  wire [3:0] mux_cond_2_shl;
  wire [19:0] mux_cond_2_pad;
  wire [17:0] mux_cond_3_shl;
  wire [19:0] mux_cond_3_pad;
  wire [13:0] mux_cond_4_shl;
  wire [19:0] mux_cond_4_pad;
  wire [3:0] mux_cond_5_shl;
  wire [19:0] mux_cond_5_pad;
  wire [1:0] mux_cond_6_shl;
  wire [19:0] mux_cond_6_pad;
  wire [13:0] mux_cond_7_shl;
  wire [19:0] mux_cond_7_pad;
  wire [16:0] mux_cond_8_shl;
  wire [19:0] mux_cond_8_pad;
  wire [3:0] mux_cond_9_shl;
  wire [19:0] mux_cond_9_pad;
  wire [9:0] mux_cond_10_shl;
  wire [19:0] mux_cond_10_pad;
  wire [3:0] mux_cond_11_shl;
  wire [19:0] mux_cond_11_pad;
  wire [17:0] mux_cond_12_shl;
  wire [19:0] mux_cond_12_pad;
  wire [8:0] mux_cond_13_shl;
  wire [19:0] mux_cond_13_pad;
  wire [4:0] mux_cond_14_shl;
  wire [19:0] mux_cond_14_pad;
  wire [11:0] mux_cond_15_shl;
  wire [19:0] mux_cond_15_pad;
  wire [12:0] mux_cond_16_shl;
  wire [19:0] mux_cond_16_pad;
  wire [5:0] mux_cond_17_shl;
  wire [19:0] mux_cond_17_pad;
  wire  mux_cond_18_shl;
  wire [19:0] mux_cond_18_pad;
  wire [1:0] mux_cond_19_shl;
  wire [19:0] mux_cond_19_pad;
  wire [2:0] mux_cond_20_shl;
  wire [19:0] mux_cond_20_pad;
  wire [5:0] mux_cond_21_shl;
  wire [19:0] mux_cond_21_pad;
  wire [16:0] mux_cond_22_shl;
  wire [19:0] mux_cond_22_pad;
  wire [13:0] mux_cond_23_shl;
  wire [19:0] mux_cond_23_pad;
  wire [19:0] mux_cond_24_shl;
  wire [19:0] mux_cond_24_pad;
  wire [14:0] mux_cond_25_shl;
  wire [19:0] mux_cond_25_pad;
  wire [8:0] mux_cond_26_shl;
  wire [19:0] mux_cond_26_pad;
  wire [18:0] mux_cond_27_shl;
  wire [19:0] mux_cond_27_pad;
  wire [5:0] mux_cond_28_shl;
  wire [19:0] mux_cond_28_pad;
  wire [12:0] cfiType_17_shl;
  wire [19:0] cfiType_17_pad;
  wire [12:0] cfiType_22_shl;
  wire [19:0] cfiType_22_pad;
  wire [12:0] cfiType_21_shl;
  wire [19:0] cfiType_21_pad;
  wire [17:0] tgtPages_4_shl;
  wire [19:0] tgtPages_4_pad;
  wire [17:0] tgtPages_6_shl;
  wire [19:0] tgtPages_6_pad;
  wire [17:0] tgtPages_11_shl;
  wire [19:0] tgtPages_11_pad;
  wire [17:0] tgtPages_7_shl;
  wire [19:0] tgtPages_7_pad;
  wire [17:0] tgtPages_20_shl;
  wire [19:0] tgtPages_20_pad;
  wire [12:0] cfiType_3_shl;
  wire [19:0] cfiType_3_pad;
  wire [17:0] tgtPages_16_shl;
  wire [19:0] tgtPages_16_pad;
  wire [12:0] cfiType_24_shl;
  wire [19:0] cfiType_24_pad;
  wire [17:0] tgtPages_17_shl;
  wire [19:0] tgtPages_17_pad;
  wire [12:0] cfiType_6_shl;
  wire [19:0] cfiType_6_pad;
  wire [17:0] tgtPages_9_shl;
  wire [19:0] tgtPages_9_pad;
  wire [17:0] tgtPages_2_shl;
  wire [19:0] tgtPages_2_pad;
  wire [12:0] cfiType_10_shl;
  wire [19:0] cfiType_10_pad;
  wire [17:0] tgtPages_18_shl;
  wire [19:0] tgtPages_18_pad;
  wire [17:0] tgtPages_0_shl;
  wire [19:0] tgtPages_0_pad;
  wire [17:0] tgtPages_25_shl;
  wire [19:0] tgtPages_25_pad;
  wire [17:0] tgtPages_22_shl;
  wire [19:0] tgtPages_22_pad;
  wire [12:0] cfiType_5_shl;
  wire [19:0] cfiType_5_pad;
  wire [12:0] cfiType_12_shl;
  wire [19:0] cfiType_12_pad;
  wire [12:0] cfiType_18_shl;
  wire [19:0] cfiType_18_pad;
  wire [17:0] tgtPages_24_shl;
  wire [19:0] tgtPages_24_pad;
  wire [17:0] tgtPages_26_shl;
  wire [19:0] tgtPages_26_pad;
  wire [17:0] tgtPages_1_shl;
  wire [19:0] tgtPages_1_pad;
  wire [17:0] tgtPages_10_shl;
  wire [19:0] tgtPages_10_pad;
  wire [12:0] cfiType_25_shl;
  wire [19:0] cfiType_25_pad;
  wire [12:0] cfiType_16_shl;
  wire [19:0] cfiType_16_pad;
  wire [17:0] tgtPages_13_shl;
  wire [19:0] tgtPages_13_pad;
  wire [12:0] cfiType_19_shl;
  wire [19:0] cfiType_19_pad;
  wire [12:0] cfiType_2_shl;
  wire [19:0] cfiType_2_pad;
  wire [12:0] cfiType_20_shl;
  wire [19:0] cfiType_20_pad;
  wire [17:0] tgtPages_15_shl;
  wire [19:0] tgtPages_15_pad;
  wire [17:0] tgtPages_8_shl;
  wire [19:0] tgtPages_8_pad;
  wire [17:0] tgtPages_5_shl;
  wire [19:0] tgtPages_5_pad;
  wire [12:0] cfiType_0_shl;
  wire [19:0] cfiType_0_pad;
  wire [17:0] tgtPages_3_shl;
  wire [19:0] tgtPages_3_pad;
  wire [17:0] tgtPages_27_shl;
  wire [19:0] tgtPages_27_pad;
  wire [12:0] cfiType_27_shl;
  wire [19:0] cfiType_27_pad;
  wire [17:0] tgtPages_14_shl;
  wire [19:0] tgtPages_14_pad;
  wire [12:0] cfiType_13_shl;
  wire [19:0] cfiType_13_pad;
  wire [12:0] cfiType_23_shl;
  wire [19:0] cfiType_23_pad;
  wire [12:0] cfiType_4_shl;
  wire [19:0] cfiType_4_pad;
  wire [12:0] cfiType_1_shl;
  wire [19:0] cfiType_1_pad;
  wire [17:0] tgtPages_21_shl;
  wire [19:0] tgtPages_21_pad;
  wire [12:0] cfiType_8_shl;
  wire [19:0] cfiType_8_pad;
  wire [17:0] tgtPages_23_shl;
  wire [19:0] tgtPages_23_pad;
  wire [17:0] tgtPages_19_shl;
  wire [19:0] tgtPages_19_pad;
  wire [12:0] cfiType_11_shl;
  wire [19:0] cfiType_11_pad;
  wire [17:0] tgtPages_12_shl;
  wire [19:0] tgtPages_12_pad;
  wire [12:0] cfiType_9_shl;
  wire [19:0] cfiType_9_pad;
  wire [12:0] cfiType_14_shl;
  wire [19:0] cfiType_14_pad;
  wire [12:0] cfiType_7_shl;
  wire [19:0] cfiType_7_pad;
  wire [12:0] cfiType_26_shl;
  wire [19:0] cfiType_26_pad;
  wire [12:0] cfiType_15_shl;
  wire [19:0] cfiType_15_pad;
  wire [19:0] BTB_xor31;
  wire [19:0] BTB_xor66;
  wire [19:0] BTB_xor32;
  wire [19:0] BTB_xor15;
  wire [19:0] BTB_xor68;
  wire [19:0] BTB_xor33;
  wire [19:0] BTB_xor70;
  wire [19:0] BTB_xor34;
  wire [19:0] BTB_xor16;
  wire [19:0] BTB_xor7;
  wire [19:0] BTB_xor72;
  wire [19:0] BTB_xor35;
  wire [19:0] BTB_xor74;
  wire [19:0] BTB_xor36;
  wire [19:0] BTB_xor17;
  wire [19:0] BTB_xor76;
  wire [19:0] BTB_xor37;
  wire [19:0] BTB_xor78;
  wire [19:0] BTB_xor38;
  wire [19:0] BTB_xor18;
  wire [19:0] BTB_xor8;
  wire [19:0] BTB_xor3;
  wire [19:0] BTB_xor39;
  wire [19:0] BTB_xor82;
  wire [19:0] BTB_xor40;
  wire [19:0] BTB_xor19;
  wire [19:0] BTB_xor84;
  wire [19:0] BTB_xor41;
  wire [19:0] BTB_xor86;
  wire [19:0] BTB_xor42;
  wire [19:0] BTB_xor20;
  wire [19:0] BTB_xor9;
  wire [19:0] BTB_xor88;
  wire [19:0] BTB_xor43;
  wire [19:0] BTB_xor90;
  wire [19:0] BTB_xor44;
  wire [19:0] BTB_xor21;
  wire [19:0] BTB_xor92;
  wire [19:0] BTB_xor45;
  wire [19:0] BTB_xor94;
  wire [19:0] BTB_xor46;
  wire [19:0] BTB_xor22;
  wire [19:0] BTB_xor10;
  wire [19:0] BTB_xor4;
  wire [19:0] BTB_xor1;
  wire [19:0] BTB_xor47;
  wire [19:0] BTB_xor98;
  wire [19:0] BTB_xor48;
  wire [19:0] BTB_xor23;
  wire [19:0] BTB_xor100;
  wire [19:0] BTB_xor49;
  wire [19:0] BTB_xor102;
  wire [19:0] BTB_xor50;
  wire [19:0] BTB_xor24;
  wire [19:0] BTB_xor11;
  wire [19:0] BTB_xor104;
  wire [19:0] BTB_xor51;
  wire [19:0] BTB_xor106;
  wire [19:0] BTB_xor52;
  wire [19:0] BTB_xor25;
  wire [19:0] BTB_xor108;
  wire [19:0] BTB_xor53;
  wire [19:0] BTB_xor110;
  wire [19:0] BTB_xor54;
  wire [19:0] BTB_xor26;
  wire [19:0] BTB_xor12;
  wire [19:0] BTB_xor5;
  wire [19:0] BTB_xor112;
  wire [19:0] BTB_xor55;
  wire [19:0] BTB_xor114;
  wire [19:0] BTB_xor56;
  wire [19:0] BTB_xor27;
  wire [19:0] BTB_xor116;
  wire [19:0] BTB_xor57;
  wire [19:0] BTB_xor118;
  wire [19:0] BTB_xor58;
  wire [19:0] BTB_xor28;
  wire [19:0] BTB_xor13;
  wire [19:0] BTB_xor120;
  wire [19:0] BTB_xor59;
  wire [19:0] BTB_xor122;
  wire [19:0] BTB_xor60;
  wire [19:0] BTB_xor29;
  wire [19:0] BTB_xor124;
  wire [19:0] BTB_xor61;
  wire [19:0] BTB_xor126;
  wire [19:0] BTB_xor62;
  wire [19:0] BTB_xor30;
  wire [19:0] BTB_xor14;
  wire [19:0] BTB_xor6;
  wire [19:0] BTB_xor2;
  wire [19:0] BTB_xor0;
  assign table__res_res_value_MPORT_addr = _res_res_value_T_3 ^ _res_res_value_T_6;
  assign table__res_res_value_MPORT_data = table_[table__res_res_value_MPORT_addr]; // @[BTB.scala 118:26]
  assign table__MPORT_data = io_bht_update_valid & _GEN_389;
  assign table__MPORT_addr = waddr_1[8:0];
  assign table__MPORT_mask = 1'h1;
  assign table__MPORT_en = io_bht_update_valid ? _GEN_387 : resetting;
  assign pagesMasked_0 = pageValid[0] ? pages_0 : 25'h0; // @[BTB.scala 207:75]
  assign pagesMasked_1 = pageValid[1] ? pages_1 : 25'h0; // @[BTB.scala 207:75]
  assign pagesMasked_2 = pageValid[2] ? pages_2 : 25'h0; // @[BTB.scala 207:75]
  assign pagesMasked_3 = pageValid[3] ? pages_3 : 25'h0; // @[BTB.scala 207:75]
  assign pagesMasked_4 = pageValid[4] ? pages_4 : 25'h0; // @[BTB.scala 207:75]
  assign pagesMasked_5 = pageValid[5] ? pages_5 : 25'h0; // @[BTB.scala 207:75]
  assign pageHit_p = io_req_bits_addr[38:14]; // @[BTB.scala 213:39]
  assign pageHit_lo_lo = pages_0 == pageHit_p; // @[BTB.scala 216:29]
  assign pageHit_lo_hi_lo = pages_1 == pageHit_p; // @[BTB.scala 216:29]
  assign pageHit_lo_hi_hi = pages_2 == pageHit_p; // @[BTB.scala 216:29]
  assign pageHit_hi_lo = pages_3 == pageHit_p; // @[BTB.scala 216:29]
  assign pageHit_hi_hi_lo = pages_4 == pageHit_p; // @[BTB.scala 216:29]
  assign pageHit_hi_hi_hi = pages_5 == pageHit_p; // @[BTB.scala 216:29]
  assign _pageHit_T = {pageHit_hi_hi_hi,pageHit_hi_hi_lo,pageHit_hi_lo,pageHit_lo_hi_hi,pageHit_lo_hi_lo,pageHit_lo_lo}; // @[Cat.scala 30:58]
  assign pageHit = pageValid & _pageHit_T; // @[BTB.scala 216:15]
  assign idxHit_idx = io_req_bits_addr[13:1]; // @[BTB.scala 219:19]
  assign idxHit_lo_lo_lo_lo = idxs_0 == idxHit_idx; // @[BTB.scala 220:16]
  assign idxHit_lo_lo_lo_hi_lo = idxs_1 == idxHit_idx; // @[BTB.scala 220:16]
  assign idxHit_lo_lo_lo_hi_hi = idxs_2 == idxHit_idx; // @[BTB.scala 220:16]
  assign idxHit_lo_lo_hi_lo_lo = idxs_3 == idxHit_idx; // @[BTB.scala 220:16]
  assign idxHit_lo_lo_hi_lo_hi = idxs_4 == idxHit_idx; // @[BTB.scala 220:16]
  assign idxHit_lo_lo_hi_hi_lo = idxs_5 == idxHit_idx; // @[BTB.scala 220:16]
  assign idxHit_lo_lo_hi_hi_hi = idxs_6 == idxHit_idx; // @[BTB.scala 220:16]
  assign idxHit_lo_hi_lo_lo = idxs_7 == idxHit_idx; // @[BTB.scala 220:16]
  assign idxHit_lo_hi_lo_hi_lo = idxs_8 == idxHit_idx; // @[BTB.scala 220:16]
  assign idxHit_lo_hi_lo_hi_hi = idxs_9 == idxHit_idx; // @[BTB.scala 220:16]
  assign idxHit_lo_hi_hi_lo_lo = idxs_10 == idxHit_idx; // @[BTB.scala 220:16]
  assign idxHit_lo_hi_hi_lo_hi = idxs_11 == idxHit_idx; // @[BTB.scala 220:16]
  assign idxHit_lo_hi_hi_hi_lo = idxs_12 == idxHit_idx; // @[BTB.scala 220:16]
  assign idxHit_lo_hi_hi_hi_hi = idxs_13 == idxHit_idx; // @[BTB.scala 220:16]
  assign idxHit_hi_lo_lo_lo = idxs_14 == idxHit_idx; // @[BTB.scala 220:16]
  assign idxHit_hi_lo_lo_hi_lo = idxs_15 == idxHit_idx; // @[BTB.scala 220:16]
  assign idxHit_hi_lo_lo_hi_hi = idxs_16 == idxHit_idx; // @[BTB.scala 220:16]
  assign idxHit_hi_lo_hi_lo_lo = idxs_17 == idxHit_idx; // @[BTB.scala 220:16]
  assign idxHit_hi_lo_hi_lo_hi = idxs_18 == idxHit_idx; // @[BTB.scala 220:16]
  assign idxHit_hi_lo_hi_hi_lo = idxs_19 == idxHit_idx; // @[BTB.scala 220:16]
  assign idxHit_hi_lo_hi_hi_hi = idxs_20 == idxHit_idx; // @[BTB.scala 220:16]
  assign idxHit_hi_hi_lo_lo = idxs_21 == idxHit_idx; // @[BTB.scala 220:16]
  assign idxHit_hi_hi_lo_hi_lo = idxs_22 == idxHit_idx; // @[BTB.scala 220:16]
  assign idxHit_hi_hi_lo_hi_hi = idxs_23 == idxHit_idx; // @[BTB.scala 220:16]
  assign idxHit_hi_hi_hi_lo_lo = idxs_24 == idxHit_idx; // @[BTB.scala 220:16]
  assign idxHit_hi_hi_hi_lo_hi = idxs_25 == idxHit_idx; // @[BTB.scala 220:16]
  assign idxHit_hi_hi_hi_hi_lo = idxs_26 == idxHit_idx; // @[BTB.scala 220:16]
  assign idxHit_hi_hi_hi_hi_hi = idxs_27 == idxHit_idx; // @[BTB.scala 220:16]
  assign idxHit_lo_lo = {idxHit_lo_lo_hi_hi_hi,idxHit_lo_lo_hi_hi_lo,idxHit_lo_lo_hi_lo_hi,idxHit_lo_lo_hi_lo_lo,idxHit_lo_lo_lo_hi_hi,idxHit_lo_lo_lo_hi_lo,idxHit_lo_lo_lo_lo}; // @[Cat.scala 30:58]
  assign idxHit_lo = {idxHit_lo_hi_hi_hi_hi,idxHit_lo_hi_hi_hi_lo,idxHit_lo_hi_hi_lo_hi,idxHit_lo_hi_hi_lo_lo,idxHit_lo_hi_lo_hi_hi,idxHit_lo_hi_lo_hi_lo,idxHit_lo_hi_lo_lo,idxHit_lo_lo}; // @[Cat.scala 30:58]
  assign idxHit_hi_lo = {idxHit_hi_lo_hi_hi_hi,idxHit_hi_lo_hi_hi_lo,idxHit_hi_lo_hi_lo_hi,idxHit_hi_lo_hi_lo_lo,idxHit_hi_lo_lo_hi_hi,idxHit_hi_lo_lo_hi_lo,idxHit_hi_lo_lo_lo}; // @[Cat.scala 30:58]
  assign _idxHit_T = {idxHit_hi_hi_hi_hi_hi,idxHit_hi_hi_hi_hi_lo,idxHit_hi_hi_hi_lo_hi,idxHit_hi_hi_hi_lo_lo,idxHit_hi_hi_lo_hi_hi,idxHit_hi_hi_lo_hi_lo,idxHit_hi_hi_lo_lo,idxHit_hi_lo,idxHit_lo}; // @[Cat.scala 30:58]
  assign idxHit = _idxHit_T & isValid; // @[BTB.scala 220:32]
  assign updatePageHit_p = r_btb_updatePipe_bits_pc[38:14]; // @[BTB.scala 213:39]
  assign updatePageHit_lo_lo = pages_0 == updatePageHit_p; // @[BTB.scala 216:29]
  assign updatePageHit_lo_hi_lo = pages_1 == updatePageHit_p; // @[BTB.scala 216:29]
  assign updatePageHit_lo_hi_hi = pages_2 == updatePageHit_p; // @[BTB.scala 216:29]
  assign updatePageHit_hi_lo = pages_3 == updatePageHit_p; // @[BTB.scala 216:29]
  assign updatePageHit_hi_hi_lo = pages_4 == updatePageHit_p; // @[BTB.scala 216:29]
  assign updatePageHit_hi_hi_hi = pages_5 == updatePageHit_p; // @[BTB.scala 216:29]
  assign _updatePageHit_T = {updatePageHit_hi_hi_hi,updatePageHit_hi_hi_lo,updatePageHit_hi_lo,updatePageHit_lo_hi_hi,updatePageHit_lo_hi_lo,updatePageHit_lo_lo}; // @[Cat.scala 30:58]
  assign updatePageHit = pageValid & _updatePageHit_T; // @[BTB.scala 216:15]
  assign updateHit = r_btb_updatePipe_bits_prediction_entry < 5'h1c; // @[BTB.scala 234:48]
  assign useUpdatePageHit = |updatePageHit; // @[BTB.scala 236:40]
  assign usePageHit = |pageHit; // @[BTB.scala 237:28]
  assign doIdxPageRepl = ~useUpdatePageHit; // @[BTB.scala 238:23]
  assign idxPageRepl_hi = pageHit[4:0]; // @[BTB.scala 240:32]
  assign idxPageRepl_lo = pageHit[5]; // @[BTB.scala 240:53]
  assign _idxPageRepl_T = {idxPageRepl_hi,idxPageRepl_lo}; // @[Cat.scala 30:58]
  assign _idxPageRepl_T_1 = 8'h1 << nextPageRepl; // @[OneHot.scala 58:35]
  assign _idxPageRepl_T_2 = usePageHit ? 8'h0 : _idxPageRepl_T_1; // @[BTB.scala 240:70]
  assign _GEN_430 = {{2'd0}, _idxPageRepl_T}; // @[BTB.scala 240:65]
  assign idxPageRepl = _GEN_430 | _idxPageRepl_T_2; // @[BTB.scala 240:65]
  assign idxPageUpdateOH = useUpdatePageHit ? {{2'd0}, updatePageHit} : idxPageRepl; // @[BTB.scala 241:28]
  assign idxPageUpdate_hi = idxPageUpdateOH[7:4]; // @[OneHot.scala 30:18]
  assign idxPageUpdate_lo = idxPageUpdateOH[3:0]; // @[OneHot.scala 31:18]
  assign idxPageUpdate_hi_1 = |idxPageUpdate_hi; // @[OneHot.scala 32:14]
  assign _idxPageUpdate_T = idxPageUpdate_hi | idxPageUpdate_lo; // @[OneHot.scala 32:28]
  assign idxPageUpdate_hi_2 = _idxPageUpdate_T[3:2]; // @[OneHot.scala 30:18]
  assign idxPageUpdate_lo_1 = _idxPageUpdate_T[1:0]; // @[OneHot.scala 31:18]
  assign idxPageUpdate_hi_3 = |idxPageUpdate_hi_2; // @[OneHot.scala 32:14]
  assign _idxPageUpdate_T_1 = idxPageUpdate_hi_2 | idxPageUpdate_lo_1; // @[OneHot.scala 32:28]
  assign idxPageUpdate_lo_2 = _idxPageUpdate_T_1[1]; // @[CircuitMath.scala 30:8]
  assign idxPageUpdate = {idxPageUpdate_hi_1,idxPageUpdate_hi_3,idxPageUpdate_lo_2}; // @[Cat.scala 30:58]
  assign idxPageReplEn = doIdxPageRepl ? idxPageRepl : 8'h0; // @[BTB.scala 243:26]
  assign samePage = updatePageHit_p == pageHit_p; // @[BTB.scala 245:45]
  assign doTgtPageRepl = ~samePage & ~usePageHit; // @[BTB.scala 246:33]
  assign tgtPageRepl_hi = idxPageUpdateOH[4:0]; // @[BTB.scala 247:71]
  assign tgtPageRepl_lo = idxPageUpdateOH[5]; // @[BTB.scala 247:100]
  assign _tgtPageRepl_T = {tgtPageRepl_hi,tgtPageRepl_lo}; // @[Cat.scala 30:58]
  assign tgtPageRepl = samePage ? idxPageUpdateOH : {{2'd0}, _tgtPageRepl_T}; // @[BTB.scala 247:24]
  assign _tgtPageUpdate_T = usePageHit ? 8'h0 : tgtPageRepl; // @[BTB.scala 248:45]
  assign _GEN_431 = {{2'd0}, pageHit}; // @[BTB.scala 248:40]
  assign _tgtPageUpdate_T_1 = _GEN_431 | _tgtPageUpdate_T; // @[BTB.scala 248:40]
  assign tgtPageUpdate_hi = _tgtPageUpdate_T_1[7:4]; // @[OneHot.scala 30:18]
  assign tgtPageUpdate_lo = _tgtPageUpdate_T_1[3:0]; // @[OneHot.scala 31:18]
  assign tgtPageUpdate_hi_1 = |tgtPageUpdate_hi; // @[OneHot.scala 32:14]
  assign _tgtPageUpdate_T_2 = tgtPageUpdate_hi | tgtPageUpdate_lo; // @[OneHot.scala 32:28]
  assign tgtPageUpdate_hi_2 = _tgtPageUpdate_T_2[3:2]; // @[OneHot.scala 30:18]
  assign tgtPageUpdate_lo_1 = _tgtPageUpdate_T_2[1:0]; // @[OneHot.scala 31:18]
  assign tgtPageUpdate_hi_3 = |tgtPageUpdate_hi_2; // @[OneHot.scala 32:14]
  assign _tgtPageUpdate_T_3 = tgtPageUpdate_hi_2 | tgtPageUpdate_lo_1; // @[OneHot.scala 32:28]
  assign tgtPageUpdate_lo_2 = _tgtPageUpdate_T_3[1]; // @[CircuitMath.scala 30:8]
  assign tgtPageUpdate = {tgtPageUpdate_hi_1,tgtPageUpdate_hi_3,tgtPageUpdate_lo_2}; // @[Cat.scala 30:58]
  assign tgtPageReplEn = doTgtPageRepl ? tgtPageRepl : 8'h0; // @[BTB.scala 249:26]
  assign _T = doIdxPageRepl | doTgtPageRepl; // @[BTB.scala 251:46]
  assign _T_1 = r_btb_updatePipe_valid & _T; // @[BTB.scala 251:28]
  assign both = doIdxPageRepl & doTgtPageRepl; // @[BTB.scala 252:30]
  assign _next_T = both ? 2'h2 : 2'h1; // @[BTB.scala 253:40]
  assign _GEN_432 = {{1'd0}, _next_T}; // @[BTB.scala 253:29]
  assign next = nextPageRepl + _GEN_432; // @[BTB.scala 253:29]
  assign _nextPageRepl_T = next >= 3'h6; // @[BTB.scala 254:30]
  assign waddr_hi = state_reg[26]; // @[Replacement.scala 243:38]
  assign waddr_left_subtree_state = state_reg[25:15]; // @[package.scala 154:13]
  assign waddr_right_subtree_state = state_reg[14:0]; // @[Replacement.scala 245:38]
  assign waddr_hi_1 = waddr_left_subtree_state[10]; // @[Replacement.scala 243:38]
  assign waddr_left_subtree_state_1 = waddr_left_subtree_state[9:7]; // @[package.scala 154:13]
  assign waddr_right_subtree_state_1 = waddr_left_subtree_state[6:0]; // @[Replacement.scala 245:38]
  assign waddr_hi_2 = waddr_left_subtree_state_1[2]; // @[Replacement.scala 243:38]
  assign waddr_left_subtree_state_2 = waddr_left_subtree_state_1[1]; // @[package.scala 154:13]
  assign waddr_right_subtree_state_2 = waddr_left_subtree_state_1[0]; // @[Replacement.scala 245:38]
  assign waddr_lo = waddr_hi_2 ? waddr_left_subtree_state_2 : waddr_right_subtree_state_2; // @[Replacement.scala 250:16]
  assign _waddr_T_2 = {waddr_hi_2,waddr_lo}; // @[Cat.scala 30:58]
  assign waddr_hi_3 = waddr_right_subtree_state_1[6]; // @[Replacement.scala 243:38]
  assign waddr_left_subtree_state_3 = waddr_right_subtree_state_1[5:3]; // @[package.scala 154:13]
  assign waddr_right_subtree_state_3 = waddr_right_subtree_state_1[2:0]; // @[Replacement.scala 245:38]
  assign waddr_hi_4 = waddr_left_subtree_state_3[2]; // @[Replacement.scala 243:38]
  assign waddr_left_subtree_state_4 = waddr_left_subtree_state_3[1]; // @[package.scala 154:13]
  assign waddr_right_subtree_state_4 = waddr_left_subtree_state_3[0]; // @[Replacement.scala 245:38]
  assign waddr_lo_1 = waddr_hi_4 ? waddr_left_subtree_state_4 : waddr_right_subtree_state_4; // @[Replacement.scala 250:16]
  assign _waddr_T_5 = {waddr_hi_4,waddr_lo_1}; // @[Cat.scala 30:58]
  assign waddr_hi_5 = waddr_right_subtree_state_3[2]; // @[Replacement.scala 243:38]
  assign waddr_left_subtree_state_5 = waddr_right_subtree_state_3[1]; // @[package.scala 154:13]
  assign waddr_right_subtree_state_5 = waddr_right_subtree_state_3[0]; // @[Replacement.scala 245:38]
  assign waddr_lo_2 = waddr_hi_5 ? waddr_left_subtree_state_5 : waddr_right_subtree_state_5; // @[Replacement.scala 250:16]
  assign _waddr_T_8 = {waddr_hi_5,waddr_lo_2}; // @[Cat.scala 30:58]
  assign waddr_lo_3 = waddr_hi_3 ? _waddr_T_5 : _waddr_T_8; // @[Replacement.scala 250:16]
  assign _waddr_T_9 = {waddr_hi_3,waddr_lo_3}; // @[Cat.scala 30:58]
  assign waddr_lo_4 = waddr_hi_1 ? {{1'd0}, _waddr_T_2} : _waddr_T_9; // @[Replacement.scala 250:16]
  assign _waddr_T_10 = {waddr_hi_1,waddr_lo_4}; // @[Cat.scala 30:58]
  assign waddr_hi_6 = waddr_right_subtree_state[14]; // @[Replacement.scala 243:38]
  assign waddr_left_subtree_state_6 = waddr_right_subtree_state[13:7]; // @[package.scala 154:13]
  assign waddr_right_subtree_state_6 = waddr_right_subtree_state[6:0]; // @[Replacement.scala 245:38]
  assign waddr_hi_7 = waddr_left_subtree_state_6[6]; // @[Replacement.scala 243:38]
  assign waddr_left_subtree_state_7 = waddr_left_subtree_state_6[5:3]; // @[package.scala 154:13]
  assign waddr_right_subtree_state_7 = waddr_left_subtree_state_6[2:0]; // @[Replacement.scala 245:38]
  assign waddr_hi_8 = waddr_left_subtree_state_7[2]; // @[Replacement.scala 243:38]
  assign waddr_left_subtree_state_8 = waddr_left_subtree_state_7[1]; // @[package.scala 154:13]
  assign waddr_right_subtree_state_8 = waddr_left_subtree_state_7[0]; // @[Replacement.scala 245:38]
  assign waddr_lo_5 = waddr_hi_8 ? waddr_left_subtree_state_8 : waddr_right_subtree_state_8; // @[Replacement.scala 250:16]
  assign _waddr_T_13 = {waddr_hi_8,waddr_lo_5}; // @[Cat.scala 30:58]
  assign waddr_hi_9 = waddr_right_subtree_state_7[2]; // @[Replacement.scala 243:38]
  assign waddr_left_subtree_state_9 = waddr_right_subtree_state_7[1]; // @[package.scala 154:13]
  assign waddr_right_subtree_state_9 = waddr_right_subtree_state_7[0]; // @[Replacement.scala 245:38]
  assign waddr_lo_6 = waddr_hi_9 ? waddr_left_subtree_state_9 : waddr_right_subtree_state_9; // @[Replacement.scala 250:16]
  assign _waddr_T_16 = {waddr_hi_9,waddr_lo_6}; // @[Cat.scala 30:58]
  assign waddr_lo_7 = waddr_hi_7 ? _waddr_T_13 : _waddr_T_16; // @[Replacement.scala 250:16]
  assign _waddr_T_17 = {waddr_hi_7,waddr_lo_7}; // @[Cat.scala 30:58]
  assign waddr_hi_10 = waddr_right_subtree_state_6[6]; // @[Replacement.scala 243:38]
  assign waddr_left_subtree_state_10 = waddr_right_subtree_state_6[5:3]; // @[package.scala 154:13]
  assign waddr_right_subtree_state_10 = waddr_right_subtree_state_6[2:0]; // @[Replacement.scala 245:38]
  assign waddr_hi_11 = waddr_left_subtree_state_10[2]; // @[Replacement.scala 243:38]
  assign waddr_left_subtree_state_11 = waddr_left_subtree_state_10[1]; // @[package.scala 154:13]
  assign waddr_right_subtree_state_11 = waddr_left_subtree_state_10[0]; // @[Replacement.scala 245:38]
  assign waddr_lo_8 = waddr_hi_11 ? waddr_left_subtree_state_11 : waddr_right_subtree_state_11; // @[Replacement.scala 250:16]
  assign _waddr_T_20 = {waddr_hi_11,waddr_lo_8}; // @[Cat.scala 30:58]
  assign waddr_hi_12 = waddr_right_subtree_state_10[2]; // @[Replacement.scala 243:38]
  assign waddr_left_subtree_state_12 = waddr_right_subtree_state_10[1]; // @[package.scala 154:13]
  assign waddr_right_subtree_state_12 = waddr_right_subtree_state_10[0]; // @[Replacement.scala 245:38]
  assign waddr_lo_9 = waddr_hi_12 ? waddr_left_subtree_state_12 : waddr_right_subtree_state_12; // @[Replacement.scala 250:16]
  assign _waddr_T_23 = {waddr_hi_12,waddr_lo_9}; // @[Cat.scala 30:58]
  assign waddr_lo_10 = waddr_hi_10 ? _waddr_T_20 : _waddr_T_23; // @[Replacement.scala 250:16]
  assign _waddr_T_24 = {waddr_hi_10,waddr_lo_10}; // @[Cat.scala 30:58]
  assign waddr_lo_11 = waddr_hi_6 ? _waddr_T_17 : _waddr_T_24; // @[Replacement.scala 250:16]
  assign _waddr_T_25 = {waddr_hi_6,waddr_lo_11}; // @[Cat.scala 30:58]
  assign waddr_lo_12 = waddr_hi ? _waddr_T_10 : _waddr_T_25; // @[Replacement.scala 250:16]
  assign _waddr_T_26 = {waddr_hi,waddr_lo_12}; // @[Cat.scala 30:58]
  assign waddr = updateHit ? r_btb_updatePipe_bits_prediction_entry : _waddr_T_26; // @[BTB.scala 258:18]
  assign _T_2 = r_respPipe_valid & r_respPipe_bits_taken; // @[BTB.scala 260:22]
  assign _T_3 = _T_2 | r_btb_updatePipe_valid; // @[BTB.scala 260:43]
  assign state_reg_touch_way_sized = r_btb_updatePipe_valid ? waddr : r_respPipe_bits_entry; // @[BTB.scala 261:20]
  assign state_reg_hi_hi = ~state_reg_touch_way_sized[4]; // @[Replacement.scala 196:33]
  assign state_reg_hi_hi_1 = ~state_reg_touch_way_sized[3]; // @[Replacement.scala 196:33]
  assign state_reg_hi_hi_2 = ~state_reg_touch_way_sized[1]; // @[Replacement.scala 196:33]
  assign state_reg_hi_lo = state_reg_hi_hi_2 ? waddr_left_subtree_state_2 : ~state_reg_touch_way_sized[0]; // @[Replacement.scala 203:16]
  assign state_reg_lo = state_reg_hi_hi_2 ? ~state_reg_touch_way_sized[0] : waddr_right_subtree_state_2; // @[Replacement.scala 206:16]
  assign _state_reg_T_8 = {state_reg_hi_hi_2,state_reg_hi_lo,state_reg_lo}; // @[Cat.scala 30:58]
  assign state_reg_hi_lo_1 = state_reg_hi_hi_1 ? waddr_left_subtree_state_1 : _state_reg_T_8; // @[Replacement.scala 203:16]
  assign state_reg_hi_hi_3 = ~state_reg_touch_way_sized[2]; // @[Replacement.scala 196:33]
  assign state_reg_hi_hi_4 = ~state_reg_touch_way_sized[1]; // @[Replacement.scala 196:33]
  assign state_reg_hi_lo_2 = state_reg_hi_hi_4 ? waddr_left_subtree_state_4 : ~state_reg_touch_way_sized[0]; // @[Replacement.scala 203:16]
  assign state_reg_lo_1 = state_reg_hi_hi_4 ? ~state_reg_touch_way_sized[0] : waddr_right_subtree_state_4; // @[Replacement.scala 206:16]
  assign _state_reg_T_17 = {state_reg_hi_hi_4,state_reg_hi_lo_2,state_reg_lo_1}; // @[Cat.scala 30:58]
  assign state_reg_hi_lo_3 = state_reg_hi_hi_3 ? waddr_left_subtree_state_3 : _state_reg_T_17; // @[Replacement.scala 203:16]
  assign state_reg_hi_lo_4 = state_reg_hi_hi_4 ? waddr_left_subtree_state_5 : ~state_reg_touch_way_sized[0]; // @[Replacement.scala 203:16]
  assign state_reg_lo_2 = state_reg_hi_hi_4 ? ~state_reg_touch_way_sized[0] : waddr_right_subtree_state_5; // @[Replacement.scala 206:16]
  assign _state_reg_T_25 = {state_reg_hi_hi_4,state_reg_hi_lo_4,state_reg_lo_2}; // @[Cat.scala 30:58]
  assign state_reg_lo_3 = state_reg_hi_hi_3 ? _state_reg_T_25 : waddr_right_subtree_state_3; // @[Replacement.scala 206:16]
  assign _state_reg_T_26 = {state_reg_hi_hi_3,state_reg_hi_lo_3,state_reg_lo_3}; // @[Cat.scala 30:58]
  assign state_reg_lo_4 = state_reg_hi_hi_1 ? _state_reg_T_26 : waddr_right_subtree_state_1; // @[Replacement.scala 206:16]
  assign _state_reg_T_27 = {state_reg_hi_hi_1,state_reg_hi_lo_1,state_reg_lo_4}; // @[Cat.scala 30:58]
  assign state_reg_hi_lo_5 = state_reg_hi_hi ? waddr_left_subtree_state : _state_reg_T_27; // @[Replacement.scala 203:16]
  assign state_reg_hi_lo_6 = state_reg_hi_hi_4 ? waddr_left_subtree_state_8 : ~state_reg_touch_way_sized[0]; // @[Replacement.scala 203:16]
  assign state_reg_lo_5 = state_reg_hi_hi_4 ? ~state_reg_touch_way_sized[0] : waddr_right_subtree_state_8; // @[Replacement.scala 206:16]
  assign _state_reg_T_37 = {state_reg_hi_hi_4,state_reg_hi_lo_6,state_reg_lo_5}; // @[Cat.scala 30:58]
  assign state_reg_hi_lo_7 = state_reg_hi_hi_3 ? waddr_left_subtree_state_7 : _state_reg_T_37; // @[Replacement.scala 203:16]
  assign state_reg_hi_lo_8 = state_reg_hi_hi_4 ? waddr_left_subtree_state_9 : ~state_reg_touch_way_sized[0]; // @[Replacement.scala 203:16]
  assign state_reg_lo_6 = state_reg_hi_hi_4 ? ~state_reg_touch_way_sized[0] : waddr_right_subtree_state_9; // @[Replacement.scala 206:16]
  assign _state_reg_T_45 = {state_reg_hi_hi_4,state_reg_hi_lo_8,state_reg_lo_6}; // @[Cat.scala 30:58]
  assign state_reg_lo_7 = state_reg_hi_hi_3 ? _state_reg_T_45 : waddr_right_subtree_state_7; // @[Replacement.scala 206:16]
  assign _state_reg_T_46 = {state_reg_hi_hi_3,state_reg_hi_lo_7,state_reg_lo_7}; // @[Cat.scala 30:58]
  assign state_reg_hi_lo_9 = state_reg_hi_hi_1 ? waddr_left_subtree_state_6 : _state_reg_T_46; // @[Replacement.scala 203:16]
  assign state_reg_hi_lo_10 = state_reg_hi_hi_4 ? waddr_left_subtree_state_11 : ~state_reg_touch_way_sized[0]; // @[Replacement.scala 203:16]
  assign state_reg_lo_8 = state_reg_hi_hi_4 ? ~state_reg_touch_way_sized[0] : waddr_right_subtree_state_11; // @[Replacement.scala 206:16]
  assign _state_reg_T_55 = {state_reg_hi_hi_4,state_reg_hi_lo_10,state_reg_lo_8}; // @[Cat.scala 30:58]
  assign state_reg_hi_lo_11 = state_reg_hi_hi_3 ? waddr_left_subtree_state_10 : _state_reg_T_55; // @[Replacement.scala 203:16]
  assign state_reg_hi_lo_12 = state_reg_hi_hi_4 ? waddr_left_subtree_state_12 : ~state_reg_touch_way_sized[0]; // @[Replacement.scala 203:16]
  assign state_reg_lo_9 = state_reg_hi_hi_4 ? ~state_reg_touch_way_sized[0] : waddr_right_subtree_state_12; // @[Replacement.scala 206:16]
  assign _state_reg_T_63 = {state_reg_hi_hi_4,state_reg_hi_lo_12,state_reg_lo_9}; // @[Cat.scala 30:58]
  assign state_reg_lo_10 = state_reg_hi_hi_3 ? _state_reg_T_63 : waddr_right_subtree_state_10; // @[Replacement.scala 206:16]
  assign _state_reg_T_64 = {state_reg_hi_hi_3,state_reg_hi_lo_11,state_reg_lo_10}; // @[Cat.scala 30:58]
  assign state_reg_lo_11 = state_reg_hi_hi_1 ? _state_reg_T_64 : waddr_right_subtree_state_6; // @[Replacement.scala 206:16]
  assign _state_reg_T_65 = {state_reg_hi_hi_1,state_reg_hi_lo_9,state_reg_lo_11}; // @[Cat.scala 30:58]
  assign state_reg_lo_12 = state_reg_hi_hi ? _state_reg_T_65 : waddr_right_subtree_state; // @[Replacement.scala 206:16]
  assign _state_reg_T_66 = {state_reg_hi_hi,state_reg_hi_lo_5,state_reg_lo_12}; // @[Cat.scala 30:58]
  assign mask = 32'h1 << waddr; // @[OneHot.scala 58:35]
  assign _idxPages_T = idxPageUpdate + 3'h1; // @[BTB.scala 268:38]
  assign _GEN_433 = {{4'd0}, isValid}; // @[BTB.scala 271:55]
  assign _isValid_T = _GEN_433 | mask; // @[BTB.scala 271:55]
  assign _isValid_T_2 = _GEN_433 & ~mask; // @[BTB.scala 271:71]
  assign _isValid_T_3 = r_btb_updatePipe_bits_isValid ? _isValid_T : _isValid_T_2; // @[BTB.scala 271:19]
  assign idxWritesEven = ~idxPageUpdate[0]; // @[BTB.scala 276:25]
  assign _T_5 = idxWritesEven ? idxPageReplEn : tgtPageReplEn; // @[BTB.scala 282:24]
  assign _T_12 = idxWritesEven ? tgtPageReplEn : idxPageReplEn; // @[BTB.scala 284:24]
  assign _GEN_435 = {{2'd0}, pageValid}; // @[BTB.scala 286:28]
  assign _pageValid_T = _GEN_435 | tgtPageReplEn; // @[BTB.scala 286:28]
  assign _pageValid_T_1 = _pageValid_T | idxPageReplEn; // @[BTB.scala 286:44]
  assign _GEN_338 = r_btb_updatePipe_valid ? _isValid_T_3 : {{4'd0}, isValid}; // @[BTB.scala 264:29]
  assign _GEN_373 = r_btb_updatePipe_valid ? _pageValid_T_1 : {{2'd0}, pageValid}; // @[BTB.scala 264:29]
  assign _io_resp_valid_T = {pageHit, 1'h0}; // @[BTB.scala 289:29]
  assign _io_resp_valid_T_29 = idxHit[0] ? idxPages_0 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_30 = idxHit[1] ? idxPages_1 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_31 = idxHit[2] ? idxPages_2 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_32 = idxHit[3] ? idxPages_3 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_33 = idxHit[4] ? idxPages_4 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_34 = idxHit[5] ? idxPages_5 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_35 = idxHit[6] ? idxPages_6 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_36 = idxHit[7] ? idxPages_7 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_37 = idxHit[8] ? idxPages_8 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_38 = idxHit[9] ? idxPages_9 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_39 = idxHit[10] ? idxPages_10 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_40 = idxHit[11] ? idxPages_11 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_41 = idxHit[12] ? idxPages_12 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_42 = idxHit[13] ? idxPages_13 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_43 = idxHit[14] ? idxPages_14 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_44 = idxHit[15] ? idxPages_15 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_45 = idxHit[16] ? idxPages_16 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_46 = idxHit[17] ? idxPages_17 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_47 = idxHit[18] ? idxPages_18 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_48 = idxHit[19] ? idxPages_19 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_49 = idxHit[20] ? idxPages_20 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_50 = idxHit[21] ? idxPages_21 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_51 = idxHit[22] ? idxPages_22 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_52 = idxHit[23] ? idxPages_23 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_53 = idxHit[24] ? idxPages_24 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_54 = idxHit[25] ? idxPages_25 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_55 = idxHit[26] ? idxPages_26 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_56 = idxHit[27] ? idxPages_27 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_57 = _io_resp_valid_T_29 | _io_resp_valid_T_30; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_58 = _io_resp_valid_T_57 | _io_resp_valid_T_31; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_59 = _io_resp_valid_T_58 | _io_resp_valid_T_32; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_60 = _io_resp_valid_T_59 | _io_resp_valid_T_33; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_61 = _io_resp_valid_T_60 | _io_resp_valid_T_34; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_62 = _io_resp_valid_T_61 | _io_resp_valid_T_35; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_63 = _io_resp_valid_T_62 | _io_resp_valid_T_36; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_64 = _io_resp_valid_T_63 | _io_resp_valid_T_37; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_65 = _io_resp_valid_T_64 | _io_resp_valid_T_38; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_66 = _io_resp_valid_T_65 | _io_resp_valid_T_39; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_67 = _io_resp_valid_T_66 | _io_resp_valid_T_40; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_68 = _io_resp_valid_T_67 | _io_resp_valid_T_41; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_69 = _io_resp_valid_T_68 | _io_resp_valid_T_42; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_70 = _io_resp_valid_T_69 | _io_resp_valid_T_43; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_71 = _io_resp_valid_T_70 | _io_resp_valid_T_44; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_72 = _io_resp_valid_T_71 | _io_resp_valid_T_45; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_73 = _io_resp_valid_T_72 | _io_resp_valid_T_46; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_74 = _io_resp_valid_T_73 | _io_resp_valid_T_47; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_75 = _io_resp_valid_T_74 | _io_resp_valid_T_48; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_76 = _io_resp_valid_T_75 | _io_resp_valid_T_49; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_77 = _io_resp_valid_T_76 | _io_resp_valid_T_50; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_78 = _io_resp_valid_T_77 | _io_resp_valid_T_51; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_79 = _io_resp_valid_T_78 | _io_resp_valid_T_52; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_80 = _io_resp_valid_T_79 | _io_resp_valid_T_53; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_81 = _io_resp_valid_T_80 | _io_resp_valid_T_54; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_82 = _io_resp_valid_T_81 | _io_resp_valid_T_55; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_83 = _io_resp_valid_T_82 | _io_resp_valid_T_56; // @[Mux.scala 27:72]
  assign _io_resp_valid_T_84 = _io_resp_valid_T >> _io_resp_valid_T_83; // @[BTB.scala 289:34]
  assign _io_resp_bits_target_T_28 = idxHit[0] ? tgtPages_0 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_29 = idxHit[1] ? tgtPages_1 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_30 = idxHit[2] ? tgtPages_2 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_31 = idxHit[3] ? tgtPages_3 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_32 = idxHit[4] ? tgtPages_4 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_33 = idxHit[5] ? tgtPages_5 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_34 = idxHit[6] ? tgtPages_6 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_35 = idxHit[7] ? tgtPages_7 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_36 = idxHit[8] ? tgtPages_8 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_37 = idxHit[9] ? tgtPages_9 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_38 = idxHit[10] ? tgtPages_10 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_39 = idxHit[11] ? tgtPages_11 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_40 = idxHit[12] ? tgtPages_12 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_41 = idxHit[13] ? tgtPages_13 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_42 = idxHit[14] ? tgtPages_14 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_43 = idxHit[15] ? tgtPages_15 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_44 = idxHit[16] ? tgtPages_16 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_45 = idxHit[17] ? tgtPages_17 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_46 = idxHit[18] ? tgtPages_18 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_47 = idxHit[19] ? tgtPages_19 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_48 = idxHit[20] ? tgtPages_20 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_49 = idxHit[21] ? tgtPages_21 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_50 = idxHit[22] ? tgtPages_22 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_51 = idxHit[23] ? tgtPages_23 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_52 = idxHit[24] ? tgtPages_24 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_53 = idxHit[25] ? tgtPages_25 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_54 = idxHit[26] ? tgtPages_26 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_55 = idxHit[27] ? tgtPages_27 : 3'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_56 = _io_resp_bits_target_T_28 | _io_resp_bits_target_T_29; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_57 = _io_resp_bits_target_T_56 | _io_resp_bits_target_T_30; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_58 = _io_resp_bits_target_T_57 | _io_resp_bits_target_T_31; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_59 = _io_resp_bits_target_T_58 | _io_resp_bits_target_T_32; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_60 = _io_resp_bits_target_T_59 | _io_resp_bits_target_T_33; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_61 = _io_resp_bits_target_T_60 | _io_resp_bits_target_T_34; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_62 = _io_resp_bits_target_T_61 | _io_resp_bits_target_T_35; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_63 = _io_resp_bits_target_T_62 | _io_resp_bits_target_T_36; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_64 = _io_resp_bits_target_T_63 | _io_resp_bits_target_T_37; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_65 = _io_resp_bits_target_T_64 | _io_resp_bits_target_T_38; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_66 = _io_resp_bits_target_T_65 | _io_resp_bits_target_T_39; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_67 = _io_resp_bits_target_T_66 | _io_resp_bits_target_T_40; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_68 = _io_resp_bits_target_T_67 | _io_resp_bits_target_T_41; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_69 = _io_resp_bits_target_T_68 | _io_resp_bits_target_T_42; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_70 = _io_resp_bits_target_T_69 | _io_resp_bits_target_T_43; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_71 = _io_resp_bits_target_T_70 | _io_resp_bits_target_T_44; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_72 = _io_resp_bits_target_T_71 | _io_resp_bits_target_T_45; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_73 = _io_resp_bits_target_T_72 | _io_resp_bits_target_T_46; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_74 = _io_resp_bits_target_T_73 | _io_resp_bits_target_T_47; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_75 = _io_resp_bits_target_T_74 | _io_resp_bits_target_T_48; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_76 = _io_resp_bits_target_T_75 | _io_resp_bits_target_T_49; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_77 = _io_resp_bits_target_T_76 | _io_resp_bits_target_T_50; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_78 = _io_resp_bits_target_T_77 | _io_resp_bits_target_T_51; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_79 = _io_resp_bits_target_T_78 | _io_resp_bits_target_T_52; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_80 = _io_resp_bits_target_T_79 | _io_resp_bits_target_T_53; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_81 = _io_resp_bits_target_T_80 | _io_resp_bits_target_T_54; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_82 = _io_resp_bits_target_T_81 | _io_resp_bits_target_T_55; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_83 = _io_resp_bits_target_T_82 == 3'h1; // @[package.scala 32:86]
  assign _io_resp_bits_target_T_84 = _io_resp_bits_target_T_83 ? pagesMasked_1 : pagesMasked_0; // @[package.scala 32:76]
  assign _io_resp_bits_target_T_85 = _io_resp_bits_target_T_82 == 3'h2; // @[package.scala 32:86]
  assign _io_resp_bits_target_T_86 = _io_resp_bits_target_T_85 ? pagesMasked_2 : _io_resp_bits_target_T_84; // @[package.scala 32:76]
  assign _io_resp_bits_target_T_87 = _io_resp_bits_target_T_82 == 3'h3; // @[package.scala 32:86]
  assign _io_resp_bits_target_T_88 = _io_resp_bits_target_T_87 ? pagesMasked_3 : _io_resp_bits_target_T_86; // @[package.scala 32:76]
  assign _io_resp_bits_target_T_89 = _io_resp_bits_target_T_82 == 3'h4; // @[package.scala 32:86]
  assign _io_resp_bits_target_T_90 = _io_resp_bits_target_T_89 ? pagesMasked_4 : _io_resp_bits_target_T_88; // @[package.scala 32:76]
  assign _io_resp_bits_target_T_91 = _io_resp_bits_target_T_82 == 3'h5; // @[package.scala 32:86]
  assign _io_resp_bits_target_T_92 = _io_resp_bits_target_T_91 ? pagesMasked_5 : _io_resp_bits_target_T_90; // @[package.scala 32:76]
  assign _io_resp_bits_target_T_93 = _io_resp_bits_target_T_82 == 3'h6; // @[package.scala 32:86]
  assign _io_resp_bits_target_T_94 = _io_resp_bits_target_T_93 ? pagesMasked_4 : _io_resp_bits_target_T_92; // @[package.scala 32:76]
  assign _io_resp_bits_target_T_95 = _io_resp_bits_target_T_82 == 3'h7; // @[package.scala 32:86]
  assign io_resp_bits_target_hi = _io_resp_bits_target_T_95 ? pagesMasked_5 : _io_resp_bits_target_T_94; // @[package.scala 32:76]
  assign _io_resp_bits_target_T_124 = idxHit[0] ? tgts_0 : 13'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_125 = idxHit[1] ? tgts_1 : 13'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_126 = idxHit[2] ? tgts_2 : 13'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_127 = idxHit[3] ? tgts_3 : 13'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_128 = idxHit[4] ? tgts_4 : 13'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_129 = idxHit[5] ? tgts_5 : 13'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_130 = idxHit[6] ? tgts_6 : 13'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_131 = idxHit[7] ? tgts_7 : 13'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_132 = idxHit[8] ? tgts_8 : 13'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_133 = idxHit[9] ? tgts_9 : 13'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_134 = idxHit[10] ? tgts_10 : 13'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_135 = idxHit[11] ? tgts_11 : 13'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_136 = idxHit[12] ? tgts_12 : 13'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_137 = idxHit[13] ? tgts_13 : 13'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_138 = idxHit[14] ? tgts_14 : 13'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_139 = idxHit[15] ? tgts_15 : 13'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_140 = idxHit[16] ? tgts_16 : 13'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_141 = idxHit[17] ? tgts_17 : 13'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_142 = idxHit[18] ? tgts_18 : 13'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_143 = idxHit[19] ? tgts_19 : 13'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_144 = idxHit[20] ? tgts_20 : 13'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_145 = idxHit[21] ? tgts_21 : 13'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_146 = idxHit[22] ? tgts_22 : 13'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_147 = idxHit[23] ? tgts_23 : 13'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_148 = idxHit[24] ? tgts_24 : 13'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_149 = idxHit[25] ? tgts_25 : 13'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_150 = idxHit[26] ? tgts_26 : 13'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_151 = idxHit[27] ? tgts_27 : 13'h0; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_152 = _io_resp_bits_target_T_124 | _io_resp_bits_target_T_125; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_153 = _io_resp_bits_target_T_152 | _io_resp_bits_target_T_126; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_154 = _io_resp_bits_target_T_153 | _io_resp_bits_target_T_127; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_155 = _io_resp_bits_target_T_154 | _io_resp_bits_target_T_128; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_156 = _io_resp_bits_target_T_155 | _io_resp_bits_target_T_129; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_157 = _io_resp_bits_target_T_156 | _io_resp_bits_target_T_130; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_158 = _io_resp_bits_target_T_157 | _io_resp_bits_target_T_131; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_159 = _io_resp_bits_target_T_158 | _io_resp_bits_target_T_132; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_160 = _io_resp_bits_target_T_159 | _io_resp_bits_target_T_133; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_161 = _io_resp_bits_target_T_160 | _io_resp_bits_target_T_134; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_162 = _io_resp_bits_target_T_161 | _io_resp_bits_target_T_135; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_163 = _io_resp_bits_target_T_162 | _io_resp_bits_target_T_136; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_164 = _io_resp_bits_target_T_163 | _io_resp_bits_target_T_137; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_165 = _io_resp_bits_target_T_164 | _io_resp_bits_target_T_138; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_166 = _io_resp_bits_target_T_165 | _io_resp_bits_target_T_139; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_167 = _io_resp_bits_target_T_166 | _io_resp_bits_target_T_140; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_168 = _io_resp_bits_target_T_167 | _io_resp_bits_target_T_141; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_169 = _io_resp_bits_target_T_168 | _io_resp_bits_target_T_142; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_170 = _io_resp_bits_target_T_169 | _io_resp_bits_target_T_143; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_171 = _io_resp_bits_target_T_170 | _io_resp_bits_target_T_144; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_172 = _io_resp_bits_target_T_171 | _io_resp_bits_target_T_145; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_173 = _io_resp_bits_target_T_172 | _io_resp_bits_target_T_146; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_174 = _io_resp_bits_target_T_173 | _io_resp_bits_target_T_147; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_175 = _io_resp_bits_target_T_174 | _io_resp_bits_target_T_148; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_176 = _io_resp_bits_target_T_175 | _io_resp_bits_target_T_149; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_177 = _io_resp_bits_target_T_176 | _io_resp_bits_target_T_150; // @[Mux.scala 27:72]
  assign _io_resp_bits_target_T_178 = _io_resp_bits_target_T_177 | _io_resp_bits_target_T_151; // @[Mux.scala 27:72]
  assign io_resp_bits_target_lo = {_io_resp_bits_target_T_178, 1'h0}; // @[BTB.scala 291:88]
  assign _io_resp_bits_target_T_179 = {io_resp_bits_target_hi,io_resp_bits_target_lo}; // @[Cat.scala 30:58]
  assign io_resp_bits_entry_hi = idxHit[27:16]; // @[OneHot.scala 30:18]
  assign io_resp_bits_entry_lo = idxHit[15:0]; // @[OneHot.scala 31:18]
  assign io_resp_bits_entry_hi_1 = |io_resp_bits_entry_hi; // @[OneHot.scala 32:14]
  assign _GEN_436 = {{4'd0}, io_resp_bits_entry_hi}; // @[OneHot.scala 32:28]
  assign _io_resp_bits_entry_T = _GEN_436 | io_resp_bits_entry_lo; // @[OneHot.scala 32:28]
  assign io_resp_bits_entry_hi_2 = _io_resp_bits_entry_T[15:8]; // @[OneHot.scala 30:18]
  assign io_resp_bits_entry_lo_1 = _io_resp_bits_entry_T[7:0]; // @[OneHot.scala 31:18]
  assign io_resp_bits_entry_hi_3 = |io_resp_bits_entry_hi_2; // @[OneHot.scala 32:14]
  assign _io_resp_bits_entry_T_1 = io_resp_bits_entry_hi_2 | io_resp_bits_entry_lo_1; // @[OneHot.scala 32:28]
  assign io_resp_bits_entry_hi_4 = _io_resp_bits_entry_T_1[7:4]; // @[OneHot.scala 30:18]
  assign io_resp_bits_entry_lo_2 = _io_resp_bits_entry_T_1[3:0]; // @[OneHot.scala 31:18]
  assign io_resp_bits_entry_hi_5 = |io_resp_bits_entry_hi_4; // @[OneHot.scala 32:14]
  assign _io_resp_bits_entry_T_2 = io_resp_bits_entry_hi_4 | io_resp_bits_entry_lo_2; // @[OneHot.scala 32:28]
  assign io_resp_bits_entry_hi_6 = _io_resp_bits_entry_T_2[3:2]; // @[OneHot.scala 30:18]
  assign io_resp_bits_entry_lo_3 = _io_resp_bits_entry_T_2[1:0]; // @[OneHot.scala 31:18]
  assign io_resp_bits_entry_hi_7 = |io_resp_bits_entry_hi_6; // @[OneHot.scala 32:14]
  assign _io_resp_bits_entry_T_3 = io_resp_bits_entry_hi_6 | io_resp_bits_entry_lo_3; // @[OneHot.scala 32:28]
  assign io_resp_bits_entry_lo_4 = _io_resp_bits_entry_T_3[1]; // @[CircuitMath.scala 30:8]
  assign io_resp_bits_entry_lo_7 = {io_resp_bits_entry_hi_3,io_resp_bits_entry_hi_5,io_resp_bits_entry_hi_7,io_resp_bits_entry_lo_4}; // @[Cat.scala 30:58]
  assign _io_resp_bits_bridx_T_28 = idxHit[0] & brIdx_0; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_29 = idxHit[1] & brIdx_1; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_30 = idxHit[2] & brIdx_2; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_31 = idxHit[3] & brIdx_3; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_32 = idxHit[4] & brIdx_4; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_33 = idxHit[5] & brIdx_5; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_34 = idxHit[6] & brIdx_6; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_35 = idxHit[7] & brIdx_7; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_36 = idxHit[8] & brIdx_8; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_37 = idxHit[9] & brIdx_9; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_38 = idxHit[10] & brIdx_10; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_39 = idxHit[11] & brIdx_11; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_40 = idxHit[12] & brIdx_12; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_41 = idxHit[13] & brIdx_13; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_42 = idxHit[14] & brIdx_14; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_43 = idxHit[15] & brIdx_15; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_44 = idxHit[16] & brIdx_16; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_45 = idxHit[17] & brIdx_17; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_46 = idxHit[18] & brIdx_18; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_47 = idxHit[19] & brIdx_19; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_48 = idxHit[20] & brIdx_20; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_49 = idxHit[21] & brIdx_21; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_50 = idxHit[22] & brIdx_22; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_51 = idxHit[23] & brIdx_23; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_52 = idxHit[24] & brIdx_24; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_53 = idxHit[25] & brIdx_25; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_54 = idxHit[26] & brIdx_26; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_55 = idxHit[27] & brIdx_27; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_56 = _io_resp_bits_bridx_T_28 | _io_resp_bits_bridx_T_29; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_57 = _io_resp_bits_bridx_T_56 | _io_resp_bits_bridx_T_30; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_58 = _io_resp_bits_bridx_T_57 | _io_resp_bits_bridx_T_31; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_59 = _io_resp_bits_bridx_T_58 | _io_resp_bits_bridx_T_32; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_60 = _io_resp_bits_bridx_T_59 | _io_resp_bits_bridx_T_33; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_61 = _io_resp_bits_bridx_T_60 | _io_resp_bits_bridx_T_34; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_62 = _io_resp_bits_bridx_T_61 | _io_resp_bits_bridx_T_35; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_63 = _io_resp_bits_bridx_T_62 | _io_resp_bits_bridx_T_36; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_64 = _io_resp_bits_bridx_T_63 | _io_resp_bits_bridx_T_37; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_65 = _io_resp_bits_bridx_T_64 | _io_resp_bits_bridx_T_38; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_66 = _io_resp_bits_bridx_T_65 | _io_resp_bits_bridx_T_39; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_67 = _io_resp_bits_bridx_T_66 | _io_resp_bits_bridx_T_40; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_68 = _io_resp_bits_bridx_T_67 | _io_resp_bits_bridx_T_41; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_69 = _io_resp_bits_bridx_T_68 | _io_resp_bits_bridx_T_42; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_70 = _io_resp_bits_bridx_T_69 | _io_resp_bits_bridx_T_43; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_71 = _io_resp_bits_bridx_T_70 | _io_resp_bits_bridx_T_44; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_72 = _io_resp_bits_bridx_T_71 | _io_resp_bits_bridx_T_45; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_73 = _io_resp_bits_bridx_T_72 | _io_resp_bits_bridx_T_46; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_74 = _io_resp_bits_bridx_T_73 | _io_resp_bits_bridx_T_47; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_75 = _io_resp_bits_bridx_T_74 | _io_resp_bits_bridx_T_48; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_76 = _io_resp_bits_bridx_T_75 | _io_resp_bits_bridx_T_49; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_77 = _io_resp_bits_bridx_T_76 | _io_resp_bits_bridx_T_50; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_78 = _io_resp_bits_bridx_T_77 | _io_resp_bits_bridx_T_51; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_79 = _io_resp_bits_bridx_T_78 | _io_resp_bits_bridx_T_52; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_80 = _io_resp_bits_bridx_T_79 | _io_resp_bits_bridx_T_53; // @[Mux.scala 27:72]
  assign _io_resp_bits_bridx_T_81 = _io_resp_bits_bridx_T_80 | _io_resp_bits_bridx_T_54; // @[Mux.scala 27:72]
  assign leftOne = idxHit[0]; // @[Misc.scala 180:37]
  assign leftOne_1 = idxHit[1]; // @[Misc.scala 180:37]
  assign rightOne = idxHit[2]; // @[Misc.scala 181:39]
  assign rightOne_1 = leftOne_1 | rightOne; // @[Misc.scala 182:16]
  assign rightTwo = leftOne_1 & rightOne; // @[Misc.scala 182:61]
  assign leftOne_2 = leftOne | rightOne_1; // @[Misc.scala 182:16]
  assign _T_29 = leftOne & rightOne_1; // @[Misc.scala 182:61]
  assign leftTwo = rightTwo | _T_29; // @[Misc.scala 182:49]
  assign leftOne_3 = idxHit[3]; // @[Misc.scala 180:37]
  assign rightOne_2 = idxHit[4]; // @[Misc.scala 181:39]
  assign leftOne_4 = leftOne_3 | rightOne_2; // @[Misc.scala 182:16]
  assign leftTwo_1 = leftOne_3 & rightOne_2; // @[Misc.scala 182:61]
  assign leftOne_5 = idxHit[5]; // @[Misc.scala 180:37]
  assign rightOne_3 = idxHit[6]; // @[Misc.scala 181:39]
  assign rightOne_4 = leftOne_5 | rightOne_3; // @[Misc.scala 182:16]
  assign rightTwo_1 = leftOne_5 & rightOne_3; // @[Misc.scala 182:61]
  assign rightOne_5 = leftOne_4 | rightOne_4; // @[Misc.scala 182:16]
  assign _T_41 = leftTwo_1 | rightTwo_1; // @[Misc.scala 182:37]
  assign _T_42 = leftOne_4 & rightOne_4; // @[Misc.scala 182:61]
  assign rightTwo_2 = _T_41 | _T_42; // @[Misc.scala 182:49]
  assign leftOne_6 = leftOne_2 | rightOne_5; // @[Misc.scala 182:16]
  assign _T_43 = leftTwo | rightTwo_2; // @[Misc.scala 182:37]
  assign _T_44 = leftOne_2 & rightOne_5; // @[Misc.scala 182:61]
  assign leftTwo_2 = _T_43 | _T_44; // @[Misc.scala 182:49]
  assign leftOne_7 = idxHit[7]; // @[Misc.scala 180:37]
  assign leftOne_8 = idxHit[8]; // @[Misc.scala 180:37]
  assign rightOne_6 = idxHit[9]; // @[Misc.scala 181:39]
  assign rightOne_7 = leftOne_8 | rightOne_6; // @[Misc.scala 182:16]
  assign rightTwo_3 = leftOne_8 & rightOne_6; // @[Misc.scala 182:61]
  assign leftOne_9 = leftOne_7 | rightOne_7; // @[Misc.scala 182:16]
  assign _T_54 = leftOne_7 & rightOne_7; // @[Misc.scala 182:61]
  assign leftTwo_3 = rightTwo_3 | _T_54; // @[Misc.scala 182:49]
  assign leftOne_10 = idxHit[10]; // @[Misc.scala 180:37]
  assign rightOne_8 = idxHit[11]; // @[Misc.scala 181:39]
  assign leftOne_11 = leftOne_10 | rightOne_8; // @[Misc.scala 182:16]
  assign leftTwo_4 = leftOne_10 & rightOne_8; // @[Misc.scala 182:61]
  assign leftOne_12 = idxHit[12]; // @[Misc.scala 180:37]
  assign rightOne_9 = idxHit[13]; // @[Misc.scala 181:39]
  assign rightOne_10 = leftOne_12 | rightOne_9; // @[Misc.scala 182:16]
  assign rightTwo_4 = leftOne_12 & rightOne_9; // @[Misc.scala 182:61]
  assign rightOne_11 = leftOne_11 | rightOne_10; // @[Misc.scala 182:16]
  assign _T_66 = leftTwo_4 | rightTwo_4; // @[Misc.scala 182:37]
  assign _T_67 = leftOne_11 & rightOne_10; // @[Misc.scala 182:61]
  assign rightTwo_5 = _T_66 | _T_67; // @[Misc.scala 182:49]
  assign rightOne_12 = leftOne_9 | rightOne_11; // @[Misc.scala 182:16]
  assign _T_68 = leftTwo_3 | rightTwo_5; // @[Misc.scala 182:37]
  assign _T_69 = leftOne_9 & rightOne_11; // @[Misc.scala 182:61]
  assign rightTwo_6 = _T_68 | _T_69; // @[Misc.scala 182:49]
  assign leftOne_13 = leftOne_6 | rightOne_12; // @[Misc.scala 182:16]
  assign _T_70 = leftTwo_2 | rightTwo_6; // @[Misc.scala 182:37]
  assign _T_71 = leftOne_6 & rightOne_12; // @[Misc.scala 182:61]
  assign leftTwo_5 = _T_70 | _T_71; // @[Misc.scala 182:49]
  assign leftOne_14 = idxHit[14]; // @[Misc.scala 180:37]
  assign leftOne_15 = idxHit[15]; // @[Misc.scala 180:37]
  assign rightOne_13 = idxHit[16]; // @[Misc.scala 181:39]
  assign rightOne_14 = leftOne_15 | rightOne_13; // @[Misc.scala 182:16]
  assign rightTwo_7 = leftOne_15 & rightOne_13; // @[Misc.scala 182:61]
  assign leftOne_16 = leftOne_14 | rightOne_14; // @[Misc.scala 182:16]
  assign _T_82 = leftOne_14 & rightOne_14; // @[Misc.scala 182:61]
  assign leftTwo_6 = rightTwo_7 | _T_82; // @[Misc.scala 182:49]
  assign leftOne_17 = idxHit[17]; // @[Misc.scala 180:37]
  assign rightOne_15 = idxHit[18]; // @[Misc.scala 181:39]
  assign leftOne_18 = leftOne_17 | rightOne_15; // @[Misc.scala 182:16]
  assign leftTwo_7 = leftOne_17 & rightOne_15; // @[Misc.scala 182:61]
  assign leftOne_19 = idxHit[19]; // @[Misc.scala 180:37]
  assign rightOne_16 = idxHit[20]; // @[Misc.scala 181:39]
  assign rightOne_17 = leftOne_19 | rightOne_16; // @[Misc.scala 182:16]
  assign rightTwo_8 = leftOne_19 & rightOne_16; // @[Misc.scala 182:61]
  assign rightOne_18 = leftOne_18 | rightOne_17; // @[Misc.scala 182:16]
  assign _T_94 = leftTwo_7 | rightTwo_8; // @[Misc.scala 182:37]
  assign _T_95 = leftOne_18 & rightOne_17; // @[Misc.scala 182:61]
  assign rightTwo_9 = _T_94 | _T_95; // @[Misc.scala 182:49]
  assign leftOne_20 = leftOne_16 | rightOne_18; // @[Misc.scala 182:16]
  assign _T_96 = leftTwo_6 | rightTwo_9; // @[Misc.scala 182:37]
  assign _T_97 = leftOne_16 & rightOne_18; // @[Misc.scala 182:61]
  assign leftTwo_8 = _T_96 | _T_97; // @[Misc.scala 182:49]
  assign leftOne_21 = idxHit[21]; // @[Misc.scala 180:37]
  assign leftOne_22 = idxHit[22]; // @[Misc.scala 180:37]
  assign rightOne_19 = idxHit[23]; // @[Misc.scala 181:39]
  assign rightOne_20 = leftOne_22 | rightOne_19; // @[Misc.scala 182:16]
  assign rightTwo_10 = leftOne_22 & rightOne_19; // @[Misc.scala 182:61]
  assign leftOne_23 = leftOne_21 | rightOne_20; // @[Misc.scala 182:16]
  assign _T_107 = leftOne_21 & rightOne_20; // @[Misc.scala 182:61]
  assign leftTwo_9 = rightTwo_10 | _T_107; // @[Misc.scala 182:49]
  assign leftOne_24 = idxHit[24]; // @[Misc.scala 180:37]
  assign rightOne_21 = idxHit[25]; // @[Misc.scala 181:39]
  assign leftOne_25 = leftOne_24 | rightOne_21; // @[Misc.scala 182:16]
  assign leftTwo_10 = leftOne_24 & rightOne_21; // @[Misc.scala 182:61]
  assign leftOne_26 = idxHit[26]; // @[Misc.scala 180:37]
  assign rightOne_22 = idxHit[27]; // @[Misc.scala 181:39]
  assign rightOne_23 = leftOne_26 | rightOne_22; // @[Misc.scala 182:16]
  assign rightTwo_11 = leftOne_26 & rightOne_22; // @[Misc.scala 182:61]
  assign rightOne_24 = leftOne_25 | rightOne_23; // @[Misc.scala 182:16]
  assign _T_119 = leftTwo_10 | rightTwo_11; // @[Misc.scala 182:37]
  assign _T_120 = leftOne_25 & rightOne_23; // @[Misc.scala 182:61]
  assign rightTwo_12 = _T_119 | _T_120; // @[Misc.scala 182:49]
  assign rightOne_25 = leftOne_23 | rightOne_24; // @[Misc.scala 182:16]
  assign _T_121 = leftTwo_9 | rightTwo_12; // @[Misc.scala 182:37]
  assign _T_122 = leftOne_23 & rightOne_24; // @[Misc.scala 182:61]
  assign rightTwo_13 = _T_121 | _T_122; // @[Misc.scala 182:49]
  assign rightOne_26 = leftOne_20 | rightOne_25; // @[Misc.scala 182:16]
  assign _T_123 = leftTwo_8 | rightTwo_13; // @[Misc.scala 182:37]
  assign _T_124 = leftOne_20 & rightOne_25; // @[Misc.scala 182:61]
  assign rightTwo_14 = _T_123 | _T_124; // @[Misc.scala 182:49]
  assign _T_126 = leftTwo_5 | rightTwo_14; // @[Misc.scala 182:37]
  assign _T_127 = leftOne_13 & rightOne_26; // @[Misc.scala 182:61]
  assign _T_128 = _T_126 | _T_127; // @[Misc.scala 182:49]
  assign _isValid_T_5 = isValid & ~idxHit; // @[BTB.scala 299:24]
  assign _GEN_374 = _T_128 ? {{4'd0}, _isValid_T_5} : _GEN_338; // @[BTB.scala 298:37]
  assign _GEN_375 = io_flush ? 32'h0 : _GEN_374; // @[BTB.scala 301:19]
  assign resetting = ~reset_waddr[9]; // @[BTB.scala 122:27]
  assign _reset_waddr_T_1 = reset_waddr + 10'h1; // @[BTB.scala 126:49]
  assign waddr_hi_13 = io_bht_update_bits_pc[38:2]; // @[BTB.scala 87:21]
  assign _GEN_437 = {{7'd0}, waddr_hi_13[10:9]}; // @[BTB.scala 88:42]
  assign _waddr_T_30 = waddr_hi_13[8:0] ^ _GEN_437; // @[BTB.scala 88:42]
  assign _waddr_T_31 = 8'hdd * io_bht_update_bits_prediction_history; // @[BTB.scala 84:12]
  assign _waddr_T_33 = {_waddr_T_31[7:5], 6'h0}; // @[BTB.scala 90:44]
  assign _waddr_T_34 = _waddr_T_30 ^ _waddr_T_33; // @[BTB.scala 90:20]
  assign _GEN_383 = resetting ? reset_waddr : {{1'd0}, _waddr_T_34}; // @[BTB.scala 100:23]
  assign _GEN_388 = io_bht_update_bits_branch ? _GEN_383 : reset_waddr; // @[BTB.scala 313:40]
  assign waddr_1 = io_bht_update_valid ? _GEN_388 : reset_waddr; // @[BTB.scala 312:32]
  assign _GEN_387 = io_bht_update_bits_branch | resetting; // @[BTB.scala 313:40]
  assign _GEN_384 = ~resetting & io_bht_update_bits_taken; // @[BTB.scala 100:23]
  assign _GEN_389 = io_bht_update_bits_branch & _GEN_384; // @[BTB.scala 313:40]
  assign isBranch_lo_lo_lo_lo = cfiType_0 == 2'h0; // @[BTB.scala 307:44]
  assign isBranch_lo_lo_lo_hi_lo = cfiType_1 == 2'h0; // @[BTB.scala 307:44]
  assign isBranch_lo_lo_lo_hi_hi = cfiType_2 == 2'h0; // @[BTB.scala 307:44]
  assign isBranch_lo_lo_hi_lo_lo = cfiType_3 == 2'h0; // @[BTB.scala 307:44]
  assign isBranch_lo_lo_hi_lo_hi = cfiType_4 == 2'h0; // @[BTB.scala 307:44]
  assign isBranch_lo_lo_hi_hi_lo = cfiType_5 == 2'h0; // @[BTB.scala 307:44]
  assign isBranch_lo_lo_hi_hi_hi = cfiType_6 == 2'h0; // @[BTB.scala 307:44]
  assign isBranch_lo_hi_lo_lo = cfiType_7 == 2'h0; // @[BTB.scala 307:44]
  assign isBranch_lo_hi_lo_hi_lo = cfiType_8 == 2'h0; // @[BTB.scala 307:44]
  assign isBranch_lo_hi_lo_hi_hi = cfiType_9 == 2'h0; // @[BTB.scala 307:44]
  assign isBranch_lo_hi_hi_lo_lo = cfiType_10 == 2'h0; // @[BTB.scala 307:44]
  assign isBranch_lo_hi_hi_lo_hi = cfiType_11 == 2'h0; // @[BTB.scala 307:44]
  assign isBranch_lo_hi_hi_hi_lo = cfiType_12 == 2'h0; // @[BTB.scala 307:44]
  assign isBranch_lo_hi_hi_hi_hi = cfiType_13 == 2'h0; // @[BTB.scala 307:44]
  assign isBranch_hi_lo_lo_lo = cfiType_14 == 2'h0; // @[BTB.scala 307:44]
  assign isBranch_hi_lo_lo_hi_lo = cfiType_15 == 2'h0; // @[BTB.scala 307:44]
  assign isBranch_hi_lo_lo_hi_hi = cfiType_16 == 2'h0; // @[BTB.scala 307:44]
  assign isBranch_hi_lo_hi_lo_lo = cfiType_17 == 2'h0; // @[BTB.scala 307:44]
  assign isBranch_hi_lo_hi_lo_hi = cfiType_18 == 2'h0; // @[BTB.scala 307:44]
  assign isBranch_hi_lo_hi_hi_lo = cfiType_19 == 2'h0; // @[BTB.scala 307:44]
  assign isBranch_hi_lo_hi_hi_hi = cfiType_20 == 2'h0; // @[BTB.scala 307:44]
  assign isBranch_hi_hi_lo_lo = cfiType_21 == 2'h0; // @[BTB.scala 307:44]
  assign isBranch_hi_hi_lo_hi_lo = cfiType_22 == 2'h0; // @[BTB.scala 307:44]
  assign isBranch_hi_hi_lo_hi_hi = cfiType_23 == 2'h0; // @[BTB.scala 307:44]
  assign isBranch_hi_hi_hi_lo_lo = cfiType_24 == 2'h0; // @[BTB.scala 307:44]
  assign isBranch_hi_hi_hi_lo_hi = cfiType_25 == 2'h0; // @[BTB.scala 307:44]
  assign isBranch_hi_hi_hi_hi_lo = cfiType_26 == 2'h0; // @[BTB.scala 307:44]
  assign isBranch_hi_hi_hi_hi_hi = cfiType_27 == 2'h0; // @[BTB.scala 307:44]
  assign isBranch_lo_lo = {isBranch_lo_lo_hi_hi_hi,isBranch_lo_lo_hi_hi_lo,isBranch_lo_lo_hi_lo_hi,isBranch_lo_lo_hi_lo_lo,isBranch_lo_lo_lo_hi_hi,isBranch_lo_lo_lo_hi_lo,isBranch_lo_lo_lo_lo}; // @[Cat.scala 30:58]
  assign isBranch_lo = {isBranch_lo_hi_hi_hi_hi,isBranch_lo_hi_hi_hi_lo,isBranch_lo_hi_hi_lo_hi,isBranch_lo_hi_hi_lo_lo,isBranch_lo_hi_lo_hi_hi,isBranch_lo_hi_lo_hi_lo,isBranch_lo_hi_lo_lo,isBranch_lo_lo}; // @[Cat.scala 30:58]
  assign isBranch_hi_lo = {isBranch_hi_lo_hi_hi_hi,isBranch_hi_lo_hi_hi_lo,isBranch_hi_lo_hi_lo_hi,isBranch_hi_lo_hi_lo_lo,isBranch_hi_lo_lo_hi_hi,isBranch_hi_lo_lo_hi_lo,isBranch_hi_lo_lo_lo}; // @[Cat.scala 30:58]
  assign _isBranch_T = {isBranch_hi_hi_hi_hi_hi,isBranch_hi_hi_hi_hi_lo,isBranch_hi_hi_hi_lo_hi,isBranch_hi_hi_hi_lo_lo,isBranch_hi_hi_lo_hi_hi,isBranch_hi_hi_lo_hi_lo,isBranch_hi_hi_lo_lo,isBranch_hi_lo,isBranch_lo}; // @[Cat.scala 30:58]
  assign _isBranch_T_1 = idxHit & _isBranch_T; // @[BTB.scala 307:28]
  assign isBranch = |_isBranch_T_1; // @[BTB.scala 307:72]
  assign res_res_value_hi = io_req_bits_addr[38:2]; // @[BTB.scala 87:21]
  assign _GEN_438 = {{7'd0}, res_res_value_hi[10:9]}; // @[BTB.scala 88:42]
  assign _res_res_value_T_3 = res_res_value_hi[8:0] ^ _GEN_438; // @[BTB.scala 88:42]
  assign _res_res_value_T_4 = 8'hdd * history; // @[BTB.scala 84:12]
  assign _res_res_value_T_6 = {_res_res_value_T_4[7:5], 6'h0}; // @[BTB.scala 90:44]
  assign res_value = resetting ? 1'h0 : table__res_res_value_MPORT_data; // @[BTB.scala 94:21]
  assign history_lo = history[7:1]; // @[BTB.scala 115:35]
  assign _history_T = {io_bht_advance_bits_bht_value,history_lo}; // @[Cat.scala 30:58]
  assign history_lo_1 = io_bht_update_bits_prediction_history[7:1]; // @[BTB.scala 112:37]
  assign _history_T_1 = {io_bht_update_bits_taken,history_lo_1}; // @[Cat.scala 30:58]
  assign _T_134 = ~res_value & isBranch; // @[BTB.scala 322:22]
  assign doPeek_lo_lo_lo_lo = cfiType_0 == 2'h3; // @[BTB.scala 328:42]
  assign doPeek_lo_lo_lo_hi_lo = cfiType_1 == 2'h3; // @[BTB.scala 328:42]
  assign doPeek_lo_lo_lo_hi_hi = cfiType_2 == 2'h3; // @[BTB.scala 328:42]
  assign doPeek_lo_lo_hi_lo_lo = cfiType_3 == 2'h3; // @[BTB.scala 328:42]
  assign doPeek_lo_lo_hi_lo_hi = cfiType_4 == 2'h3; // @[BTB.scala 328:42]
  assign doPeek_lo_lo_hi_hi_lo = cfiType_5 == 2'h3; // @[BTB.scala 328:42]
  assign doPeek_lo_lo_hi_hi_hi = cfiType_6 == 2'h3; // @[BTB.scala 328:42]
  assign doPeek_lo_hi_lo_lo = cfiType_7 == 2'h3; // @[BTB.scala 328:42]
  assign doPeek_lo_hi_lo_hi_lo = cfiType_8 == 2'h3; // @[BTB.scala 328:42]
  assign doPeek_lo_hi_lo_hi_hi = cfiType_9 == 2'h3; // @[BTB.scala 328:42]
  assign doPeek_lo_hi_hi_lo_lo = cfiType_10 == 2'h3; // @[BTB.scala 328:42]
  assign doPeek_lo_hi_hi_lo_hi = cfiType_11 == 2'h3; // @[BTB.scala 328:42]
  assign doPeek_lo_hi_hi_hi_lo = cfiType_12 == 2'h3; // @[BTB.scala 328:42]
  assign doPeek_lo_hi_hi_hi_hi = cfiType_13 == 2'h3; // @[BTB.scala 328:42]
  assign doPeek_hi_lo_lo_lo = cfiType_14 == 2'h3; // @[BTB.scala 328:42]
  assign doPeek_hi_lo_lo_hi_lo = cfiType_15 == 2'h3; // @[BTB.scala 328:42]
  assign doPeek_hi_lo_lo_hi_hi = cfiType_16 == 2'h3; // @[BTB.scala 328:42]
  assign doPeek_hi_lo_hi_lo_lo = cfiType_17 == 2'h3; // @[BTB.scala 328:42]
  assign doPeek_hi_lo_hi_lo_hi = cfiType_18 == 2'h3; // @[BTB.scala 328:42]
  assign doPeek_hi_lo_hi_hi_lo = cfiType_19 == 2'h3; // @[BTB.scala 328:42]
  assign doPeek_hi_lo_hi_hi_hi = cfiType_20 == 2'h3; // @[BTB.scala 328:42]
  assign doPeek_hi_hi_lo_lo = cfiType_21 == 2'h3; // @[BTB.scala 328:42]
  assign doPeek_hi_hi_lo_hi_lo = cfiType_22 == 2'h3; // @[BTB.scala 328:42]
  assign doPeek_hi_hi_lo_hi_hi = cfiType_23 == 2'h3; // @[BTB.scala 328:42]
  assign doPeek_hi_hi_hi_lo_lo = cfiType_24 == 2'h3; // @[BTB.scala 328:42]
  assign doPeek_hi_hi_hi_lo_hi = cfiType_25 == 2'h3; // @[BTB.scala 328:42]
  assign doPeek_hi_hi_hi_hi_lo = cfiType_26 == 2'h3; // @[BTB.scala 328:42]
  assign doPeek_hi_hi_hi_hi_hi = cfiType_27 == 2'h3; // @[BTB.scala 328:42]
  assign doPeek_lo_lo = {doPeek_lo_lo_hi_hi_hi,doPeek_lo_lo_hi_hi_lo,doPeek_lo_lo_hi_lo_hi,doPeek_lo_lo_hi_lo_lo,doPeek_lo_lo_lo_hi_hi,doPeek_lo_lo_lo_hi_lo,doPeek_lo_lo_lo_lo}; // @[Cat.scala 30:58]
  assign doPeek_lo = {doPeek_lo_hi_hi_hi_hi,doPeek_lo_hi_hi_hi_lo,doPeek_lo_hi_hi_lo_hi,doPeek_lo_hi_hi_lo_lo,doPeek_lo_hi_lo_hi_hi,doPeek_lo_hi_lo_hi_lo,doPeek_lo_hi_lo_lo,doPeek_lo_lo}; // @[Cat.scala 30:58]
  assign doPeek_hi_lo = {doPeek_hi_lo_hi_hi_hi,doPeek_hi_lo_hi_hi_lo,doPeek_hi_lo_hi_lo_hi,doPeek_hi_lo_hi_lo_lo,doPeek_hi_lo_lo_hi_hi,doPeek_hi_lo_lo_hi_lo,doPeek_hi_lo_lo_lo}; // @[Cat.scala 30:58]
  assign _doPeek_T = {doPeek_hi_hi_hi_hi_hi,doPeek_hi_hi_hi_hi_lo,doPeek_hi_hi_hi_lo_hi,doPeek_hi_hi_hi_lo_lo,doPeek_hi_hi_lo_hi_hi,doPeek_hi_hi_lo_hi_lo,doPeek_hi_hi_lo_lo,doPeek_hi_lo,doPeek_lo}; // @[Cat.scala 30:58]
  assign _doPeek_T_1 = idxHit & _doPeek_T; // @[BTB.scala 328:26]
  assign doPeek = |_doPeek_T_1; // @[BTB.scala 328:67]
  assign _io_ras_head_valid_T = count == 3'h0; // @[BTB.scala 56:29]
  assign _GEN_397 = 3'h1 == pos ? stack_1 : stack_0; // @[BTB.scala 330:22]
  assign _GEN_398 = 3'h2 == pos ? stack_2 : _GEN_397; // @[BTB.scala 330:22]
  assign _GEN_399 = 3'h3 == pos ? stack_3 : _GEN_398; // @[BTB.scala 330:22]
  assign _GEN_400 = 3'h4 == pos ? stack_4 : _GEN_399; // @[BTB.scala 330:22]
  assign _GEN_401 = 3'h5 == pos ? stack_5 : _GEN_400; // @[BTB.scala 330:22]
  assign _T_137 = ~_io_ras_head_valid_T & doPeek; // @[BTB.scala 331:24]
  assign _T_138 = io_ras_update_bits_cfiType == 2'h2; // @[BTB.scala 335:40]
  assign _T_139 = count < 3'h6; // @[BTB.scala 45:17]
  assign _count_T_1 = count + 3'h1; // @[BTB.scala 45:42]
  assign _nextPos_T = pos < 3'h5; // @[BTB.scala 46:49]
  assign _nextPos_T_3 = pos + 3'h1; // @[BTB.scala 46:62]
  assign nextPos = _nextPos_T ? _nextPos_T_3 : 3'h0; // @[BTB.scala 46:22]
  assign _T_140 = io_ras_update_bits_cfiType == 2'h3; // @[BTB.scala 337:46]
  assign _count_T_3 = count - 3'h1; // @[BTB.scala 52:20]
  assign _pos_T = pos > 3'h0; // @[BTB.scala 53:42]
  assign _pos_T_3 = pos - 3'h1; // @[BTB.scala 53:50]
  assign io_resp_valid = _io_resp_valid_T_84[0]; // @[BTB.scala 289:17]
  assign io_resp_bits_taken = _T_134 ? 1'h0 : 1'h1; // @[BTB.scala 290:22 BTB.scala 322:56]
  assign io_resp_bits_bridx = _io_resp_bits_bridx_T_81 | _io_resp_bits_bridx_T_55; // @[BTB.scala 293:22]
  assign io_resp_bits_target = _T_137 ? _GEN_401 : _io_resp_bits_target_T_179; // @[BTB.scala 291:23 BTB.scala 332:27]
  assign io_resp_bits_entry = {io_resp_bits_entry_hi_1,io_resp_bits_entry_lo_7}; // @[BTB.scala 292:22]
  assign io_resp_bits_bht_history = history; // @[BTB.scala 323:22]
  assign io_resp_bits_bht_value = resetting ? 1'h0 : table__res_res_value_MPORT_data; // @[BTB.scala 323:22]
  assign io_ras_head_valid = ~_io_ras_head_valid_T; // @[BTB.scala 329:23]
  assign io_ras_head_bits = 3'h5 == pos ? stack_5 : _GEN_400; // @[BTB.scala 330:22]
  assign BTB_cov_read_addr = BTB_state;
  assign BTB_cov_read_data = BTB_cov[BTB_cov_read_addr]; // @[Coverage map for BTB]
  assign BTB_cov_write_data = 1'h1;
  assign BTB_cov_write_addr = BTB_state;
  assign BTB_cov_write_mask = 1'h1;
  assign BTB_cov_write_en = 1'h1;
  assign mux_cond_0 = idxHit[19];
  assign mux_cond_1 = idxHit[20];
  assign mux_cond_2 = idxHit[27];
  assign mux_cond_3 = idxHit[5];
  assign mux_cond_4 = idxHit[6];
  assign mux_cond_5 = idxHit[15];
  assign mux_cond_6 = idxHit[23];
  assign mux_cond_7 = idxHit[1];
  assign mux_cond_8 = idxHit[10];
  assign mux_cond_9 = idxHit[26];
  assign mux_cond_10 = idxHit[13];
  assign mux_cond_11 = idxHit[24];
  assign mux_cond_12 = idxHit[2];
  assign mux_cond_13 = idxHit[12];
  assign mux_cond_14 = idxHit[17];
  assign mux_cond_15 = idxHit[0];
  assign mux_cond_16 = idxHit[4];
  assign mux_cond_17 = idxHit[22];
  assign mux_cond_18 = idxHit[3];
  assign mux_cond_19 = idxHit[18];
  assign mux_cond_20 = idxHit[11];
  assign mux_cond_21 = idxHit[8];
  assign mux_cond_22 = idxHit[21];
  assign mux_cond_23 = idxHit[25];
  assign mux_cond_24 = _T_128;
  assign mux_cond_25 = idxHit[7];
  assign mux_cond_26 = idxHit[14];
  assign mux_cond_27 = idxHit[16];
  assign mux_cond_28 = idxHit[9];
  assign nextPageRepl_shl = {nextPageRepl, 7'h0};
  assign nextPageRepl_pad = {10'h0,nextPageRepl_shl};
  assign r_respPipe_bits_taken_shl = {r_respPipe_bits_taken, 3'h0};
  assign r_respPipe_bits_taken_pad = {16'h0,r_respPipe_bits_taken_shl};
  assign r_btb_updatePipe_valid_shl = {r_btb_updatePipe_valid, 16'h0};
  assign r_btb_updatePipe_valid_pad = {3'h0,r_btb_updatePipe_valid_shl};
  assign count_shl = {count, 12'h0};
  assign count_pad = {5'h0,count_shl};
  assign r_respPipe_valid_shl = {r_respPipe_valid, 13'h0};
  assign r_respPipe_valid_pad = {6'h0,r_respPipe_valid_shl};
  assign pos_shl = {pos, 1'h0};
  assign pos_pad = {16'h0,pos_shl};
  assign pageValid_shl = {pageValid, 8'h0};
  assign pageValid_pad = {6'h0,pageValid_shl};
  assign r_btb_updatePipe_bits_isValid_shl = {r_btb_updatePipe_bits_isValid, 17'h0};
  assign r_btb_updatePipe_bits_isValid_pad = {2'h0,r_btb_updatePipe_bits_isValid_shl};
  assign mux_cond_0_shl = {mux_cond_0, 14'h0};
  assign mux_cond_0_pad = {5'h0,mux_cond_0_shl};
  assign mux_cond_1_shl = {mux_cond_1, 17'h0};
  assign mux_cond_1_pad = {2'h0,mux_cond_1_shl};
  assign mux_cond_2_shl = {mux_cond_2, 3'h0};
  assign mux_cond_2_pad = {16'h0,mux_cond_2_shl};
  assign mux_cond_3_shl = {mux_cond_3, 17'h0};
  assign mux_cond_3_pad = {2'h0,mux_cond_3_shl};
  assign mux_cond_4_shl = {mux_cond_4, 13'h0};
  assign mux_cond_4_pad = {6'h0,mux_cond_4_shl};
  assign mux_cond_5_shl = {mux_cond_5, 3'h0};
  assign mux_cond_5_pad = {16'h0,mux_cond_5_shl};
  assign mux_cond_6_shl = {mux_cond_6, 1'h0};
  assign mux_cond_6_pad = {18'h0,mux_cond_6_shl};
  assign mux_cond_7_shl = {mux_cond_7, 13'h0};
  assign mux_cond_7_pad = {6'h0,mux_cond_7_shl};
  assign mux_cond_8_shl = {mux_cond_8, 16'h0};
  assign mux_cond_8_pad = {3'h0,mux_cond_8_shl};
  assign mux_cond_9_shl = {mux_cond_9, 3'h0};
  assign mux_cond_9_pad = {16'h0,mux_cond_9_shl};
  assign mux_cond_10_shl = {mux_cond_10, 9'h0};
  assign mux_cond_10_pad = {10'h0,mux_cond_10_shl};
  assign mux_cond_11_shl = {mux_cond_11, 3'h0};
  assign mux_cond_11_pad = {16'h0,mux_cond_11_shl};
  assign mux_cond_12_shl = {mux_cond_12, 17'h0};
  assign mux_cond_12_pad = {2'h0,mux_cond_12_shl};
  assign mux_cond_13_shl = {mux_cond_13, 8'h0};
  assign mux_cond_13_pad = {11'h0,mux_cond_13_shl};
  assign mux_cond_14_shl = {mux_cond_14, 4'h0};
  assign mux_cond_14_pad = {15'h0,mux_cond_14_shl};
  assign mux_cond_15_shl = {mux_cond_15, 11'h0};
  assign mux_cond_15_pad = {8'h0,mux_cond_15_shl};
  assign mux_cond_16_shl = {mux_cond_16, 12'h0};
  assign mux_cond_16_pad = {7'h0,mux_cond_16_shl};
  assign mux_cond_17_shl = {mux_cond_17, 5'h0};
  assign mux_cond_17_pad = {14'h0,mux_cond_17_shl};
  assign mux_cond_18_shl = mux_cond_18;
  assign mux_cond_18_pad = {19'h0,mux_cond_18_shl};
  assign mux_cond_19_shl = {mux_cond_19, 1'h0};
  assign mux_cond_19_pad = {18'h0,mux_cond_19_shl};
  assign mux_cond_20_shl = {mux_cond_20, 2'h0};
  assign mux_cond_20_pad = {17'h0,mux_cond_20_shl};
  assign mux_cond_21_shl = {mux_cond_21, 5'h0};
  assign mux_cond_21_pad = {14'h0,mux_cond_21_shl};
  assign mux_cond_22_shl = {mux_cond_22, 16'h0};
  assign mux_cond_22_pad = {3'h0,mux_cond_22_shl};
  assign mux_cond_23_shl = {mux_cond_23, 13'h0};
  assign mux_cond_23_pad = {6'h0,mux_cond_23_shl};
  assign mux_cond_24_shl = {mux_cond_24, 19'h0};
  assign mux_cond_24_pad = mux_cond_24_shl;
  assign mux_cond_25_shl = {mux_cond_25, 14'h0};
  assign mux_cond_25_pad = {5'h0,mux_cond_25_shl};
  assign mux_cond_26_shl = {mux_cond_26, 8'h0};
  assign mux_cond_26_pad = {11'h0,mux_cond_26_shl};
  assign mux_cond_27_shl = {mux_cond_27, 18'h0};
  assign mux_cond_27_pad = {1'h0,mux_cond_27_shl};
  assign mux_cond_28_shl = {mux_cond_28, 5'h0};
  assign mux_cond_28_pad = {14'h0,mux_cond_28_shl};
  assign cfiType_17_shl = {cfiType_17, 11'h0};
  assign cfiType_17_pad = {7'h0,cfiType_17_shl};
  assign cfiType_22_shl = {cfiType_22, 11'h0};
  assign cfiType_22_pad = {7'h0,cfiType_22_shl};
  assign cfiType_21_shl = {cfiType_21, 11'h0};
  assign cfiType_21_pad = {7'h0,cfiType_21_shl};
  assign tgtPages_4_shl = {tgtPages_4, 15'h0};
  assign tgtPages_4_pad = {2'h0,tgtPages_4_shl};
  assign tgtPages_6_shl = {tgtPages_6, 15'h0};
  assign tgtPages_6_pad = {2'h0,tgtPages_6_shl};
  assign tgtPages_11_shl = {tgtPages_11, 15'h0};
  assign tgtPages_11_pad = {2'h0,tgtPages_11_shl};
  assign tgtPages_7_shl = {tgtPages_7, 15'h0};
  assign tgtPages_7_pad = {2'h0,tgtPages_7_shl};
  assign tgtPages_20_shl = {tgtPages_20, 15'h0};
  assign tgtPages_20_pad = {2'h0,tgtPages_20_shl};
  assign cfiType_3_shl = {cfiType_3, 11'h0};
  assign cfiType_3_pad = {7'h0,cfiType_3_shl};
  assign tgtPages_16_shl = {tgtPages_16, 15'h0};
  assign tgtPages_16_pad = {2'h0,tgtPages_16_shl};
  assign cfiType_24_shl = {cfiType_24, 11'h0};
  assign cfiType_24_pad = {7'h0,cfiType_24_shl};
  assign tgtPages_17_shl = {tgtPages_17, 15'h0};
  assign tgtPages_17_pad = {2'h0,tgtPages_17_shl};
  assign cfiType_6_shl = {cfiType_6, 11'h0};
  assign cfiType_6_pad = {7'h0,cfiType_6_shl};
  assign tgtPages_9_shl = {tgtPages_9, 15'h0};
  assign tgtPages_9_pad = {2'h0,tgtPages_9_shl};
  assign tgtPages_2_shl = {tgtPages_2, 15'h0};
  assign tgtPages_2_pad = {2'h0,tgtPages_2_shl};
  assign cfiType_10_shl = {cfiType_10, 11'h0};
  assign cfiType_10_pad = {7'h0,cfiType_10_shl};
  assign tgtPages_18_shl = {tgtPages_18, 15'h0};
  assign tgtPages_18_pad = {2'h0,tgtPages_18_shl};
  assign tgtPages_0_shl = {tgtPages_0, 15'h0};
  assign tgtPages_0_pad = {2'h0,tgtPages_0_shl};
  assign tgtPages_25_shl = {tgtPages_25, 15'h0};
  assign tgtPages_25_pad = {2'h0,tgtPages_25_shl};
  assign tgtPages_22_shl = {tgtPages_22, 15'h0};
  assign tgtPages_22_pad = {2'h0,tgtPages_22_shl};
  assign cfiType_5_shl = {cfiType_5, 11'h0};
  assign cfiType_5_pad = {7'h0,cfiType_5_shl};
  assign cfiType_12_shl = {cfiType_12, 11'h0};
  assign cfiType_12_pad = {7'h0,cfiType_12_shl};
  assign cfiType_18_shl = {cfiType_18, 11'h0};
  assign cfiType_18_pad = {7'h0,cfiType_18_shl};
  assign tgtPages_24_shl = {tgtPages_24, 15'h0};
  assign tgtPages_24_pad = {2'h0,tgtPages_24_shl};
  assign tgtPages_26_shl = {tgtPages_26, 15'h0};
  assign tgtPages_26_pad = {2'h0,tgtPages_26_shl};
  assign tgtPages_1_shl = {tgtPages_1, 15'h0};
  assign tgtPages_1_pad = {2'h0,tgtPages_1_shl};
  assign tgtPages_10_shl = {tgtPages_10, 15'h0};
  assign tgtPages_10_pad = {2'h0,tgtPages_10_shl};
  assign cfiType_25_shl = {cfiType_25, 11'h0};
  assign cfiType_25_pad = {7'h0,cfiType_25_shl};
  assign cfiType_16_shl = {cfiType_16, 11'h0};
  assign cfiType_16_pad = {7'h0,cfiType_16_shl};
  assign tgtPages_13_shl = {tgtPages_13, 15'h0};
  assign tgtPages_13_pad = {2'h0,tgtPages_13_shl};
  assign cfiType_19_shl = {cfiType_19, 11'h0};
  assign cfiType_19_pad = {7'h0,cfiType_19_shl};
  assign cfiType_2_shl = {cfiType_2, 11'h0};
  assign cfiType_2_pad = {7'h0,cfiType_2_shl};
  assign cfiType_20_shl = {cfiType_20, 11'h0};
  assign cfiType_20_pad = {7'h0,cfiType_20_shl};
  assign tgtPages_15_shl = {tgtPages_15, 15'h0};
  assign tgtPages_15_pad = {2'h0,tgtPages_15_shl};
  assign tgtPages_8_shl = {tgtPages_8, 15'h0};
  assign tgtPages_8_pad = {2'h0,tgtPages_8_shl};
  assign tgtPages_5_shl = {tgtPages_5, 15'h0};
  assign tgtPages_5_pad = {2'h0,tgtPages_5_shl};
  assign cfiType_0_shl = {cfiType_0, 11'h0};
  assign cfiType_0_pad = {7'h0,cfiType_0_shl};
  assign tgtPages_3_shl = {tgtPages_3, 15'h0};
  assign tgtPages_3_pad = {2'h0,tgtPages_3_shl};
  assign tgtPages_27_shl = {tgtPages_27, 15'h0};
  assign tgtPages_27_pad = {2'h0,tgtPages_27_shl};
  assign cfiType_27_shl = {cfiType_27, 11'h0};
  assign cfiType_27_pad = {7'h0,cfiType_27_shl};
  assign tgtPages_14_shl = {tgtPages_14, 15'h0};
  assign tgtPages_14_pad = {2'h0,tgtPages_14_shl};
  assign cfiType_13_shl = {cfiType_13, 11'h0};
  assign cfiType_13_pad = {7'h0,cfiType_13_shl};
  assign cfiType_23_shl = {cfiType_23, 11'h0};
  assign cfiType_23_pad = {7'h0,cfiType_23_shl};
  assign cfiType_4_shl = {cfiType_4, 11'h0};
  assign cfiType_4_pad = {7'h0,cfiType_4_shl};
  assign cfiType_1_shl = {cfiType_1, 11'h0};
  assign cfiType_1_pad = {7'h0,cfiType_1_shl};
  assign tgtPages_21_shl = {tgtPages_21, 15'h0};
  assign tgtPages_21_pad = {2'h0,tgtPages_21_shl};
  assign cfiType_8_shl = {cfiType_8, 11'h0};
  assign cfiType_8_pad = {7'h0,cfiType_8_shl};
  assign tgtPages_23_shl = {tgtPages_23, 15'h0};
  assign tgtPages_23_pad = {2'h0,tgtPages_23_shl};
  assign tgtPages_19_shl = {tgtPages_19, 15'h0};
  assign tgtPages_19_pad = {2'h0,tgtPages_19_shl};
  assign cfiType_11_shl = {cfiType_11, 11'h0};
  assign cfiType_11_pad = {7'h0,cfiType_11_shl};
  assign tgtPages_12_shl = {tgtPages_12, 15'h0};
  assign tgtPages_12_pad = {2'h0,tgtPages_12_shl};
  assign cfiType_9_shl = {cfiType_9, 11'h0};
  assign cfiType_9_pad = {7'h0,cfiType_9_shl};
  assign cfiType_14_shl = {cfiType_14, 11'h0};
  assign cfiType_14_pad = {7'h0,cfiType_14_shl};
  assign cfiType_7_shl = {cfiType_7, 11'h0};
  assign cfiType_7_pad = {7'h0,cfiType_7_shl};
  assign cfiType_26_shl = {cfiType_26, 11'h0};
  assign cfiType_26_pad = {7'h0,cfiType_26_shl};
  assign cfiType_15_shl = {cfiType_15, 11'h0};
  assign cfiType_15_pad = {7'h0,cfiType_15_shl};
  assign BTB_xor31 = nextPageRepl_pad ^ r_respPipe_bits_taken_pad;
  assign BTB_xor66 = count_pad ^ r_respPipe_valid_pad;
  assign BTB_xor32 = r_btb_updatePipe_valid_pad ^ BTB_xor66;
  assign BTB_xor15 = BTB_xor31 ^ BTB_xor32;
  assign BTB_xor68 = pageValid_pad ^ r_btb_updatePipe_bits_isValid_pad;
  assign BTB_xor33 = pos_pad ^ BTB_xor68;
  assign BTB_xor70 = mux_cond_1_pad ^ mux_cond_2_pad;
  assign BTB_xor34 = mux_cond_0_pad ^ BTB_xor70;
  assign BTB_xor16 = BTB_xor33 ^ BTB_xor34;
  assign BTB_xor7 = BTB_xor15 ^ BTB_xor16;
  assign BTB_xor72 = mux_cond_4_pad ^ mux_cond_5_pad;
  assign BTB_xor35 = mux_cond_3_pad ^ BTB_xor72;
  assign BTB_xor74 = mux_cond_7_pad ^ mux_cond_8_pad;
  assign BTB_xor36 = mux_cond_6_pad ^ BTB_xor74;
  assign BTB_xor17 = BTB_xor35 ^ BTB_xor36;
  assign BTB_xor76 = mux_cond_10_pad ^ mux_cond_11_pad;
  assign BTB_xor37 = mux_cond_9_pad ^ BTB_xor76;
  assign BTB_xor78 = mux_cond_13_pad ^ mux_cond_14_pad;
  assign BTB_xor38 = mux_cond_12_pad ^ BTB_xor78;
  assign BTB_xor18 = BTB_xor37 ^ BTB_xor38;
  assign BTB_xor8 = BTB_xor17 ^ BTB_xor18;
  assign BTB_xor3 = BTB_xor7 ^ BTB_xor8;
  assign BTB_xor39 = mux_cond_15_pad ^ mux_cond_16_pad;
  assign BTB_xor82 = mux_cond_18_pad ^ mux_cond_19_pad;
  assign BTB_xor40 = mux_cond_17_pad ^ BTB_xor82;
  assign BTB_xor19 = BTB_xor39 ^ BTB_xor40;
  assign BTB_xor84 = mux_cond_21_pad ^ mux_cond_22_pad;
  assign BTB_xor41 = mux_cond_20_pad ^ BTB_xor84;
  assign BTB_xor86 = mux_cond_24_pad ^ mux_cond_25_pad;
  assign BTB_xor42 = mux_cond_23_pad ^ BTB_xor86;
  assign BTB_xor20 = BTB_xor41 ^ BTB_xor42;
  assign BTB_xor9 = BTB_xor19 ^ BTB_xor20;
  assign BTB_xor88 = mux_cond_27_pad ^ mux_cond_28_pad;
  assign BTB_xor43 = mux_cond_26_pad ^ BTB_xor88;
  assign BTB_xor90 = cfiType_22_pad ^ cfiType_21_pad;
  assign BTB_xor44 = cfiType_17_pad ^ BTB_xor90;
  assign BTB_xor21 = BTB_xor43 ^ BTB_xor44;
  assign BTB_xor92 = tgtPages_6_pad ^ tgtPages_11_pad;
  assign BTB_xor45 = tgtPages_4_pad ^ BTB_xor92;
  assign BTB_xor94 = tgtPages_20_pad ^ cfiType_3_pad;
  assign BTB_xor46 = tgtPages_7_pad ^ BTB_xor94;
  assign BTB_xor22 = BTB_xor45 ^ BTB_xor46;
  assign BTB_xor10 = BTB_xor21 ^ BTB_xor22;
  assign BTB_xor4 = BTB_xor9 ^ BTB_xor10;
  assign BTB_xor1 = BTB_xor3 ^ BTB_xor4;
  assign BTB_xor47 = tgtPages_16_pad ^ cfiType_24_pad;
  assign BTB_xor98 = cfiType_6_pad ^ tgtPages_9_pad;
  assign BTB_xor48 = tgtPages_17_pad ^ BTB_xor98;
  assign BTB_xor23 = BTB_xor47 ^ BTB_xor48;
  assign BTB_xor100 = cfiType_10_pad ^ tgtPages_18_pad;
  assign BTB_xor49 = tgtPages_2_pad ^ BTB_xor100;
  assign BTB_xor102 = tgtPages_25_pad ^ tgtPages_22_pad;
  assign BTB_xor50 = tgtPages_0_pad ^ BTB_xor102;
  assign BTB_xor24 = BTB_xor49 ^ BTB_xor50;
  assign BTB_xor11 = BTB_xor23 ^ BTB_xor24;
  assign BTB_xor104 = cfiType_12_pad ^ cfiType_18_pad;
  assign BTB_xor51 = cfiType_5_pad ^ BTB_xor104;
  assign BTB_xor106 = tgtPages_26_pad ^ tgtPages_1_pad;
  assign BTB_xor52 = tgtPages_24_pad ^ BTB_xor106;
  assign BTB_xor25 = BTB_xor51 ^ BTB_xor52;
  assign BTB_xor108 = cfiType_25_pad ^ cfiType_16_pad;
  assign BTB_xor53 = tgtPages_10_pad ^ BTB_xor108;
  assign BTB_xor110 = cfiType_19_pad ^ cfiType_2_pad;
  assign BTB_xor54 = tgtPages_13_pad ^ BTB_xor110;
  assign BTB_xor26 = BTB_xor53 ^ BTB_xor54;
  assign BTB_xor12 = BTB_xor25 ^ BTB_xor26;
  assign BTB_xor5 = BTB_xor11 ^ BTB_xor12;
  assign BTB_xor112 = tgtPages_15_pad ^ tgtPages_8_pad;
  assign BTB_xor55 = cfiType_20_pad ^ BTB_xor112;
  assign BTB_xor114 = cfiType_0_pad ^ tgtPages_3_pad;
  assign BTB_xor56 = tgtPages_5_pad ^ BTB_xor114;
  assign BTB_xor27 = BTB_xor55 ^ BTB_xor56;
  assign BTB_xor116 = cfiType_27_pad ^ tgtPages_14_pad;
  assign BTB_xor57 = tgtPages_27_pad ^ BTB_xor116;
  assign BTB_xor118 = cfiType_23_pad ^ cfiType_4_pad;
  assign BTB_xor58 = cfiType_13_pad ^ BTB_xor118;
  assign BTB_xor28 = BTB_xor57 ^ BTB_xor58;
  assign BTB_xor13 = BTB_xor27 ^ BTB_xor28;
  assign BTB_xor120 = tgtPages_21_pad ^ cfiType_8_pad;
  assign BTB_xor59 = cfiType_1_pad ^ BTB_xor120;
  assign BTB_xor122 = tgtPages_19_pad ^ cfiType_11_pad;
  assign BTB_xor60 = tgtPages_23_pad ^ BTB_xor122;
  assign BTB_xor29 = BTB_xor59 ^ BTB_xor60;
  assign BTB_xor124 = cfiType_9_pad ^ cfiType_14_pad;
  assign BTB_xor61 = tgtPages_12_pad ^ BTB_xor124;
  assign BTB_xor126 = cfiType_26_pad ^ cfiType_15_pad;
  assign BTB_xor62 = cfiType_7_pad ^ BTB_xor126;
  assign BTB_xor30 = BTB_xor61 ^ BTB_xor62;
  assign BTB_xor14 = BTB_xor29 ^ BTB_xor30;
  assign BTB_xor6 = BTB_xor13 ^ BTB_xor14;
  assign BTB_xor2 = BTB_xor5 ^ BTB_xor6;
  assign BTB_xor0 = BTB_xor1 ^ BTB_xor2;
  assign io_covSum = BTB_covSum;
  assign metaAssert = 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    table_[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  idxs_0 = _RAND_1[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  idxs_1 = _RAND_2[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  idxs_2 = _RAND_3[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  idxs_3 = _RAND_4[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  idxs_4 = _RAND_5[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  idxs_5 = _RAND_6[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  idxs_6 = _RAND_7[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  idxs_7 = _RAND_8[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  idxs_8 = _RAND_9[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  idxs_9 = _RAND_10[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  idxs_10 = _RAND_11[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  idxs_11 = _RAND_12[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  idxs_12 = _RAND_13[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  idxs_13 = _RAND_14[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  idxs_14 = _RAND_15[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  idxs_15 = _RAND_16[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  idxs_16 = _RAND_17[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  idxs_17 = _RAND_18[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  idxs_18 = _RAND_19[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  idxs_19 = _RAND_20[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  idxs_20 = _RAND_21[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  idxs_21 = _RAND_22[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  idxs_22 = _RAND_23[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  idxs_23 = _RAND_24[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  idxs_24 = _RAND_25[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  idxs_25 = _RAND_26[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  idxs_26 = _RAND_27[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  idxs_27 = _RAND_28[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  idxPages_0 = _RAND_29[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  idxPages_1 = _RAND_30[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  idxPages_2 = _RAND_31[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  idxPages_3 = _RAND_32[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  idxPages_4 = _RAND_33[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  idxPages_5 = _RAND_34[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  idxPages_6 = _RAND_35[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  idxPages_7 = _RAND_36[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  idxPages_8 = _RAND_37[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  idxPages_9 = _RAND_38[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  idxPages_10 = _RAND_39[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  idxPages_11 = _RAND_40[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  idxPages_12 = _RAND_41[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  idxPages_13 = _RAND_42[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  idxPages_14 = _RAND_43[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  idxPages_15 = _RAND_44[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  idxPages_16 = _RAND_45[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  idxPages_17 = _RAND_46[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  idxPages_18 = _RAND_47[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  idxPages_19 = _RAND_48[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  idxPages_20 = _RAND_49[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  idxPages_21 = _RAND_50[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  idxPages_22 = _RAND_51[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  idxPages_23 = _RAND_52[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  idxPages_24 = _RAND_53[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  idxPages_25 = _RAND_54[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  idxPages_26 = _RAND_55[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  idxPages_27 = _RAND_56[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  tgts_0 = _RAND_57[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  tgts_1 = _RAND_58[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  tgts_2 = _RAND_59[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  tgts_3 = _RAND_60[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  tgts_4 = _RAND_61[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  tgts_5 = _RAND_62[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  tgts_6 = _RAND_63[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  tgts_7 = _RAND_64[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  tgts_8 = _RAND_65[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  tgts_9 = _RAND_66[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  tgts_10 = _RAND_67[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  tgts_11 = _RAND_68[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  tgts_12 = _RAND_69[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  tgts_13 = _RAND_70[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  tgts_14 = _RAND_71[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  tgts_15 = _RAND_72[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  tgts_16 = _RAND_73[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  tgts_17 = _RAND_74[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  tgts_18 = _RAND_75[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  tgts_19 = _RAND_76[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  tgts_20 = _RAND_77[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  tgts_21 = _RAND_78[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  tgts_22 = _RAND_79[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  tgts_23 = _RAND_80[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  tgts_24 = _RAND_81[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  tgts_25 = _RAND_82[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  tgts_26 = _RAND_83[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  tgts_27 = _RAND_84[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  tgtPages_0 = _RAND_85[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  tgtPages_1 = _RAND_86[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  tgtPages_2 = _RAND_87[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  tgtPages_3 = _RAND_88[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  tgtPages_4 = _RAND_89[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  tgtPages_5 = _RAND_90[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  tgtPages_6 = _RAND_91[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  tgtPages_7 = _RAND_92[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  tgtPages_8 = _RAND_93[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  tgtPages_9 = _RAND_94[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  tgtPages_10 = _RAND_95[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  tgtPages_11 = _RAND_96[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  tgtPages_12 = _RAND_97[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  tgtPages_13 = _RAND_98[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  tgtPages_14 = _RAND_99[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  tgtPages_15 = _RAND_100[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  tgtPages_16 = _RAND_101[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  tgtPages_17 = _RAND_102[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  tgtPages_18 = _RAND_103[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  tgtPages_19 = _RAND_104[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  tgtPages_20 = _RAND_105[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  tgtPages_21 = _RAND_106[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  tgtPages_22 = _RAND_107[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  tgtPages_23 = _RAND_108[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  tgtPages_24 = _RAND_109[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  tgtPages_25 = _RAND_110[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  tgtPages_26 = _RAND_111[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  tgtPages_27 = _RAND_112[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  pages_0 = _RAND_113[24:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  pages_1 = _RAND_114[24:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  pages_2 = _RAND_115[24:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  pages_3 = _RAND_116[24:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  pages_4 = _RAND_117[24:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  pages_5 = _RAND_118[24:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  pageValid = _RAND_119[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  isValid = _RAND_120[27:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  cfiType_0 = _RAND_121[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  cfiType_1 = _RAND_122[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  cfiType_2 = _RAND_123[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  cfiType_3 = _RAND_124[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  cfiType_4 = _RAND_125[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  cfiType_5 = _RAND_126[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  cfiType_6 = _RAND_127[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  cfiType_7 = _RAND_128[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  cfiType_8 = _RAND_129[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  cfiType_9 = _RAND_130[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  cfiType_10 = _RAND_131[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  cfiType_11 = _RAND_132[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  cfiType_12 = _RAND_133[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  cfiType_13 = _RAND_134[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  cfiType_14 = _RAND_135[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  cfiType_15 = _RAND_136[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  cfiType_16 = _RAND_137[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  cfiType_17 = _RAND_138[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  cfiType_18 = _RAND_139[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  cfiType_19 = _RAND_140[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  cfiType_20 = _RAND_141[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  cfiType_21 = _RAND_142[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  cfiType_22 = _RAND_143[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  cfiType_23 = _RAND_144[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  cfiType_24 = _RAND_145[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  cfiType_25 = _RAND_146[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  cfiType_26 = _RAND_147[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  cfiType_27 = _RAND_148[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  brIdx_0 = _RAND_149[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  brIdx_1 = _RAND_150[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  brIdx_2 = _RAND_151[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  brIdx_3 = _RAND_152[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  brIdx_4 = _RAND_153[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  brIdx_5 = _RAND_154[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  brIdx_6 = _RAND_155[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  brIdx_7 = _RAND_156[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  brIdx_8 = _RAND_157[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  brIdx_9 = _RAND_158[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  brIdx_10 = _RAND_159[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  brIdx_11 = _RAND_160[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  brIdx_12 = _RAND_161[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  brIdx_13 = _RAND_162[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  brIdx_14 = _RAND_163[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  brIdx_15 = _RAND_164[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  brIdx_16 = _RAND_165[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  brIdx_17 = _RAND_166[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  brIdx_18 = _RAND_167[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  brIdx_19 = _RAND_168[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  brIdx_20 = _RAND_169[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  brIdx_21 = _RAND_170[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  brIdx_22 = _RAND_171[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  brIdx_23 = _RAND_172[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  brIdx_24 = _RAND_173[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  brIdx_25 = _RAND_174[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  brIdx_26 = _RAND_175[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  brIdx_27 = _RAND_176[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  r_btb_updatePipe_valid = _RAND_177[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  r_btb_updatePipe_bits_prediction_entry = _RAND_178[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {2{`RANDOM}};
  r_btb_updatePipe_bits_pc = _RAND_179[38:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  r_btb_updatePipe_bits_isValid = _RAND_180[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {2{`RANDOM}};
  r_btb_updatePipe_bits_br_pc = _RAND_181[38:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  r_btb_updatePipe_bits_cfiType = _RAND_182[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  nextPageRepl = _RAND_183[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  state_reg = _RAND_184[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  r_respPipe_valid = _RAND_185[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  r_respPipe_bits_taken = _RAND_186[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  r_respPipe_bits_entry = _RAND_187[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  history = _RAND_188[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  reset_waddr = _RAND_189[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  count = _RAND_190[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  pos = _RAND_191[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {2{`RANDOM}};
  stack_0 = _RAND_192[38:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {2{`RANDOM}};
  stack_1 = _RAND_193[38:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {2{`RANDOM}};
  stack_2 = _RAND_194[38:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {2{`RANDOM}};
  stack_3 = _RAND_195[38:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {2{`RANDOM}};
  stack_4 = _RAND_196[38:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {2{`RANDOM}};
  stack_5 = _RAND_197[38:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  BTB_state = _RAND_198[19:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1048576; initvar = initvar+1)
    BTB_cov[initvar] = _RAND_199[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  BTB_covSum = _RAND_200[29:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(table__MPORT_en & table__MPORT_mask) begin
      table_[table__MPORT_addr] <= table__MPORT_data; // @[BTB.scala 118:26]
    end
    if (metaReset) begin
      idxs_0 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h0 == waddr) begin
        idxs_0 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_1 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h1 == waddr) begin
        idxs_1 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_2 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h2 == waddr) begin
        idxs_2 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_3 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h3 == waddr) begin
        idxs_3 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_4 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h4 == waddr) begin
        idxs_4 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_5 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h5 == waddr) begin
        idxs_5 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_6 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h6 == waddr) begin
        idxs_6 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_7 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h7 == waddr) begin
        idxs_7 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_8 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h8 == waddr) begin
        idxs_8 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_9 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h9 == waddr) begin
        idxs_9 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_10 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'ha == waddr) begin
        idxs_10 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_11 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hb == waddr) begin
        idxs_11 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_12 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hc == waddr) begin
        idxs_12 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_13 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hd == waddr) begin
        idxs_13 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_14 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'he == waddr) begin
        idxs_14 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_15 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hf == waddr) begin
        idxs_15 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_16 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h10 == waddr) begin
        idxs_16 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_17 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h11 == waddr) begin
        idxs_17 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_18 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h12 == waddr) begin
        idxs_18 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_19 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h13 == waddr) begin
        idxs_19 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_20 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h14 == waddr) begin
        idxs_20 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_21 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h15 == waddr) begin
        idxs_21 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_22 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h16 == waddr) begin
        idxs_22 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_23 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h17 == waddr) begin
        idxs_23 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_24 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h18 == waddr) begin
        idxs_24 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_25 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h19 == waddr) begin
        idxs_25 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_26 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h1a == waddr) begin
        idxs_26 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxs_27 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h1b == waddr) begin
        idxs_27 <= r_btb_updatePipe_bits_pc[13:1];
      end
    end
    if (metaReset) begin
      idxPages_0 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h0 == waddr) begin
        idxPages_0 <= _idxPages_T[2:0];
      end
    end
    if (metaReset) begin
      idxPages_1 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h1 == waddr) begin
        idxPages_1 <= _idxPages_T[2:0];
      end
    end
    if (metaReset) begin
      idxPages_2 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h2 == waddr) begin
        idxPages_2 <= _idxPages_T[2:0];
      end
    end
    if (metaReset) begin
      idxPages_3 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h3 == waddr) begin
        idxPages_3 <= _idxPages_T[2:0];
      end
    end
    if (metaReset) begin
      idxPages_4 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h4 == waddr) begin
        idxPages_4 <= _idxPages_T[2:0];
      end
    end
    if (metaReset) begin
      idxPages_5 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h5 == waddr) begin
        idxPages_5 <= _idxPages_T[2:0];
      end
    end
    if (metaReset) begin
      idxPages_6 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h6 == waddr) begin
        idxPages_6 <= _idxPages_T[2:0];
      end
    end
    if (metaReset) begin
      idxPages_7 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h7 == waddr) begin
        idxPages_7 <= _idxPages_T[2:0];
      end
    end
    if (metaReset) begin
      idxPages_8 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h8 == waddr) begin
        idxPages_8 <= _idxPages_T[2:0];
      end
    end
    if (metaReset) begin
      idxPages_9 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h9 == waddr) begin
        idxPages_9 <= _idxPages_T[2:0];
      end
    end
    if (metaReset) begin
      idxPages_10 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'ha == waddr) begin
        idxPages_10 <= _idxPages_T[2:0];
      end
    end
    if (metaReset) begin
      idxPages_11 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hb == waddr) begin
        idxPages_11 <= _idxPages_T[2:0];
      end
    end
    if (metaReset) begin
      idxPages_12 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hc == waddr) begin
        idxPages_12 <= _idxPages_T[2:0];
      end
    end
    if (metaReset) begin
      idxPages_13 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hd == waddr) begin
        idxPages_13 <= _idxPages_T[2:0];
      end
    end
    if (metaReset) begin
      idxPages_14 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'he == waddr) begin
        idxPages_14 <= _idxPages_T[2:0];
      end
    end
    if (metaReset) begin
      idxPages_15 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hf == waddr) begin
        idxPages_15 <= _idxPages_T[2:0];
      end
    end
    if (metaReset) begin
      idxPages_16 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h10 == waddr) begin
        idxPages_16 <= _idxPages_T[2:0];
      end
    end
    if (metaReset) begin
      idxPages_17 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h11 == waddr) begin
        idxPages_17 <= _idxPages_T[2:0];
      end
    end
    if (metaReset) begin
      idxPages_18 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h12 == waddr) begin
        idxPages_18 <= _idxPages_T[2:0];
      end
    end
    if (metaReset) begin
      idxPages_19 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h13 == waddr) begin
        idxPages_19 <= _idxPages_T[2:0];
      end
    end
    if (metaReset) begin
      idxPages_20 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h14 == waddr) begin
        idxPages_20 <= _idxPages_T[2:0];
      end
    end
    if (metaReset) begin
      idxPages_21 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h15 == waddr) begin
        idxPages_21 <= _idxPages_T[2:0];
      end
    end
    if (metaReset) begin
      idxPages_22 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h16 == waddr) begin
        idxPages_22 <= _idxPages_T[2:0];
      end
    end
    if (metaReset) begin
      idxPages_23 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h17 == waddr) begin
        idxPages_23 <= _idxPages_T[2:0];
      end
    end
    if (metaReset) begin
      idxPages_24 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h18 == waddr) begin
        idxPages_24 <= _idxPages_T[2:0];
      end
    end
    if (metaReset) begin
      idxPages_25 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h19 == waddr) begin
        idxPages_25 <= _idxPages_T[2:0];
      end
    end
    if (metaReset) begin
      idxPages_26 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h1a == waddr) begin
        idxPages_26 <= _idxPages_T[2:0];
      end
    end
    if (metaReset) begin
      idxPages_27 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h1b == waddr) begin
        idxPages_27 <= _idxPages_T[2:0];
      end
    end
    if (metaReset) begin
      tgts_0 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h0 == waddr) begin
        tgts_0 <= idxHit_idx;
      end
    end
    if (metaReset) begin
      tgts_1 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h1 == waddr) begin
        tgts_1 <= idxHit_idx;
      end
    end
    if (metaReset) begin
      tgts_2 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h2 == waddr) begin
        tgts_2 <= idxHit_idx;
      end
    end
    if (metaReset) begin
      tgts_3 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h3 == waddr) begin
        tgts_3 <= idxHit_idx;
      end
    end
    if (metaReset) begin
      tgts_4 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h4 == waddr) begin
        tgts_4 <= idxHit_idx;
      end
    end
    if (metaReset) begin
      tgts_5 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h5 == waddr) begin
        tgts_5 <= idxHit_idx;
      end
    end
    if (metaReset) begin
      tgts_6 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h6 == waddr) begin
        tgts_6 <= idxHit_idx;
      end
    end
    if (metaReset) begin
      tgts_7 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h7 == waddr) begin
        tgts_7 <= idxHit_idx;
      end
    end
    if (metaReset) begin
      tgts_8 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h8 == waddr) begin
        tgts_8 <= idxHit_idx;
      end
    end
    if (metaReset) begin
      tgts_9 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h9 == waddr) begin
        tgts_9 <= idxHit_idx;
      end
    end
    if (metaReset) begin
      tgts_10 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'ha == waddr) begin
        tgts_10 <= idxHit_idx;
      end
    end
    if (metaReset) begin
      tgts_11 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hb == waddr) begin
        tgts_11 <= idxHit_idx;
      end
    end
    if (metaReset) begin
      tgts_12 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hc == waddr) begin
        tgts_12 <= idxHit_idx;
      end
    end
    if (metaReset) begin
      tgts_13 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hd == waddr) begin
        tgts_13 <= idxHit_idx;
      end
    end
    if (metaReset) begin
      tgts_14 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'he == waddr) begin
        tgts_14 <= idxHit_idx;
      end
    end
    if (metaReset) begin
      tgts_15 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hf == waddr) begin
        tgts_15 <= idxHit_idx;
      end
    end
    if (metaReset) begin
      tgts_16 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h10 == waddr) begin
        tgts_16 <= idxHit_idx;
      end
    end
    if (metaReset) begin
      tgts_17 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h11 == waddr) begin
        tgts_17 <= idxHit_idx;
      end
    end
    if (metaReset) begin
      tgts_18 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h12 == waddr) begin
        tgts_18 <= idxHit_idx;
      end
    end
    if (metaReset) begin
      tgts_19 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h13 == waddr) begin
        tgts_19 <= idxHit_idx;
      end
    end
    if (metaReset) begin
      tgts_20 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h14 == waddr) begin
        tgts_20 <= idxHit_idx;
      end
    end
    if (metaReset) begin
      tgts_21 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h15 == waddr) begin
        tgts_21 <= idxHit_idx;
      end
    end
    if (metaReset) begin
      tgts_22 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h16 == waddr) begin
        tgts_22 <= idxHit_idx;
      end
    end
    if (metaReset) begin
      tgts_23 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h17 == waddr) begin
        tgts_23 <= idxHit_idx;
      end
    end
    if (metaReset) begin
      tgts_24 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h18 == waddr) begin
        tgts_24 <= idxHit_idx;
      end
    end
    if (metaReset) begin
      tgts_25 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h19 == waddr) begin
        tgts_25 <= idxHit_idx;
      end
    end
    if (metaReset) begin
      tgts_26 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h1a == waddr) begin
        tgts_26 <= idxHit_idx;
      end
    end
    if (metaReset) begin
      tgts_27 <= 13'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h1b == waddr) begin
        tgts_27 <= idxHit_idx;
      end
    end
    if (metaReset) begin
      tgtPages_0 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h0 == waddr) begin
        tgtPages_0 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_1 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h1 == waddr) begin
        tgtPages_1 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_2 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h2 == waddr) begin
        tgtPages_2 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_3 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h3 == waddr) begin
        tgtPages_3 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_4 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h4 == waddr) begin
        tgtPages_4 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_5 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h5 == waddr) begin
        tgtPages_5 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_6 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h6 == waddr) begin
        tgtPages_6 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_7 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h7 == waddr) begin
        tgtPages_7 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_8 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h8 == waddr) begin
        tgtPages_8 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_9 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h9 == waddr) begin
        tgtPages_9 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_10 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'ha == waddr) begin
        tgtPages_10 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_11 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hb == waddr) begin
        tgtPages_11 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_12 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hc == waddr) begin
        tgtPages_12 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_13 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hd == waddr) begin
        tgtPages_13 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_14 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'he == waddr) begin
        tgtPages_14 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_15 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hf == waddr) begin
        tgtPages_15 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_16 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h10 == waddr) begin
        tgtPages_16 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_17 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h11 == waddr) begin
        tgtPages_17 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_18 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h12 == waddr) begin
        tgtPages_18 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_19 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h13 == waddr) begin
        tgtPages_19 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_20 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h14 == waddr) begin
        tgtPages_20 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_21 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h15 == waddr) begin
        tgtPages_21 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_22 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h16 == waddr) begin
        tgtPages_22 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_23 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h17 == waddr) begin
        tgtPages_23 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_24 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h18 == waddr) begin
        tgtPages_24 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_25 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h19 == waddr) begin
        tgtPages_25 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_26 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h1a == waddr) begin
        tgtPages_26 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      tgtPages_27 <= 3'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h1b == waddr) begin
        tgtPages_27 <= tgtPageUpdate;
      end
    end
    if (metaReset) begin
      pages_0 <= 25'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (_T_5[0]) begin
        if (idxWritesEven) begin
          pages_0 <= updatePageHit_p;
        end else begin
          pages_0 <= pageHit_p;
        end
      end
    end
    if (metaReset) begin
      pages_1 <= 25'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (_T_12[1]) begin
        if (idxWritesEven) begin
          pages_1 <= pageHit_p;
        end else begin
          pages_1 <= updatePageHit_p;
        end
      end
    end
    if (metaReset) begin
      pages_2 <= 25'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (_T_5[2]) begin
        if (idxWritesEven) begin
          pages_2 <= updatePageHit_p;
        end else begin
          pages_2 <= pageHit_p;
        end
      end
    end
    if (metaReset) begin
      pages_3 <= 25'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (_T_12[3]) begin
        if (idxWritesEven) begin
          pages_3 <= pageHit_p;
        end else begin
          pages_3 <= updatePageHit_p;
        end
      end
    end
    if (metaReset) begin
      pages_4 <= 25'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (_T_5[4]) begin
        if (idxWritesEven) begin
          pages_4 <= updatePageHit_p;
        end else begin
          pages_4 <= pageHit_p;
        end
      end
    end
    if (metaReset) begin
      pages_5 <= 25'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (_T_12[5]) begin
        if (idxWritesEven) begin
          pages_5 <= pageHit_p;
        end else begin
          pages_5 <= updatePageHit_p;
        end
      end
    end
    if (metaReset) begin
      pageValid <= 6'h0;
    end else if (reset) begin
      pageValid <= 6'h0;
    end else begin
      pageValid <= _GEN_373[5:0];
    end
    if (metaReset) begin
      isValid <= 28'h0;
    end else if (reset) begin
      isValid <= 28'h0;
    end else begin
      isValid <= _GEN_375[27:0];
    end
    if (metaReset) begin
      cfiType_0 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h0 == waddr) begin
        cfiType_0 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_1 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h1 == waddr) begin
        cfiType_1 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_2 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h2 == waddr) begin
        cfiType_2 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_3 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h3 == waddr) begin
        cfiType_3 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_4 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h4 == waddr) begin
        cfiType_4 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_5 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h5 == waddr) begin
        cfiType_5 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_6 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h6 == waddr) begin
        cfiType_6 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_7 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h7 == waddr) begin
        cfiType_7 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_8 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h8 == waddr) begin
        cfiType_8 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_9 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h9 == waddr) begin
        cfiType_9 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_10 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'ha == waddr) begin
        cfiType_10 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_11 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hb == waddr) begin
        cfiType_11 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_12 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hc == waddr) begin
        cfiType_12 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_13 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hd == waddr) begin
        cfiType_13 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_14 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'he == waddr) begin
        cfiType_14 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_15 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hf == waddr) begin
        cfiType_15 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_16 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h10 == waddr) begin
        cfiType_16 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_17 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h11 == waddr) begin
        cfiType_17 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_18 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h12 == waddr) begin
        cfiType_18 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_19 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h13 == waddr) begin
        cfiType_19 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_20 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h14 == waddr) begin
        cfiType_20 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_21 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h15 == waddr) begin
        cfiType_21 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_22 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h16 == waddr) begin
        cfiType_22 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_23 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h17 == waddr) begin
        cfiType_23 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_24 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h18 == waddr) begin
        cfiType_24 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_25 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h19 == waddr) begin
        cfiType_25 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_26 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h1a == waddr) begin
        cfiType_26 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      cfiType_27 <= 2'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h1b == waddr) begin
        cfiType_27 <= r_btb_updatePipe_bits_cfiType;
      end
    end
    if (metaReset) begin
      brIdx_0 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h0 == waddr) begin
        brIdx_0 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_1 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h1 == waddr) begin
        brIdx_1 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_2 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h2 == waddr) begin
        brIdx_2 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_3 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h3 == waddr) begin
        brIdx_3 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_4 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h4 == waddr) begin
        brIdx_4 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_5 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h5 == waddr) begin
        brIdx_5 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_6 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h6 == waddr) begin
        brIdx_6 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_7 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h7 == waddr) begin
        brIdx_7 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_8 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h8 == waddr) begin
        brIdx_8 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_9 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h9 == waddr) begin
        brIdx_9 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_10 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'ha == waddr) begin
        brIdx_10 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_11 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hb == waddr) begin
        brIdx_11 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_12 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hc == waddr) begin
        brIdx_12 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_13 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hd == waddr) begin
        brIdx_13 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_14 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'he == waddr) begin
        brIdx_14 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_15 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'hf == waddr) begin
        brIdx_15 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_16 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h10 == waddr) begin
        brIdx_16 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_17 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h11 == waddr) begin
        brIdx_17 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_18 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h12 == waddr) begin
        brIdx_18 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_19 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h13 == waddr) begin
        brIdx_19 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_20 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h14 == waddr) begin
        brIdx_20 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_21 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h15 == waddr) begin
        brIdx_21 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_22 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h16 == waddr) begin
        brIdx_22 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_23 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h17 == waddr) begin
        brIdx_23 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_24 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h18 == waddr) begin
        brIdx_24 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_25 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h19 == waddr) begin
        brIdx_25 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_26 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h1a == waddr) begin
        brIdx_26 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      brIdx_27 <= 1'h0;
    end else if (r_btb_updatePipe_valid) begin
      if (5'h1b == waddr) begin
        brIdx_27 <= r_btb_updatePipe_bits_br_pc[1];
      end
    end
    if (metaReset) begin
      r_btb_updatePipe_valid <= 1'h0;
    end else if (reset) begin
      r_btb_updatePipe_valid <= 1'h0;
    end else begin
      r_btb_updatePipe_valid <= io_btb_update_valid;
    end
    if (metaReset) begin
      r_btb_updatePipe_bits_prediction_entry <= 5'h0;
    end else if (io_btb_update_valid) begin
      r_btb_updatePipe_bits_prediction_entry <= io_btb_update_bits_prediction_entry;
    end
    if (metaReset) begin
      r_btb_updatePipe_bits_pc <= 39'h0;
    end else if (io_btb_update_valid) begin
      r_btb_updatePipe_bits_pc <= io_btb_update_bits_pc;
    end
    if (metaReset) begin
      r_btb_updatePipe_bits_isValid <= 1'h0;
    end else if (io_btb_update_valid) begin
      r_btb_updatePipe_bits_isValid <= io_btb_update_bits_isValid;
    end
    if (metaReset) begin
      r_btb_updatePipe_bits_br_pc <= 39'h0;
    end else if (io_btb_update_valid) begin
      r_btb_updatePipe_bits_br_pc <= io_btb_update_bits_br_pc;
    end
    if (metaReset) begin
      r_btb_updatePipe_bits_cfiType <= 2'h0;
    end else if (io_btb_update_valid) begin
      r_btb_updatePipe_bits_cfiType <= io_btb_update_bits_cfiType;
    end
    if (metaReset) begin
      nextPageRepl <= 3'h0;
    end else if (reset) begin
      nextPageRepl <= 3'h0;
    end else if (_T_1) begin
      if (_nextPageRepl_T) begin
        nextPageRepl <= {{2'd0}, next[0]};
      end else begin
        nextPageRepl <= next;
      end
    end
    if (metaReset) begin
      state_reg <= 27'h0;
    end else if (reset) begin
      state_reg <= 27'h0;
    end else if (_T_3) begin
      state_reg <= _state_reg_T_66;
    end
    if (metaReset) begin
      r_respPipe_valid <= 1'h0;
    end else if (reset) begin
      r_respPipe_valid <= 1'h0;
    end else begin
      r_respPipe_valid <= io_resp_valid;
    end
    if (metaReset) begin
      r_respPipe_bits_taken <= 1'h0;
    end else if (io_resp_valid) begin
      r_respPipe_bits_taken <= io_resp_bits_taken;
    end
    if (metaReset) begin
      r_respPipe_bits_entry <= 5'h0;
    end else if (io_resp_valid) begin
      r_respPipe_bits_entry <= io_resp_bits_entry;
    end
    if (metaReset) begin
      history <= 8'h0;
    end else if (reset) begin
      history <= 8'h0;
    end else if (io_bht_update_valid) begin
      if (io_bht_update_bits_branch) begin
        if (io_bht_update_bits_mispredict) begin
          history <= _history_T_1;
        end else if (io_bht_advance_valid) begin
          history <= _history_T;
        end
      end else if (io_bht_update_bits_mispredict) begin
        history <= io_bht_update_bits_prediction_history;
      end else if (io_bht_advance_valid) begin
        history <= _history_T;
      end
    end else if (io_bht_advance_valid) begin
      history <= _history_T;
    end
    if (metaReset) begin
      reset_waddr <= 10'h0;
    end else if (reset) begin
      reset_waddr <= 10'h0;
    end else if (resetting) begin
      reset_waddr <= _reset_waddr_T_1;
    end
    if (metaReset) begin
      count <= 3'h0;
    end else if (reset) begin
      count <= 3'h0;
    end else if (io_ras_update_valid) begin
      if (_T_138) begin
        if (_T_139) begin
          count <= _count_T_1;
        end
      end else if (_T_140) begin
        if (~_io_ras_head_valid_T) begin
          count <= _count_T_3;
        end
      end
    end
    if (metaReset) begin
      pos <= 3'h0;
    end else if (reset) begin
      pos <= 3'h0;
    end else if (io_ras_update_valid) begin
      if (_T_138) begin
        if (_nextPos_T) begin
          pos <= _nextPos_T_3;
        end else begin
          pos <= 3'h0;
        end
      end else if (_T_140) begin
        if (~_io_ras_head_valid_T) begin
          if (_pos_T) begin
            pos <= _pos_T_3;
          end else begin
            pos <= 3'h5;
          end
        end
      end
    end
    if (metaReset) begin
      stack_0 <= 39'h0;
    end else if (io_ras_update_valid) begin
      if (_T_138) begin
        if (3'h0 == nextPos) begin
          stack_0 <= io_ras_update_bits_returnAddr;
        end
      end
    end
    if (metaReset) begin
      stack_1 <= 39'h0;
    end else if (io_ras_update_valid) begin
      if (_T_138) begin
        if (3'h1 == nextPos) begin
          stack_1 <= io_ras_update_bits_returnAddr;
        end
      end
    end
    if (metaReset) begin
      stack_2 <= 39'h0;
    end else if (io_ras_update_valid) begin
      if (_T_138) begin
        if (3'h2 == nextPos) begin
          stack_2 <= io_ras_update_bits_returnAddr;
        end
      end
    end
    if (metaReset) begin
      stack_3 <= 39'h0;
    end else if (io_ras_update_valid) begin
      if (_T_138) begin
        if (3'h3 == nextPos) begin
          stack_3 <= io_ras_update_bits_returnAddr;
        end
      end
    end
    if (metaReset) begin
      stack_4 <= 39'h0;
    end else if (io_ras_update_valid) begin
      if (_T_138) begin
        if (3'h4 == nextPos) begin
          stack_4 <= io_ras_update_bits_returnAddr;
        end
      end
    end
    if (metaReset) begin
      stack_5 <= 39'h0;
    end else if (io_ras_update_valid) begin
      if (_T_138) begin
        if (3'h5 == nextPos) begin
          stack_5 <= io_ras_update_bits_returnAddr;
        end
      end
    end
    BTB_state <= BTB_xor0;
    if (!(BTB_cov_read_data)) begin
      BTB_covSum <= BTB_covSum + 1'h1;
    end
  end
  always @(posedge clock) begin
    if(BTB_cov_write_en & BTB_cov_write_mask) begin
      BTB_cov[BTB_cov_write_addr] <= BTB_cov_write_data; // @[Coverage map for BTB]
    end
  end
endmodule
module FPUDecoder(
  input  [31:0] io_inst,
  output        io_sigs_wen,
  output        io_sigs_ren1,
  output        io_sigs_ren2,
  output        io_sigs_ren3,
  output        io_sigs_swap12,
  output        io_sigs_swap23,
  output [1:0]  io_sigs_typeTagIn,
  output [1:0]  io_sigs_typeTagOut,
  output        io_sigs_fromint,
  output        io_sigs_toint,
  output        io_sigs_fastpipe,
  output        io_sigs_fma,
  output        io_sigs_div,
  output        io_sigs_sqrt,
  output        io_sigs_wflags,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire [31:0] _decoder_T; // @[Decode.scala 14:65]
  wire  decoder_0; // @[Decode.scala 14:121]
  wire [31:0] _decoder_T_2; // @[Decode.scala 14:65]
  wire  _decoder_T_3; // @[Decode.scala 14:121]
  wire [31:0] _decoder_T_4; // @[Decode.scala 14:65]
  wire  _decoder_T_5; // @[Decode.scala 14:121]
  wire [31:0] _decoder_T_6; // @[Decode.scala 14:65]
  wire  _decoder_T_7; // @[Decode.scala 14:121]
  wire  _decoder_T_9; // @[Decode.scala 15:30]
  wire [31:0] _decoder_T_10; // @[Decode.scala 14:65]
  wire  _decoder_T_11; // @[Decode.scala 14:121]
  wire [31:0] _decoder_T_12; // @[Decode.scala 14:65]
  wire  _decoder_T_13; // @[Decode.scala 14:121]
  wire [31:0] _decoder_T_14; // @[Decode.scala 14:65]
  wire  decoder_4; // @[Decode.scala 14:121]
  wire  _decoder_T_17; // @[Decode.scala 15:30]
  wire [31:0] _decoder_T_18; // @[Decode.scala 14:65]
  wire  _decoder_T_19; // @[Decode.scala 14:121]
  wire [31:0] _decoder_T_20; // @[Decode.scala 14:65]
  wire  _decoder_T_21; // @[Decode.scala 14:121]
  wire  _decoder_T_23; // @[Decode.scala 15:30]
  wire [31:0] _decoder_T_24; // @[Decode.scala 14:65]
  wire [31:0] _decoder_T_26; // @[Decode.scala 14:65]
  wire  _decoder_T_27; // @[Decode.scala 14:121]
  wire [31:0] _decoder_T_28; // @[Decode.scala 14:65]
  wire  _decoder_T_29; // @[Decode.scala 14:121]
  wire [31:0] _decoder_T_30; // @[Decode.scala 14:65]
  wire  _decoder_T_31; // @[Decode.scala 14:121]
  wire [31:0] _decoder_T_32; // @[Decode.scala 14:65]
  wire  _decoder_T_33; // @[Decode.scala 14:121]
  wire [31:0] _decoder_T_34; // @[Decode.scala 14:65]
  wire  _decoder_T_35; // @[Decode.scala 14:121]
  wire [31:0] _decoder_T_36; // @[Decode.scala 14:65]
  wire  _decoder_T_37; // @[Decode.scala 14:121]
  wire  _decoder_T_39; // @[Decode.scala 15:30]
  wire  _decoder_T_40; // @[Decode.scala 15:30]
  wire  _decoder_T_41; // @[Decode.scala 15:30]
  wire  _decoder_T_42; // @[Decode.scala 15:30]
  wire  _decoder_T_43; // @[Decode.scala 15:30]
  wire  decoder_7; // @[Decode.scala 15:30]
  wire [31:0] _decoder_T_44; // @[Decode.scala 14:65]
  wire  _decoder_T_45; // @[Decode.scala 14:121]
  wire [31:0] _decoder_T_46; // @[Decode.scala 14:65]
  wire  _decoder_T_47; // @[Decode.scala 14:121]
  wire  _decoder_T_49; // @[Decode.scala 14:121]
  wire  _decoder_T_51; // @[Decode.scala 15:30]
  wire  decoder_8; // @[Decode.scala 15:30]
  wire [31:0] _decoder_T_52; // @[Decode.scala 14:65]
  wire  _decoder_T_55; // @[Decode.scala 14:121]
  wire [31:0] _decoder_T_57; // @[Decode.scala 14:65]
  wire  _decoder_T_58; // @[Decode.scala 14:121]
  wire [31:0] _decoder_T_59; // @[Decode.scala 14:65]
  wire  _decoder_T_60; // @[Decode.scala 14:121]
  wire [31:0] _decoder_T_62; // @[Decode.scala 14:65]
  wire  _decoder_T_63; // @[Decode.scala 14:121]
  wire [31:0] _decoder_T_64; // @[Decode.scala 14:65]
  wire  _decoder_T_65; // @[Decode.scala 14:121]
  wire  _decoder_T_67; // @[Decode.scala 15:30]
  wire [31:0] _decoder_T_68; // @[Decode.scala 14:65]
  wire [31:0] _decoder_T_72; // @[Decode.scala 14:65]
  wire  _decoder_T_73; // @[Decode.scala 14:121]
  wire [31:0] _decoder_T_74; // @[Decode.scala 14:65]
  wire  _decoder_T_75; // @[Decode.scala 14:121]
  wire [31:0] _decoder_T_76; // @[Decode.scala 14:65]
  wire  _decoder_T_77; // @[Decode.scala 14:121]
  wire  _decoder_T_79; // @[Decode.scala 15:30]
  wire  _decoder_T_80; // @[Decode.scala 15:30]
  wire [29:0] FPUDecoder_covSum;
  assign _decoder_T = io_inst & 32'h40; // @[Decode.scala 14:65]
  assign decoder_0 = _decoder_T == 32'h0; // @[Decode.scala 14:121]
  assign _decoder_T_2 = io_inst & 32'h80000020; // @[Decode.scala 14:65]
  assign _decoder_T_3 = _decoder_T_2 == 32'h0; // @[Decode.scala 14:121]
  assign _decoder_T_4 = io_inst & 32'h30; // @[Decode.scala 14:65]
  assign _decoder_T_5 = _decoder_T_4 == 32'h0; // @[Decode.scala 14:121]
  assign _decoder_T_6 = io_inst & 32'h10000020; // @[Decode.scala 14:65]
  assign _decoder_T_7 = _decoder_T_6 == 32'h10000000; // @[Decode.scala 14:121]
  assign _decoder_T_9 = _decoder_T_3 | _decoder_T_5; // @[Decode.scala 15:30]
  assign _decoder_T_10 = io_inst & 32'h80000004; // @[Decode.scala 14:65]
  assign _decoder_T_11 = _decoder_T_10 == 32'h0; // @[Decode.scala 14:121]
  assign _decoder_T_12 = io_inst & 32'h10000004; // @[Decode.scala 14:65]
  assign _decoder_T_13 = _decoder_T_12 == 32'h0; // @[Decode.scala 14:121]
  assign _decoder_T_14 = io_inst & 32'h50; // @[Decode.scala 14:65]
  assign decoder_4 = _decoder_T_14 == 32'h40; // @[Decode.scala 14:121]
  assign _decoder_T_17 = _decoder_T_11 | _decoder_T_13; // @[Decode.scala 15:30]
  assign _decoder_T_18 = io_inst & 32'h40000004; // @[Decode.scala 14:65]
  assign _decoder_T_19 = _decoder_T_18 == 32'h0; // @[Decode.scala 14:121]
  assign _decoder_T_20 = io_inst & 32'h20; // @[Decode.scala 14:65]
  assign _decoder_T_21 = _decoder_T_20 == 32'h20; // @[Decode.scala 14:121]
  assign _decoder_T_23 = _decoder_T_19 | _decoder_T_21; // @[Decode.scala 15:30]
  assign _decoder_T_24 = io_inst & 32'h30000010; // @[Decode.scala 14:65]
  assign _decoder_T_26 = io_inst & 32'h42000000; // @[Decode.scala 14:65]
  assign _decoder_T_27 = _decoder_T_26 == 32'h2000000; // @[Decode.scala 14:121]
  assign _decoder_T_28 = io_inst & 32'h2000010; // @[Decode.scala 14:65]
  assign _decoder_T_29 = _decoder_T_28 == 32'h2000000; // @[Decode.scala 14:121]
  assign _decoder_T_30 = io_inst & 32'h12000000; // @[Decode.scala 14:65]
  assign _decoder_T_31 = _decoder_T_30 == 32'h12000000; // @[Decode.scala 14:121]
  assign _decoder_T_32 = io_inst & 32'hd2000010; // @[Decode.scala 14:65]
  assign _decoder_T_33 = _decoder_T_32 == 32'h40000010; // @[Decode.scala 14:121]
  assign _decoder_T_34 = io_inst & 32'h70001010; // @[Decode.scala 14:65]
  assign _decoder_T_35 = _decoder_T_34 == 32'h60000010; // @[Decode.scala 14:121]
  assign _decoder_T_36 = io_inst & 32'h82000000; // @[Decode.scala 14:65]
  assign _decoder_T_37 = _decoder_T_36 == 32'h82000000; // @[Decode.scala 14:121]
  assign _decoder_T_39 = decoder_0 | _decoder_T_27; // @[Decode.scala 15:30]
  assign _decoder_T_40 = _decoder_T_39 | _decoder_T_29; // @[Decode.scala 15:30]
  assign _decoder_T_41 = _decoder_T_40 | _decoder_T_31; // @[Decode.scala 15:30]
  assign _decoder_T_42 = _decoder_T_41 | _decoder_T_33; // @[Decode.scala 15:30]
  assign _decoder_T_43 = _decoder_T_42 | _decoder_T_35; // @[Decode.scala 15:30]
  assign decoder_7 = _decoder_T_43 | _decoder_T_37; // @[Decode.scala 15:30]
  assign _decoder_T_44 = io_inst & 32'h1040; // @[Decode.scala 14:65]
  assign _decoder_T_45 = _decoder_T_44 == 32'h1000; // @[Decode.scala 14:121]
  assign _decoder_T_46 = io_inst & 32'h2000020; // @[Decode.scala 14:65]
  assign _decoder_T_47 = _decoder_T_46 == 32'h2000000; // @[Decode.scala 14:121]
  assign _decoder_T_49 = _decoder_T_24 == 32'h30000010; // @[Decode.scala 14:121]
  assign _decoder_T_51 = _decoder_T_45 | _decoder_T_47; // @[Decode.scala 15:30]
  assign decoder_8 = _decoder_T_51 | _decoder_T_49; // @[Decode.scala 15:30]
  assign _decoder_T_52 = io_inst & 32'h90000010; // @[Decode.scala 14:65]
  assign _decoder_T_55 = _decoder_T_52 == 32'h80000010; // @[Decode.scala 14:121]
  assign _decoder_T_57 = io_inst & 32'ha0000010; // @[Decode.scala 14:65]
  assign _decoder_T_58 = _decoder_T_57 == 32'h20000010; // @[Decode.scala 14:121]
  assign _decoder_T_59 = io_inst & 32'hd0000010; // @[Decode.scala 14:65]
  assign _decoder_T_60 = _decoder_T_59 == 32'h40000010; // @[Decode.scala 14:121]
  assign _decoder_T_62 = io_inst & 32'h70000004; // @[Decode.scala 14:65]
  assign _decoder_T_63 = _decoder_T_62 == 32'h0; // @[Decode.scala 14:121]
  assign _decoder_T_64 = io_inst & 32'h68000004; // @[Decode.scala 14:65]
  assign _decoder_T_65 = _decoder_T_64 == 32'h0; // @[Decode.scala 14:121]
  assign _decoder_T_67 = _decoder_T_63 | _decoder_T_65; // @[Decode.scala 15:30]
  assign _decoder_T_68 = io_inst & 32'h58000010; // @[Decode.scala 14:65]
  assign _decoder_T_72 = io_inst & 32'h20000004; // @[Decode.scala 14:65]
  assign _decoder_T_73 = _decoder_T_72 == 32'h0; // @[Decode.scala 14:121]
  assign _decoder_T_74 = io_inst & 32'h8002000; // @[Decode.scala 14:65]
  assign _decoder_T_75 = _decoder_T_74 == 32'h8000000; // @[Decode.scala 14:121]
  assign _decoder_T_76 = io_inst & 32'hc0000004; // @[Decode.scala 14:65]
  assign _decoder_T_77 = _decoder_T_76 == 32'h80000000; // @[Decode.scala 14:121]
  assign _decoder_T_79 = _decoder_T_73 | decoder_4; // @[Decode.scala 15:30]
  assign _decoder_T_80 = _decoder_T_79 | _decoder_T_75; // @[Decode.scala 15:30]
  assign io_sigs_wen = _decoder_T_9 | _decoder_T_7; // @[FPU.scala 174:40]
  assign io_sigs_ren1 = _decoder_T_17 | decoder_4; // @[FPU.scala 174:40]
  assign io_sigs_ren2 = _decoder_T_23 | decoder_4; // @[FPU.scala 174:40]
  assign io_sigs_ren3 = _decoder_T_14 == 32'h40; // @[FPU.scala 174:40]
  assign io_sigs_swap12 = _decoder_T == 32'h0; // @[FPU.scala 174:40]
  assign io_sigs_swap23 = _decoder_T_24 == 32'h10; // @[FPU.scala 174:40]
  assign io_sigs_typeTagIn = {{1'd0}, decoder_7}; // @[FPU.scala 174:40]
  assign io_sigs_typeTagOut = {{1'd0}, decoder_8}; // @[FPU.scala 174:40]
  assign io_sigs_fromint = _decoder_T_52 == 32'h90000010; // @[FPU.scala 174:40]
  assign io_sigs_toint = _decoder_T_21 | _decoder_T_55; // @[FPU.scala 174:40]
  assign io_sigs_fastpipe = _decoder_T_58 | _decoder_T_60; // @[FPU.scala 174:40]
  assign io_sigs_fma = _decoder_T_67 | decoder_4; // @[FPU.scala 174:40]
  assign io_sigs_div = _decoder_T_68 == 32'h18000010; // @[FPU.scala 174:40]
  assign io_sigs_sqrt = _decoder_T_59 == 32'h50000010; // @[FPU.scala 174:40]
  assign io_sigs_wflags = _decoder_T_80 | _decoder_T_77; // @[FPU.scala 174:40]
  assign FPUDecoder_covSum = 30'h0;
  assign io_covSum = FPUDecoder_covSum;
  assign metaAssert = 1'h0;
endmodule
module FPUFMAPipe(
  input         clock,
  input         reset,
  input         io_in_valid,
  input         io_in_bits_ren3,
  input         io_in_bits_swap23,
  input  [2:0]  io_in_bits_rm,
  input  [1:0]  io_in_bits_fmaCmd,
  input  [64:0] io_in_bits_in1,
  input  [64:0] io_in_bits_in2,
  input  [64:0] io_in_bits_in3,
  output [64:0] io_out_bits_data,
  output [4:0]  io_out_bits_exc,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset,
  input         fma_halt
);
  wire  fma_clock; // @[FPU.scala 712:19]
  wire  fma_reset; // @[FPU.scala 712:19]
  wire  fma_io_validin; // @[FPU.scala 712:19]
  wire [1:0] fma_io_op; // @[FPU.scala 712:19]
  wire [32:0] fma_io_a; // @[FPU.scala 712:19]
  wire [32:0] fma_io_b; // @[FPU.scala 712:19]
  wire [32:0] fma_io_c; // @[FPU.scala 712:19]
  wire [2:0] fma_io_roundingMode; // @[FPU.scala 712:19]
  wire [32:0] fma_io_out; // @[FPU.scala 712:19]
  wire [4:0] fma_io_exceptionFlags; // @[FPU.scala 712:19]
  wire [29:0] fma_io_covSum; // @[FPU.scala 712:19]
  wire  fma_metaAssert; // @[FPU.scala 712:19]
  wire  fma_metaReset; // @[FPU.scala 712:19]
  reg  valid; // @[FPU.scala 700:18]
  reg [31:0] _RAND_0;
  reg [2:0] in_rm; // @[FPU.scala 701:15]
  reg [31:0] _RAND_1;
  reg [1:0] in_fmaCmd; // @[FPU.scala 701:15]
  reg [31:0] _RAND_2;
  reg [64:0] in_in1; // @[FPU.scala 701:15]
  reg [95:0] _RAND_3;
  reg [64:0] in_in2; // @[FPU.scala 701:15]
  reg [95:0] _RAND_4;
  reg [64:0] in_in3; // @[FPU.scala 701:15]
  reg [95:0] _RAND_5;
  wire [64:0] _zero_T; // @[FPU.scala 704:32]
  wire [64:0] zero; // @[FPU.scala 704:50]
  wire  _T; // @[FPU.scala 709:21]
  wire [29:0] FPUFMAPipe_covSum;
  wire [29:0] fma_sum;
  wire  fma_metaAssert_wire;
  reg  FPUFMAPipe_metaAssert;
  reg [31:0] _RAND_6;
  MulAddRecFNPipe fma ( // @[FPU.scala 712:19]
    .clock(fma_clock),
    .reset(fma_reset),
    .io_validin(fma_io_validin),
    .io_op(fma_io_op),
    .io_a(fma_io_a),
    .io_b(fma_io_b),
    .io_c(fma_io_c),
    .io_roundingMode(fma_io_roundingMode),
    .io_out(fma_io_out),
    .io_exceptionFlags(fma_io_exceptionFlags),
    .io_covSum(fma_io_covSum),
    .metaAssert(fma_metaAssert),
    .metaReset(fma_metaReset)
  );
  assign _zero_T = io_in_bits_in1 ^ io_in_bits_in2; // @[FPU.scala 704:32]
  assign zero = _zero_T & 65'h100000000; // @[FPU.scala 704:50]
  assign _T = io_in_bits_ren3 | io_in_bits_swap23; // @[FPU.scala 709:21]
  assign io_out_bits_data = {{32'd0}, fma_io_out}; // @[FPU.scala 725:10]
  assign io_out_bits_exc = fma_io_exceptionFlags; // @[FPU.scala 725:10]
  assign fma_clock = clock;
  assign fma_reset = reset;
  assign fma_io_validin = valid; // @[FPU.scala 713:18]
  assign fma_io_op = in_fmaCmd; // @[FPU.scala 714:13]
  assign fma_io_a = in_in1[32:0]; // @[FPU.scala 717:12]
  assign fma_io_b = in_in2[32:0]; // @[FPU.scala 718:12]
  assign fma_io_c = in_in3[32:0]; // @[FPU.scala 719:12]
  assign fma_io_roundingMode = in_rm; // @[FPU.scala 715:23]
  assign FPUFMAPipe_covSum = 30'h0;
  assign fma_sum = FPUFMAPipe_covSum + fma_io_covSum;
  assign io_covSum = fma_sum;
  assign fma_metaAssert_wire = fma_metaAssert;
  assign metaAssert = FPUFMAPipe_metaAssert;
  assign fma_metaReset = metaReset | fma_halt;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  valid = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  in_rm = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  in_fmaCmd = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {3{`RANDOM}};
  in_in1 = _RAND_3[64:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {3{`RANDOM}};
  in_in2 = _RAND_4[64:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {3{`RANDOM}};
  in_in3 = _RAND_5[64:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  FPUFMAPipe_metaAssert = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      valid <= 1'h0;
    end else begin
      valid <= io_in_valid;
    end
    if (metaReset) begin
      in_rm <= 3'h0;
    end else if (io_in_valid) begin
      in_rm <= io_in_bits_rm;
    end
    if (metaReset) begin
      in_fmaCmd <= 2'h0;
    end else if (io_in_valid) begin
      in_fmaCmd <= io_in_bits_fmaCmd;
    end
    if (metaReset) begin
      in_in1 <= 65'h0;
    end else if (io_in_valid) begin
      in_in1 <= io_in_bits_in1;
    end
    if (metaReset) begin
      in_in2 <= 65'h0;
    end else if (io_in_valid) begin
      if (io_in_bits_swap23) begin
        in_in2 <= 65'h80000000;
      end else begin
        in_in2 <= io_in_bits_in2;
      end
    end
    if (metaReset) begin
      in_in3 <= 65'h0;
    end else if (io_in_valid) begin
      if (~_T) begin
        in_in3 <= zero;
      end else begin
        in_in3 <= io_in_bits_in3;
      end
    end
    if (metaReset) begin
      FPUFMAPipe_metaAssert <= 1'h0;
    end else begin
      FPUFMAPipe_metaAssert <= FPUFMAPipe_metaAssert | fma_metaAssert_wire;
    end
  end
endmodule
module FPToInt(
  input         clock,
  input         io_in_valid,
  input         io_in_bits_ren2,
  input  [1:0]  io_in_bits_typeTagIn,
  input  [1:0]  io_in_bits_typeTagOut,
  input         io_in_bits_wflags,
  input  [2:0]  io_in_bits_rm,
  input  [1:0]  io_in_bits_typ,
  input  [1:0]  io_in_bits_fmt,
  input  [64:0] io_in_bits_in1,
  input  [64:0] io_in_bits_in2,
  output [2:0]  io_out_bits_in_rm,
  output [64:0] io_out_bits_in_in1,
  output [64:0] io_out_bits_in_in2,
  output        io_out_bits_lt,
  output [63:0] io_out_bits_store,
  output [63:0] io_out_bits_toint,
  output [4:0]  io_out_bits_exc,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  wire [64:0] dcmp_io_a; // @[FPU.scala 465:20]
  wire [64:0] dcmp_io_b; // @[FPU.scala 465:20]
  wire  dcmp_io_signaling; // @[FPU.scala 465:20]
  wire  dcmp_io_lt; // @[FPU.scala 465:20]
  wire  dcmp_io_eq; // @[FPU.scala 465:20]
  wire [4:0] dcmp_io_exceptionFlags; // @[FPU.scala 465:20]
  wire [29:0] dcmp_io_covSum; // @[FPU.scala 465:20]
  wire  dcmp_metaAssert; // @[FPU.scala 465:20]
  wire [64:0] conv_io_in; // @[FPU.scala 493:24]
  wire [2:0] conv_io_roundingMode; // @[FPU.scala 493:24]
  wire  conv_io_signedOut; // @[FPU.scala 493:24]
  wire [63:0] conv_io_out; // @[FPU.scala 493:24]
  wire [2:0] conv_io_intExceptionFlags; // @[FPU.scala 493:24]
  wire [29:0] conv_io_covSum; // @[FPU.scala 493:24]
  wire  conv_metaAssert; // @[FPU.scala 493:24]
  wire [64:0] narrow_io_in; // @[FPU.scala 503:30]
  wire [2:0] narrow_io_roundingMode; // @[FPU.scala 503:30]
  wire  narrow_io_signedOut; // @[FPU.scala 503:30]
  wire [2:0] narrow_io_intExceptionFlags; // @[FPU.scala 503:30]
  wire [29:0] narrow_io_covSum; // @[FPU.scala 503:30]
  wire  narrow_metaAssert; // @[FPU.scala 503:30]
  reg  in_ren2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  reg [1:0] in_typeTagOut; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  reg  in_wflags; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [2:0] in_rm; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg [1:0] in_typ; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg [1:0] in_fmt; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg [64:0] in_in1; // @[Reg.scala 15:16]
  reg [95:0] _RAND_6;
  reg [64:0] in_in2; // @[Reg.scala 15:16]
  reg [95:0] _RAND_7;
  wire [11:0] store_unrecoded_rawIn_exp; // @[rawFloatFromRecFN.scala 50:21]
  wire  store_unrecoded_rawIn_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  store_unrecoded_rawIn_isSpecial; // @[rawFloatFromRecFN.scala 52:54]
  wire  store_unrecoded_rawIn__isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  store_unrecoded_rawIn__isInf; // @[rawFloatFromRecFN.scala 56:33]
  wire  store_unrecoded_rawIn__sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [12:0] store_unrecoded_rawIn__sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire  store_unrecoded_rawIn_out_sig_hi_lo; // @[rawFloatFromRecFN.scala 60:39]
  wire [51:0] store_unrecoded_rawIn_out_sig_lo; // @[rawFloatFromRecFN.scala 60:51]
  wire [53:0] store_unrecoded_rawIn__sig; // @[Cat.scala 30:58]
  wire  store_unrecoded_isSubnormal; // @[fNFromRecFN.scala 50:39]
  wire [5:0] store_unrecoded_denormShiftDist; // @[fNFromRecFN.scala 51:39]
  wire [52:0] _store_unrecoded_denormFract_T_1; // @[fNFromRecFN.scala 52:42]
  wire [51:0] store_unrecoded_denormFract; // @[fNFromRecFN.scala 52:60]
  wire [10:0] _store_unrecoded_expOut_T_2; // @[fNFromRecFN.scala 57:45]
  wire [10:0] _store_unrecoded_expOut_T_3; // @[fNFromRecFN.scala 55:16]
  wire  _store_unrecoded_expOut_T_4; // @[fNFromRecFN.scala 59:44]
  wire [10:0] _store_unrecoded_expOut_T_6; // @[Bitwise.scala 72:12]
  wire [10:0] store_unrecoded_hi_lo; // @[fNFromRecFN.scala 59:15]
  wire [51:0] _store_unrecoded_fractOut_T_1; // @[fNFromRecFN.scala 63:20]
  wire [51:0] store_unrecoded_lo; // @[fNFromRecFN.scala 61:16]
  wire [63:0] store_unrecoded; // @[Cat.scala 30:58]
  wire  store_prevRecoded_hi_hi; // @[FPU.scala 437:10]
  wire  store_prevRecoded_hi_lo; // @[FPU.scala 438:10]
  wire [30:0] store_prevRecoded_lo; // @[FPU.scala 439:10]
  wire [32:0] store_prevRecoded; // @[Cat.scala 30:58]
  wire [8:0] store_prevUnrecoded_rawIn_exp; // @[rawFloatFromRecFN.scala 50:21]
  wire  store_prevUnrecoded_rawIn_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  store_prevUnrecoded_rawIn_isSpecial; // @[rawFloatFromRecFN.scala 52:54]
  wire  store_prevUnrecoded_rawIn__isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  store_prevUnrecoded_rawIn__isInf; // @[rawFloatFromRecFN.scala 56:33]
  wire  store_prevUnrecoded_rawIn__sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [9:0] store_prevUnrecoded_rawIn__sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire  store_prevUnrecoded_rawIn_out_sig_hi_lo; // @[rawFloatFromRecFN.scala 60:39]
  wire [22:0] store_prevUnrecoded_rawIn_out_sig_lo; // @[rawFloatFromRecFN.scala 60:51]
  wire [24:0] store_prevUnrecoded_rawIn__sig; // @[Cat.scala 30:58]
  wire  store_prevUnrecoded_isSubnormal; // @[fNFromRecFN.scala 50:39]
  wire [4:0] store_prevUnrecoded_denormShiftDist; // @[fNFromRecFN.scala 51:39]
  wire [23:0] _store_prevUnrecoded_denormFract_T_1; // @[fNFromRecFN.scala 52:42]
  wire [22:0] store_prevUnrecoded_denormFract; // @[fNFromRecFN.scala 52:60]
  wire [7:0] _store_prevUnrecoded_expOut_T_2; // @[fNFromRecFN.scala 57:45]
  wire [7:0] _store_prevUnrecoded_expOut_T_3; // @[fNFromRecFN.scala 55:16]
  wire  _store_prevUnrecoded_expOut_T_4; // @[fNFromRecFN.scala 59:44]
  wire [7:0] _store_prevUnrecoded_expOut_T_6; // @[Bitwise.scala 72:12]
  wire [7:0] store_prevUnrecoded_hi_lo; // @[fNFromRecFN.scala 59:15]
  wire [22:0] _store_prevUnrecoded_fractOut_T_1; // @[fNFromRecFN.scala 63:20]
  wire [22:0] store_prevUnrecoded_lo; // @[fNFromRecFN.scala 61:16]
  wire [31:0] store_prevUnrecoded; // @[Cat.scala 30:58]
  wire [31:0] store_hi; // @[FPU.scala 441:21]
  wire  _store_T_1; // @[FPU.scala 243:56]
  wire [31:0] store_lo; // @[FPU.scala 441:44]
  wire [63:0] _store_T_3; // @[Cat.scala 30:58]
  wire [31:0] store_hi_1; // @[FPU.scala 472:104]
  wire [63:0] _store_T_4; // @[Cat.scala 30:58]
  wire  store_truncIdx; // @[package.scala 31:49]
  wire [63:0] store; // @[package.scala 32:76]
  wire  intType_x6; // @[FPU.scala 474:35]
  wire  cvtType; // @[package.scala 154:13]
  wire  io_out_bits_exc_hi_hi_1; // @[FPU.scala 510:54]
  wire [31:0] toint_hi; // @[FPU.scala 511:53]
  wire  excSign; // @[FPU.scala 508:59]
  wire  excOut_hi; // @[FPU.scala 509:46]
  wire [30:0] excOut_lo; // @[Bitwise.scala 72:12]
  wire [63:0] _toint_T_10; // @[Cat.scala 30:58]
  wire [63:0] _GEN_25; // @[FPU.scala 511:26]
  wire [63:0] _GEN_26; // @[FPU.scala 502:30]
  wire [1:0] _toint_T_4; // @[Cat.scala 30:58]
  wire [2:0] _GEN_34; // @[FPU.scala 486:22]
  wire [2:0] _toint_T_5; // @[FPU.scala 486:22]
  wire  _toint_T_6; // @[FPU.scala 486:53]
  wire [63:0] _toint_T_8; // @[FPU.scala 486:77]
  wire [63:0] _GEN_35; // @[FPU.scala 486:57]
  wire [63:0] _toint_T_9; // @[FPU.scala 486:57]
  wire [63:0] _GEN_29; // @[FPU.scala 490:21]
  wire  classify_out_hi_hi_hi_hi_1; // @[FPU.scala 259:24]
  wire  classify_out_hi_hi_hi_lo_1; // @[FPU.scala 258:24]
  wire [1:0] classify_out_codeHi_1; // @[FPU.scala 249:22]
  wire  classify_out_isSpecial_1; // @[FPU.scala 250:28]
  wire  classify_out_isInf_1; // @[FPU.scala 256:27]
  wire  classify_out_hi_hi_lo_1; // @[FPU.scala 261:31]
  wire  _classify_out_isNormal_T_4; // @[FPU.scala 254:27]
  wire  classify_out_isHighSubnormalIn_1; // @[FPU.scala 252:55]
  wire  _classify_out_isNormal_T_6; // @[FPU.scala 254:39]
  wire  _classify_out_isNormal_T_7; // @[FPU.scala 254:71]
  wire  classify_out_isNormal_1; // @[FPU.scala 254:61]
  wire  classify_out_hi_lo_hi_1; // @[FPU.scala 261:50]
  wire  _classify_out_isSubnormal_T_3; // @[FPU.scala 253:28]
  wire  _classify_out_isSubnormal_T_5; // @[FPU.scala 253:62]
  wire  classify_out_isSubnormal_1; // @[FPU.scala 253:40]
  wire  classify_out_hi_lo_lo_1; // @[FPU.scala 262:21]
  wire  classify_out_isZero_1; // @[FPU.scala 255:23]
  wire  classify_out_lo_hi_hi_hi_1; // @[FPU.scala 262:38]
  wire  classify_out_lo_hi_hi_lo_1; // @[FPU.scala 262:55]
  wire  classify_out_lo_hi_lo_1; // @[FPU.scala 263:21]
  wire  classify_out_lo_lo_hi_1; // @[FPU.scala 263:39]
  wire  classify_out_lo_lo_lo_1; // @[FPU.scala 263:54]
  wire [9:0] _classify_out_T_10; // @[Cat.scala 30:58]
  wire  _classify_out_expOut_T_1; // @[FPU.scala 275:36]
  wire  _classify_out_expOut_T_2; // @[FPU.scala 275:25]
  wire [11:0] _classify_out_expOut_commonCase_T_1; // @[FPU.scala 274:31]
  wire [11:0] classify_out_expOut_commonCase; // @[FPU.scala 274:48]
  wire [5:0] classify_out_expOut_lo; // @[FPU.scala 275:65]
  wire [8:0] _classify_out_expOut_T_3; // @[Cat.scala 30:58]
  wire [8:0] classify_out_hi_lo; // @[FPU.scala 275:10]
  wire [75:0] _classify_out_fractOut_T; // @[FPU.scala 271:28]
  wire [22:0] classify_out_lo; // @[FPU.scala 271:38]
  wire [32:0] _classify_out_T; // @[Cat.scala 30:58]
  wire [2:0] classify_out_code; // @[FPU.scala 248:17]
  wire  classify_out_isNaN; // @[FPU.scala 257:22]
  wire  classify_out_hi_hi_hi_hi; // @[FPU.scala 259:24]
  wire  classify_out_hi_hi_hi_lo; // @[FPU.scala 258:24]
  wire [1:0] classify_out_codeHi; // @[FPU.scala 249:22]
  wire  classify_out_isSpecial; // @[FPU.scala 250:28]
  wire  classify_out_isInf; // @[FPU.scala 256:27]
  wire  classify_out_sign; // @[FPU.scala 247:17]
  wire  classify_out_hi_hi_lo; // @[FPU.scala 261:31]
  wire  _classify_out_isNormal_T; // @[FPU.scala 254:27]
  wire  classify_out_isHighSubnormalIn; // @[FPU.scala 252:55]
  wire  _classify_out_isNormal_T_2; // @[FPU.scala 254:39]
  wire  _classify_out_isNormal_T_3; // @[FPU.scala 254:71]
  wire  classify_out_isNormal; // @[FPU.scala 254:61]
  wire  classify_out_hi_lo_hi; // @[FPU.scala 261:50]
  wire  _classify_out_isSubnormal_T; // @[FPU.scala 253:28]
  wire  _classify_out_isSubnormal_T_2; // @[FPU.scala 253:62]
  wire  classify_out_isSubnormal; // @[FPU.scala 253:40]
  wire  classify_out_hi_lo_lo; // @[FPU.scala 262:21]
  wire  classify_out_isZero; // @[FPU.scala 255:23]
  wire  classify_out_lo_hi_hi_hi; // @[FPU.scala 262:38]
  wire  classify_out_lo_hi_hi_lo; // @[FPU.scala 262:55]
  wire  classify_out_lo_hi_lo; // @[FPU.scala 263:21]
  wire  classify_out_lo_lo_hi; // @[FPU.scala 263:39]
  wire  classify_out_lo_lo_lo; // @[FPU.scala 263:54]
  wire [9:0] _classify_out_T_5; // @[Cat.scala 30:58]
  wire [9:0] classify_out; // @[package.scala 32:76]
  wire [63:0] _GEN_36; // @[FPU.scala 481:27]
  wire [63:0] _toint_T_2; // @[FPU.scala 481:27]
  wire [63:0] _GEN_23; // @[FPU.scala 479:19]
  wire [63:0] toint; // @[FPU.scala 485:20]
  wire [31:0] io_out_bits_toint_lo; // @[FPU.scala 476:59]
  wire [31:0] io_out_bits_toint_hi; // @[Bitwise.scala 72:12]
  wire [63:0] _io_out_bits_toint_T_2; // @[Cat.scala 30:58]
  wire  _GEN_28; // @[FPU.scala 490:21]
  wire  _GEN_24; // @[FPU.scala 479:19]
  wire  intType; // @[FPU.scala 485:20]
  wire  io_out_bits_exc_hi_hi; // @[FPU.scala 498:62]
  wire  io_out_bits_exc_lo; // @[FPU.scala 498:104]
  wire [4:0] _io_out_bits_exc_T_1; // @[Cat.scala 30:58]
  wire  io_out_bits_exc_lo_1; // @[FPU.scala 512:64]
  wire [4:0] _io_out_bits_exc_T_4; // @[Cat.scala 30:58]
  wire [4:0] _GEN_27; // @[FPU.scala 502:30]
  wire [4:0] _GEN_30; // @[FPU.scala 490:21]
  wire  _io_out_bits_lt_T_1; // @[FPU.scala 519:53]
  wire  _io_out_bits_lt_T_3; // @[FPU.scala 519:79]
  wire  _io_out_bits_lt_T_4; // @[FPU.scala 519:59]
  reg [3:0] FPToInt_state; // @[Register tracking FPToInt state]
  reg [31:0] _RAND_8;
  reg  FPToInt_cov [0:15]; // @[Coverage map for FPToInt]
  reg [31:0] _RAND_9;
  wire  FPToInt_cov_read_data; // @[Coverage map for FPToInt]
  wire [3:0] FPToInt_cov_read_addr; // @[Coverage map for FPToInt]
  wire  FPToInt_cov_write_data; // @[Coverage map for FPToInt]
  wire [3:0] FPToInt_cov_write_addr; // @[Coverage map for FPToInt]
  wire  FPToInt_cov_write_mask; // @[Coverage map for FPToInt]
  wire  FPToInt_cov_write_en; // @[Coverage map for FPToInt]
  reg [29:0] FPToInt_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_10;
  wire  in_wflags_shl;
  wire [3:0] in_wflags_pad;
  wire [2:0] in_typ_shl;
  wire [3:0] in_typ_pad;
  wire [3:0] in_ren2_shl;
  wire [3:0] in_ren2_pad;
  wire [3:0] FPToInt_xor2;
  wire [3:0] FPToInt_xor0;
  wire [29:0] dcmp_sum;
  wire [29:0] conv_sum;
  wire [29:0] narrow_sum;
  wire  dcmp_metaAssert_wire;
  wire  conv_metaAssert_wire;
  wire  narrow_metaAssert_wire;
  wire  FPToInt_or2;
  wire  FPToInt_or0;
  CompareRecFN dcmp ( // @[FPU.scala 465:20]
    .io_a(dcmp_io_a),
    .io_b(dcmp_io_b),
    .io_signaling(dcmp_io_signaling),
    .io_lt(dcmp_io_lt),
    .io_eq(dcmp_io_eq),
    .io_exceptionFlags(dcmp_io_exceptionFlags),
    .io_covSum(dcmp_io_covSum),
    .metaAssert(dcmp_metaAssert)
  );
  RecFNToIN conv ( // @[FPU.scala 493:24]
    .io_in(conv_io_in),
    .io_roundingMode(conv_io_roundingMode),
    .io_signedOut(conv_io_signedOut),
    .io_out(conv_io_out),
    .io_intExceptionFlags(conv_io_intExceptionFlags),
    .io_covSum(conv_io_covSum),
    .metaAssert(conv_metaAssert)
  );
  RecFNToIN_1 narrow ( // @[FPU.scala 503:30]
    .io_in(narrow_io_in),
    .io_roundingMode(narrow_io_roundingMode),
    .io_signedOut(narrow_io_signedOut),
    .io_intExceptionFlags(narrow_io_intExceptionFlags),
    .io_covSum(narrow_io_covSum),
    .metaAssert(narrow_metaAssert)
  );
  assign store_unrecoded_rawIn_exp = in_in1[63:52]; // @[rawFloatFromRecFN.scala 50:21]
  assign store_unrecoded_rawIn_isZero = store_unrecoded_rawIn_exp[11:9] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign store_unrecoded_rawIn_isSpecial = store_unrecoded_rawIn_exp[11:10] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign store_unrecoded_rawIn__isNaN = store_unrecoded_rawIn_isSpecial & store_unrecoded_rawIn_exp[9]; // @[rawFloatFromRecFN.scala 55:33]
  assign store_unrecoded_rawIn__isInf = store_unrecoded_rawIn_isSpecial & ~store_unrecoded_rawIn_exp[9]; // @[rawFloatFromRecFN.scala 56:33]
  assign store_unrecoded_rawIn__sign = in_in1[64]; // @[rawFloatFromRecFN.scala 58:25]
  assign store_unrecoded_rawIn__sExp = {1'b0,$signed(store_unrecoded_rawIn_exp)}; // @[rawFloatFromRecFN.scala 59:27]
  assign store_unrecoded_rawIn_out_sig_hi_lo = ~store_unrecoded_rawIn_isZero; // @[rawFloatFromRecFN.scala 60:39]
  assign store_unrecoded_rawIn_out_sig_lo = in_in1[51:0]; // @[rawFloatFromRecFN.scala 60:51]
  assign store_unrecoded_rawIn__sig = {1'h0,store_unrecoded_rawIn_out_sig_hi_lo,store_unrecoded_rawIn_out_sig_lo}; // @[Cat.scala 30:58]
  assign store_unrecoded_isSubnormal = $signed(store_unrecoded_rawIn__sExp) < 13'sh402; // @[fNFromRecFN.scala 50:39]
  assign store_unrecoded_denormShiftDist = 6'h1 - store_unrecoded_rawIn__sExp[5:0]; // @[fNFromRecFN.scala 51:39]
  assign _store_unrecoded_denormFract_T_1 = store_unrecoded_rawIn__sig[53:1] >> store_unrecoded_denormShiftDist; // @[fNFromRecFN.scala 52:42]
  assign store_unrecoded_denormFract = _store_unrecoded_denormFract_T_1[51:0]; // @[fNFromRecFN.scala 52:60]
  assign _store_unrecoded_expOut_T_2 = store_unrecoded_rawIn__sExp[10:0] - 11'h401; // @[fNFromRecFN.scala 57:45]
  assign _store_unrecoded_expOut_T_3 = store_unrecoded_isSubnormal ? 11'h0 : _store_unrecoded_expOut_T_2; // @[fNFromRecFN.scala 55:16]
  assign _store_unrecoded_expOut_T_4 = store_unrecoded_rawIn__isNaN | store_unrecoded_rawIn__isInf; // @[fNFromRecFN.scala 59:44]
  assign _store_unrecoded_expOut_T_6 = _store_unrecoded_expOut_T_4 ? 11'h7ff : 11'h0; // @[Bitwise.scala 72:12]
  assign store_unrecoded_hi_lo = _store_unrecoded_expOut_T_3 | _store_unrecoded_expOut_T_6; // @[fNFromRecFN.scala 59:15]
  assign _store_unrecoded_fractOut_T_1 = store_unrecoded_rawIn__isInf ? 52'h0 : store_unrecoded_rawIn__sig[51:0]; // @[fNFromRecFN.scala 63:20]
  assign store_unrecoded_lo = store_unrecoded_isSubnormal ? store_unrecoded_denormFract : _store_unrecoded_fractOut_T_1; // @[fNFromRecFN.scala 61:16]
  assign store_unrecoded = {store_unrecoded_rawIn__sign,store_unrecoded_hi_lo,store_unrecoded_lo}; // @[Cat.scala 30:58]
  assign store_prevRecoded_hi_hi = in_in1[31]; // @[FPU.scala 437:10]
  assign store_prevRecoded_hi_lo = in_in1[52]; // @[FPU.scala 438:10]
  assign store_prevRecoded_lo = in_in1[30:0]; // @[FPU.scala 439:10]
  assign store_prevRecoded = {store_prevRecoded_hi_hi,store_prevRecoded_hi_lo,store_prevRecoded_lo}; // @[Cat.scala 30:58]
  assign store_prevUnrecoded_rawIn_exp = store_prevRecoded[31:23]; // @[rawFloatFromRecFN.scala 50:21]
  assign store_prevUnrecoded_rawIn_isZero = store_prevUnrecoded_rawIn_exp[8:6] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign store_prevUnrecoded_rawIn_isSpecial = store_prevUnrecoded_rawIn_exp[8:7] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign store_prevUnrecoded_rawIn__isNaN = store_prevUnrecoded_rawIn_isSpecial & store_prevUnrecoded_rawIn_exp[6]; // @[rawFloatFromRecFN.scala 55:33]
  assign store_prevUnrecoded_rawIn__isInf = store_prevUnrecoded_rawIn_isSpecial & ~store_prevUnrecoded_rawIn_exp[6]; // @[rawFloatFromRecFN.scala 56:33]
  assign store_prevUnrecoded_rawIn__sign = store_prevRecoded[32]; // @[rawFloatFromRecFN.scala 58:25]
  assign store_prevUnrecoded_rawIn__sExp = {1'b0,$signed(store_prevUnrecoded_rawIn_exp)}; // @[rawFloatFromRecFN.scala 59:27]
  assign store_prevUnrecoded_rawIn_out_sig_hi_lo = ~store_prevUnrecoded_rawIn_isZero; // @[rawFloatFromRecFN.scala 60:39]
  assign store_prevUnrecoded_rawIn_out_sig_lo = store_prevRecoded[22:0]; // @[rawFloatFromRecFN.scala 60:51]
  assign store_prevUnrecoded_rawIn__sig = {1'h0,store_prevUnrecoded_rawIn_out_sig_hi_lo,store_prevUnrecoded_rawIn_out_sig_lo}; // @[Cat.scala 30:58]
  assign store_prevUnrecoded_isSubnormal = $signed(store_prevUnrecoded_rawIn__sExp) < 10'sh82; // @[fNFromRecFN.scala 50:39]
  assign store_prevUnrecoded_denormShiftDist = 5'h1 - store_prevUnrecoded_rawIn__sExp[4:0]; // @[fNFromRecFN.scala 51:39]
  assign _store_prevUnrecoded_denormFract_T_1 = store_prevUnrecoded_rawIn__sig[24:1] >> store_prevUnrecoded_denormShiftDist; // @[fNFromRecFN.scala 52:42]
  assign store_prevUnrecoded_denormFract = _store_prevUnrecoded_denormFract_T_1[22:0]; // @[fNFromRecFN.scala 52:60]
  assign _store_prevUnrecoded_expOut_T_2 = store_prevUnrecoded_rawIn__sExp[7:0] - 8'h81; // @[fNFromRecFN.scala 57:45]
  assign _store_prevUnrecoded_expOut_T_3 = store_prevUnrecoded_isSubnormal ? 8'h0 : _store_prevUnrecoded_expOut_T_2; // @[fNFromRecFN.scala 55:16]
  assign _store_prevUnrecoded_expOut_T_4 = store_prevUnrecoded_rawIn__isNaN | store_prevUnrecoded_rawIn__isInf; // @[fNFromRecFN.scala 59:44]
  assign _store_prevUnrecoded_expOut_T_6 = _store_prevUnrecoded_expOut_T_4 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign store_prevUnrecoded_hi_lo = _store_prevUnrecoded_expOut_T_3 | _store_prevUnrecoded_expOut_T_6; // @[fNFromRecFN.scala 59:15]
  assign _store_prevUnrecoded_fractOut_T_1 = store_prevUnrecoded_rawIn__isInf ? 23'h0 : store_prevUnrecoded_rawIn__sig[22:0]; // @[fNFromRecFN.scala 63:20]
  assign store_prevUnrecoded_lo = store_prevUnrecoded_isSubnormal ? store_prevUnrecoded_denormFract : _store_prevUnrecoded_fractOut_T_1; // @[fNFromRecFN.scala 61:16]
  assign store_prevUnrecoded = {store_prevUnrecoded_rawIn__sign,store_prevUnrecoded_hi_lo,store_prevUnrecoded_lo}; // @[Cat.scala 30:58]
  assign store_hi = store_unrecoded[63:32]; // @[FPU.scala 441:21]
  assign _store_T_1 = &in_in1[63:61]; // @[FPU.scala 243:56]
  assign store_lo = _store_T_1 ? store_prevUnrecoded : store_unrecoded[31:0]; // @[FPU.scala 441:44]
  assign _store_T_3 = {store_hi,store_lo}; // @[Cat.scala 30:58]
  assign store_hi_1 = _store_T_3[31:0]; // @[FPU.scala 472:104]
  assign _store_T_4 = {store_hi_1,store_hi_1}; // @[Cat.scala 30:58]
  assign store_truncIdx = in_typeTagOut[0]; // @[package.scala 31:49]
  assign store = store_truncIdx ? _store_T_3 : _store_T_4; // @[package.scala 32:76]
  assign intType_x6 = in_fmt[0]; // @[FPU.scala 474:35]
  assign cvtType = in_typ[1]; // @[package.scala 154:13]
  assign io_out_bits_exc_hi_hi_1 = conv_io_intExceptionFlags[2] | narrow_io_intExceptionFlags[1]; // @[FPU.scala 510:54]
  assign toint_hi = conv_io_out[63:32]; // @[FPU.scala 511:53]
  assign excSign = store_unrecoded_rawIn__sign & ~_store_T_1; // @[FPU.scala 508:59]
  assign excOut_hi = conv_io_signedOut == excSign; // @[FPU.scala 509:46]
  assign excOut_lo = excSign ? 31'h0 : 31'h7fffffff; // @[Bitwise.scala 72:12]
  assign _toint_T_10 = {toint_hi,excOut_hi,excOut_lo}; // @[Cat.scala 30:58]
  assign _GEN_25 = io_out_bits_exc_hi_hi_1 ? _toint_T_10 : conv_io_out; // @[FPU.scala 511:26]
  assign _GEN_26 = cvtType ? conv_io_out : _GEN_25; // @[FPU.scala 502:30]
  assign _toint_T_4 = {dcmp_io_lt,dcmp_io_eq}; // @[Cat.scala 30:58]
  assign _GEN_34 = {{1'd0}, _toint_T_4}; // @[FPU.scala 486:22]
  assign _toint_T_5 = ~in_rm & _GEN_34; // @[FPU.scala 486:22]
  assign _toint_T_6 = |_toint_T_5; // @[FPU.scala 486:53]
  assign _toint_T_8 = {store[63:32], 32'h0}; // @[FPU.scala 486:77]
  assign _GEN_35 = {{63'd0}, _toint_T_6}; // @[FPU.scala 486:57]
  assign _toint_T_9 = _GEN_35 | _toint_T_8; // @[FPU.scala 486:57]
  assign _GEN_29 = in_ren2 ? _toint_T_9 : _GEN_26; // @[FPU.scala 490:21]
  assign classify_out_hi_hi_hi_hi_1 = _store_T_1 & in_in1[51]; // @[FPU.scala 259:24]
  assign classify_out_hi_hi_hi_lo_1 = _store_T_1 & ~in_in1[51]; // @[FPU.scala 258:24]
  assign classify_out_codeHi_1 = in_in1[63:62]; // @[FPU.scala 249:22]
  assign classify_out_isSpecial_1 = classify_out_codeHi_1 == 2'h3; // @[FPU.scala 250:28]
  assign classify_out_isInf_1 = classify_out_isSpecial_1 & ~in_in1[61]; // @[FPU.scala 256:27]
  assign classify_out_hi_hi_lo_1 = classify_out_isInf_1 & ~store_unrecoded_rawIn__sign; // @[FPU.scala 261:31]
  assign _classify_out_isNormal_T_4 = classify_out_codeHi_1 == 2'h1; // @[FPU.scala 254:27]
  assign classify_out_isHighSubnormalIn_1 = in_in1[61:52] < 10'h2; // @[FPU.scala 252:55]
  assign _classify_out_isNormal_T_6 = _classify_out_isNormal_T_4 & ~classify_out_isHighSubnormalIn_1; // @[FPU.scala 254:39]
  assign _classify_out_isNormal_T_7 = classify_out_codeHi_1 == 2'h2; // @[FPU.scala 254:71]
  assign classify_out_isNormal_1 = _classify_out_isNormal_T_6 | _classify_out_isNormal_T_7; // @[FPU.scala 254:61]
  assign classify_out_hi_lo_hi_1 = classify_out_isNormal_1 & ~store_unrecoded_rawIn__sign; // @[FPU.scala 261:50]
  assign _classify_out_isSubnormal_T_3 = in_in1[63:61] == 3'h1; // @[FPU.scala 253:28]
  assign _classify_out_isSubnormal_T_5 = _classify_out_isNormal_T_4 & classify_out_isHighSubnormalIn_1; // @[FPU.scala 253:62]
  assign classify_out_isSubnormal_1 = _classify_out_isSubnormal_T_3 | _classify_out_isSubnormal_T_5; // @[FPU.scala 253:40]
  assign classify_out_hi_lo_lo_1 = classify_out_isSubnormal_1 & ~store_unrecoded_rawIn__sign; // @[FPU.scala 262:21]
  assign classify_out_isZero_1 = in_in1[63:61] == 3'h0; // @[FPU.scala 255:23]
  assign classify_out_lo_hi_hi_hi_1 = classify_out_isZero_1 & ~store_unrecoded_rawIn__sign; // @[FPU.scala 262:38]
  assign classify_out_lo_hi_hi_lo_1 = classify_out_isZero_1 & store_unrecoded_rawIn__sign; // @[FPU.scala 262:55]
  assign classify_out_lo_hi_lo_1 = classify_out_isSubnormal_1 & store_unrecoded_rawIn__sign; // @[FPU.scala 263:21]
  assign classify_out_lo_lo_hi_1 = classify_out_isNormal_1 & store_unrecoded_rawIn__sign; // @[FPU.scala 263:39]
  assign classify_out_lo_lo_lo_1 = classify_out_isInf_1 & store_unrecoded_rawIn__sign; // @[FPU.scala 263:54]
  assign _classify_out_T_10 = {classify_out_hi_hi_hi_hi_1,classify_out_hi_hi_hi_lo_1,classify_out_hi_hi_lo_1,classify_out_hi_lo_hi_1,classify_out_hi_lo_lo_1,classify_out_lo_hi_hi_hi_1,classify_out_lo_hi_hi_lo_1,classify_out_lo_hi_lo_1,classify_out_lo_lo_hi_1,classify_out_lo_lo_lo_1}; // @[Cat.scala 30:58]
  assign _classify_out_expOut_T_1 = store_unrecoded_rawIn_exp[11:9] >= 3'h6; // @[FPU.scala 275:36]
  assign _classify_out_expOut_T_2 = store_unrecoded_rawIn_isZero | _classify_out_expOut_T_1; // @[FPU.scala 275:25]
  assign _classify_out_expOut_commonCase_T_1 = store_unrecoded_rawIn_exp + 12'h100; // @[FPU.scala 274:31]
  assign classify_out_expOut_commonCase = _classify_out_expOut_commonCase_T_1 - 12'h800; // @[FPU.scala 274:48]
  assign classify_out_expOut_lo = classify_out_expOut_commonCase[5:0]; // @[FPU.scala 275:65]
  assign _classify_out_expOut_T_3 = {store_unrecoded_rawIn_exp[11:9],classify_out_expOut_lo}; // @[Cat.scala 30:58]
  assign classify_out_hi_lo = _classify_out_expOut_T_2 ? _classify_out_expOut_T_3 : classify_out_expOut_commonCase[8:0]; // @[FPU.scala 275:10]
  assign _classify_out_fractOut_T = {store_unrecoded_rawIn_out_sig_lo, 24'h0}; // @[FPU.scala 271:28]
  assign classify_out_lo = _classify_out_fractOut_T[75:53]; // @[FPU.scala 271:38]
  assign _classify_out_T = {store_unrecoded_rawIn__sign,classify_out_hi_lo,classify_out_lo}; // @[Cat.scala 30:58]
  assign classify_out_code = _classify_out_T[31:29]; // @[FPU.scala 248:17]
  assign classify_out_isNaN = &classify_out_code; // @[FPU.scala 257:22]
  assign classify_out_hi_hi_hi_hi = classify_out_isNaN & _classify_out_T[22]; // @[FPU.scala 259:24]
  assign classify_out_hi_hi_hi_lo = classify_out_isNaN & ~_classify_out_T[22]; // @[FPU.scala 258:24]
  assign classify_out_codeHi = classify_out_code[2:1]; // @[FPU.scala 249:22]
  assign classify_out_isSpecial = classify_out_codeHi == 2'h3; // @[FPU.scala 250:28]
  assign classify_out_isInf = classify_out_isSpecial & ~classify_out_code[0]; // @[FPU.scala 256:27]
  assign classify_out_sign = _classify_out_T[32]; // @[FPU.scala 247:17]
  assign classify_out_hi_hi_lo = classify_out_isInf & ~classify_out_sign; // @[FPU.scala 261:31]
  assign _classify_out_isNormal_T = classify_out_codeHi == 2'h1; // @[FPU.scala 254:27]
  assign classify_out_isHighSubnormalIn = _classify_out_T[29:23] < 7'h2; // @[FPU.scala 252:55]
  assign _classify_out_isNormal_T_2 = _classify_out_isNormal_T & ~classify_out_isHighSubnormalIn; // @[FPU.scala 254:39]
  assign _classify_out_isNormal_T_3 = classify_out_codeHi == 2'h2; // @[FPU.scala 254:71]
  assign classify_out_isNormal = _classify_out_isNormal_T_2 | _classify_out_isNormal_T_3; // @[FPU.scala 254:61]
  assign classify_out_hi_lo_hi = classify_out_isNormal & ~classify_out_sign; // @[FPU.scala 261:50]
  assign _classify_out_isSubnormal_T = classify_out_code == 3'h1; // @[FPU.scala 253:28]
  assign _classify_out_isSubnormal_T_2 = _classify_out_isNormal_T & classify_out_isHighSubnormalIn; // @[FPU.scala 253:62]
  assign classify_out_isSubnormal = _classify_out_isSubnormal_T | _classify_out_isSubnormal_T_2; // @[FPU.scala 253:40]
  assign classify_out_hi_lo_lo = classify_out_isSubnormal & ~classify_out_sign; // @[FPU.scala 262:21]
  assign classify_out_isZero = classify_out_code == 3'h0; // @[FPU.scala 255:23]
  assign classify_out_lo_hi_hi_hi = classify_out_isZero & ~classify_out_sign; // @[FPU.scala 262:38]
  assign classify_out_lo_hi_hi_lo = classify_out_isZero & classify_out_sign; // @[FPU.scala 262:55]
  assign classify_out_lo_hi_lo = classify_out_isSubnormal & classify_out_sign; // @[FPU.scala 263:21]
  assign classify_out_lo_lo_hi = classify_out_isNormal & classify_out_sign; // @[FPU.scala 263:39]
  assign classify_out_lo_lo_lo = classify_out_isInf & classify_out_sign; // @[FPU.scala 263:54]
  assign _classify_out_T_5 = {classify_out_hi_hi_hi_hi,classify_out_hi_hi_hi_lo,classify_out_hi_hi_lo,classify_out_hi_lo_hi,classify_out_hi_lo_lo,classify_out_lo_hi_hi_hi,classify_out_lo_hi_hi_lo,classify_out_lo_hi_lo,classify_out_lo_lo_hi,classify_out_lo_lo_lo}; // @[Cat.scala 30:58]
  assign classify_out = store_truncIdx ? _classify_out_T_10 : _classify_out_T_5; // @[package.scala 32:76]
  assign _GEN_36 = {{54'd0}, classify_out}; // @[FPU.scala 481:27]
  assign _toint_T_2 = _GEN_36 | _toint_T_8; // @[FPU.scala 481:27]
  assign _GEN_23 = in_rm[0] ? _toint_T_2 : store; // @[FPU.scala 479:19]
  assign toint = in_wflags ? _GEN_29 : _GEN_23; // @[FPU.scala 485:20]
  assign io_out_bits_toint_lo = toint[31:0]; // @[FPU.scala 476:59]
  assign io_out_bits_toint_hi = io_out_bits_toint_lo[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  assign _io_out_bits_toint_T_2 = {io_out_bits_toint_hi,io_out_bits_toint_lo}; // @[Cat.scala 30:58]
  assign _GEN_28 = ~in_ren2 & cvtType; // @[FPU.scala 490:21]
  assign _GEN_24 = in_rm[0] ? 1'h0 : intType_x6; // @[FPU.scala 479:19]
  assign intType = in_wflags ? _GEN_28 : _GEN_24; // @[FPU.scala 485:20]
  assign io_out_bits_exc_hi_hi = |conv_io_intExceptionFlags[2:1]; // @[FPU.scala 498:62]
  assign io_out_bits_exc_lo = conv_io_intExceptionFlags[0]; // @[FPU.scala 498:104]
  assign _io_out_bits_exc_T_1 = {io_out_bits_exc_hi_hi,3'h0,io_out_bits_exc_lo}; // @[Cat.scala 30:58]
  assign io_out_bits_exc_lo_1 = ~io_out_bits_exc_hi_hi_1 & io_out_bits_exc_lo; // @[FPU.scala 512:64]
  assign _io_out_bits_exc_T_4 = {io_out_bits_exc_hi_hi_1,3'h0,io_out_bits_exc_lo_1}; // @[Cat.scala 30:58]
  assign _GEN_27 = cvtType ? _io_out_bits_exc_T_1 : _io_out_bits_exc_T_4; // @[FPU.scala 502:30]
  assign _GEN_30 = in_ren2 ? dcmp_io_exceptionFlags : _GEN_27; // @[FPU.scala 490:21]
  assign _io_out_bits_lt_T_1 = $signed(dcmp_io_a) < 65'sh0; // @[FPU.scala 519:53]
  assign _io_out_bits_lt_T_3 = $signed(dcmp_io_b) >= 65'sh0; // @[FPU.scala 519:79]
  assign _io_out_bits_lt_T_4 = _io_out_bits_lt_T_1 & _io_out_bits_lt_T_3; // @[FPU.scala 519:59]
  assign io_out_bits_in_rm = in_rm; // @[FPU.scala 520:18]
  assign io_out_bits_in_in1 = in_in1; // @[FPU.scala 520:18]
  assign io_out_bits_in_in2 = in_in2; // @[FPU.scala 520:18]
  assign io_out_bits_lt = dcmp_io_lt | _io_out_bits_lt_T_4; // @[FPU.scala 519:18]
  assign io_out_bits_store = store_truncIdx ? _store_T_3 : _store_T_4; // @[FPU.scala 475:21]
  assign io_out_bits_toint = intType ? toint : _io_out_bits_toint_T_2; // @[FPU.scala 476:21]
  assign io_out_bits_exc = in_wflags ? _GEN_30 : 5'h0; // @[FPU.scala 477:19 FPU.scala 487:21 FPU.scala 498:23 FPU.scala 512:27]
  assign dcmp_io_a = in_in1; // @[FPU.scala 466:13]
  assign dcmp_io_b = in_in2; // @[FPU.scala 467:13]
  assign dcmp_io_signaling = ~in_rm[1]; // @[FPU.scala 468:21]
  assign conv_io_in = in_in1; // @[FPU.scala 494:18]
  assign conv_io_roundingMode = in_rm; // @[FPU.scala 495:28]
  assign conv_io_signedOut = ~in_typ[0]; // @[FPU.scala 496:25]
  assign narrow_io_in = in_in1; // @[FPU.scala 504:24]
  assign narrow_io_roundingMode = in_rm; // @[FPU.scala 505:34]
  assign narrow_io_signedOut = ~in_typ[0]; // @[FPU.scala 506:31]
  assign FPToInt_cov_read_addr = FPToInt_state;
  assign FPToInt_cov_read_data = FPToInt_cov[FPToInt_cov_read_addr]; // @[Coverage map for FPToInt]
  assign FPToInt_cov_write_data = 1'h1;
  assign FPToInt_cov_write_addr = FPToInt_state;
  assign FPToInt_cov_write_mask = 1'h1;
  assign FPToInt_cov_write_en = 1'h1;
  assign in_wflags_shl = in_wflags;
  assign in_wflags_pad = {3'h0,in_wflags_shl};
  assign in_typ_shl = {in_typ, 1'h0};
  assign in_typ_pad = {1'h0,in_typ_shl};
  assign in_ren2_shl = {in_ren2, 3'h0};
  assign in_ren2_pad = in_ren2_shl;
  assign FPToInt_xor2 = in_typ_pad ^ in_ren2_pad;
  assign FPToInt_xor0 = in_wflags_pad ^ FPToInt_xor2;
  assign dcmp_sum = FPToInt_covSum + dcmp_io_covSum;
  assign conv_sum = dcmp_sum + conv_io_covSum;
  assign narrow_sum = conv_sum + narrow_io_covSum;
  assign io_covSum = narrow_sum;
  assign dcmp_metaAssert_wire = dcmp_metaAssert;
  assign conv_metaAssert_wire = conv_metaAssert;
  assign narrow_metaAssert_wire = narrow_metaAssert;
  assign FPToInt_or2 = conv_metaAssert_wire | narrow_metaAssert_wire;
  assign FPToInt_or0 = dcmp_metaAssert_wire | FPToInt_or2;
  assign metaAssert = FPToInt_or0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  in_ren2 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  in_typeTagOut = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  in_wflags = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  in_rm = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  in_typ = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  in_fmt = _RAND_5[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {3{`RANDOM}};
  in_in1 = _RAND_6[64:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {3{`RANDOM}};
  in_in2 = _RAND_7[64:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  FPToInt_state = _RAND_8[3:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    FPToInt_cov[initvar] = _RAND_9[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  FPToInt_covSum = _RAND_10[29:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      in_ren2 <= 1'h0;
    end else if (io_in_valid) begin
      in_ren2 <= io_in_bits_ren2;
    end
    if (metaReset) begin
      in_typeTagOut <= 2'h0;
    end else if (io_in_valid) begin
      in_typeTagOut <= io_in_bits_typeTagOut;
    end
    if (metaReset) begin
      in_wflags <= 1'h0;
    end else if (io_in_valid) begin
      in_wflags <= io_in_bits_wflags;
    end
    if (metaReset) begin
      in_rm <= 3'h0;
    end else if (io_in_valid) begin
      in_rm <= io_in_bits_rm;
    end
    if (metaReset) begin
      in_typ <= 2'h0;
    end else if (io_in_valid) begin
      in_typ <= io_in_bits_typ;
    end
    if (metaReset) begin
      in_fmt <= 2'h0;
    end else if (io_in_valid) begin
      in_fmt <= io_in_bits_fmt;
    end
    if (metaReset) begin
      in_in1 <= 65'h0;
    end else if (io_in_valid) begin
      in_in1 <= io_in_bits_in1;
    end
    if (metaReset) begin
      in_in2 <= 65'h0;
    end else if (io_in_valid) begin
      in_in2 <= io_in_bits_in2;
    end
    FPToInt_state <= FPToInt_xor0;
    if (!(FPToInt_cov_read_data)) begin
      FPToInt_covSum <= FPToInt_covSum + 1'h1;
    end
  end
  always @(posedge clock) begin
    if(FPToInt_cov_write_en & FPToInt_cov_write_mask) begin
      FPToInt_cov[FPToInt_cov_write_addr] <= FPToInt_cov_write_data; // @[Coverage map for FPToInt]
    end
  end
endmodule
module IntToFP(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [1:0]  io_in_bits_typeTagIn,
  input         io_in_bits_wflags,
  input  [2:0]  io_in_bits_rm,
  input  [1:0]  io_in_bits_typ,
  input  [63:0] io_in_bits_in1,
  output [64:0] io_out_bits_data,
  output [4:0]  io_out_bits_exc,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  wire  i2f_io_signedIn; // @[FPU.scala 551:23]
  wire [63:0] i2f_io_in; // @[FPU.scala 551:23]
  wire [2:0] i2f_io_roundingMode; // @[FPU.scala 551:23]
  wire [32:0] i2f_io_out; // @[FPU.scala 551:23]
  wire [4:0] i2f_io_exceptionFlags; // @[FPU.scala 551:23]
  wire [29:0] i2f_io_covSum; // @[FPU.scala 551:23]
  wire  i2f_metaAssert; // @[FPU.scala 551:23]
  wire  i2f_1_io_signedIn; // @[FPU.scala 551:23]
  wire [63:0] i2f_1_io_in; // @[FPU.scala 551:23]
  wire [2:0] i2f_1_io_roundingMode; // @[FPU.scala 551:23]
  wire [64:0] i2f_1_io_out; // @[FPU.scala 551:23]
  wire [4:0] i2f_1_io_exceptionFlags; // @[FPU.scala 551:23]
  wire [29:0] i2f_1_io_covSum; // @[FPU.scala 551:23]
  wire  i2f_1_metaAssert; // @[FPU.scala 551:23]
  reg  inPipe_valid; // @[Valid.scala 117:22]
  reg [31:0] _RAND_0;
  reg [1:0] inPipe_bits_typeTagIn; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  reg  inPipe_bits_wflags; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [2:0] inPipe_bits_rm; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg [1:0] inPipe_bits_typ; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg [63:0] inPipe_bits_in1; // @[Reg.scala 15:16]
  reg [63:0] _RAND_5;
  wire  mux_data_truncIdx; // @[package.scala 31:49]
  wire [63:0] _mux_data_T_1; // @[package.scala 32:76]
  wire [63:0] _mux_data_T_2; // @[FPU.scala 426:23]
  wire  mux_data_rawIn_sign; // @[rawFloatFromFN.scala 46:22]
  wire [10:0] mux_data_rawIn_expIn; // @[rawFloatFromFN.scala 47:23]
  wire [51:0] mux_data_rawIn_fractIn; // @[rawFloatFromFN.scala 48:25]
  wire  mux_data_rawIn_isZeroExpIn; // @[rawFloatFromFN.scala 50:34]
  wire  mux_data_rawIn_isZeroFractIn; // @[rawFloatFromFN.scala 51:38]
  wire [5:0] _mux_data_rawIn_normDist_T_52; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_53; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_54; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_55; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_56; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_57; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_58; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_59; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_60; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_61; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_62; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_63; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_64; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_65; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_66; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_67; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_68; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_69; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_70; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_71; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_72; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_73; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_74; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_75; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_76; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_77; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_78; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_79; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_80; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_81; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_82; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_83; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_84; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_85; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_86; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_87; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_88; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_89; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_90; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_91; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_92; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_93; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_94; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_95; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_96; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_97; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_98; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_99; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_100; // @[Mux.scala 47:69]
  wire [5:0] _mux_data_rawIn_normDist_T_101; // @[Mux.scala 47:69]
  wire [5:0] mux_data_rawIn_normDist; // @[Mux.scala 47:69]
  wire [114:0] _GEN_24; // @[rawFloatFromFN.scala 54:36]
  wire [114:0] _mux_data_rawIn_subnormFract_T; // @[rawFloatFromFN.scala 54:36]
  wire [51:0] mux_data_rawIn_subnormFract; // @[rawFloatFromFN.scala 54:64]
  wire [11:0] _GEN_25; // @[rawFloatFromFN.scala 57:26]
  wire [11:0] _mux_data_rawIn_adjustedExp_T; // @[rawFloatFromFN.scala 57:26]
  wire [11:0] _mux_data_rawIn_adjustedExp_T_1; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _mux_data_rawIn_adjustedExp_T_2; // @[rawFloatFromFN.scala 60:27]
  wire [10:0] _GEN_26; // @[rawFloatFromFN.scala 60:22]
  wire [10:0] _mux_data_rawIn_adjustedExp_T_3; // @[rawFloatFromFN.scala 60:22]
  wire [11:0] _GEN_27; // @[rawFloatFromFN.scala 59:15]
  wire [11:0] mux_data_rawIn_adjustedExp; // @[rawFloatFromFN.scala 59:15]
  wire  mux_data_rawIn_isZero; // @[rawFloatFromFN.scala 62:34]
  wire  mux_data_rawIn_isSpecial; // @[rawFloatFromFN.scala 63:62]
  wire  mux_data_rawIn__isNaN; // @[rawFloatFromFN.scala 66:33]
  wire [12:0] mux_data_rawIn__sExp; // @[rawFloatFromFN.scala 70:48]
  wire  mux_data_rawIn_out_sig_hi_lo; // @[rawFloatFromFN.scala 72:29]
  wire [51:0] mux_data_rawIn_out_sig_lo; // @[rawFloatFromFN.scala 72:42]
  wire [53:0] mux_data_rawIn__sig; // @[Cat.scala 30:58]
  wire [2:0] _mux_data_T_4; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_28; // @[recFNFromFN.scala 48:79]
  wire [2:0] mux_data_hi_lo; // @[recFNFromFN.scala 48:79]
  wire [8:0] mux_data_lo_hi; // @[recFNFromFN.scala 50:23]
  wire [51:0] mux_data_lo_lo; // @[recFNFromFN.scala 51:22]
  wire [64:0] _mux_data_T_6; // @[Cat.scala 30:58]
  wire  mux_data_rawIn_sign_1; // @[rawFloatFromFN.scala 46:22]
  wire [7:0] mux_data_rawIn_expIn_1; // @[rawFloatFromFN.scala 47:23]
  wire [22:0] mux_data_rawIn_fractIn_1; // @[rawFloatFromFN.scala 48:25]
  wire  mux_data_rawIn_isZeroExpIn_1; // @[rawFloatFromFN.scala 50:34]
  wire  mux_data_rawIn_isZeroFractIn_1; // @[rawFloatFromFN.scala 51:38]
  wire [4:0] _mux_data_rawIn_normDist_T_125; // @[Mux.scala 47:69]
  wire [4:0] _mux_data_rawIn_normDist_T_126; // @[Mux.scala 47:69]
  wire [4:0] _mux_data_rawIn_normDist_T_127; // @[Mux.scala 47:69]
  wire [4:0] _mux_data_rawIn_normDist_T_128; // @[Mux.scala 47:69]
  wire [4:0] _mux_data_rawIn_normDist_T_129; // @[Mux.scala 47:69]
  wire [4:0] _mux_data_rawIn_normDist_T_130; // @[Mux.scala 47:69]
  wire [4:0] _mux_data_rawIn_normDist_T_131; // @[Mux.scala 47:69]
  wire [4:0] _mux_data_rawIn_normDist_T_132; // @[Mux.scala 47:69]
  wire [4:0] _mux_data_rawIn_normDist_T_133; // @[Mux.scala 47:69]
  wire [4:0] _mux_data_rawIn_normDist_T_134; // @[Mux.scala 47:69]
  wire [4:0] _mux_data_rawIn_normDist_T_135; // @[Mux.scala 47:69]
  wire [4:0] _mux_data_rawIn_normDist_T_136; // @[Mux.scala 47:69]
  wire [4:0] _mux_data_rawIn_normDist_T_137; // @[Mux.scala 47:69]
  wire [4:0] _mux_data_rawIn_normDist_T_138; // @[Mux.scala 47:69]
  wire [4:0] _mux_data_rawIn_normDist_T_139; // @[Mux.scala 47:69]
  wire [4:0] _mux_data_rawIn_normDist_T_140; // @[Mux.scala 47:69]
  wire [4:0] _mux_data_rawIn_normDist_T_141; // @[Mux.scala 47:69]
  wire [4:0] _mux_data_rawIn_normDist_T_142; // @[Mux.scala 47:69]
  wire [4:0] _mux_data_rawIn_normDist_T_143; // @[Mux.scala 47:69]
  wire [4:0] _mux_data_rawIn_normDist_T_144; // @[Mux.scala 47:69]
  wire [4:0] _mux_data_rawIn_normDist_T_145; // @[Mux.scala 47:69]
  wire [4:0] mux_data_rawIn_normDist_1; // @[Mux.scala 47:69]
  wire [53:0] _GEN_29; // @[rawFloatFromFN.scala 54:36]
  wire [53:0] _mux_data_rawIn_subnormFract_T_2; // @[rawFloatFromFN.scala 54:36]
  wire [22:0] mux_data_rawIn_subnormFract_1; // @[rawFloatFromFN.scala 54:64]
  wire [8:0] _GEN_30; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _mux_data_rawIn_adjustedExp_T_5; // @[rawFloatFromFN.scala 57:26]
  wire [8:0] _mux_data_rawIn_adjustedExp_T_6; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _mux_data_rawIn_adjustedExp_T_7; // @[rawFloatFromFN.scala 60:27]
  wire [7:0] _GEN_31; // @[rawFloatFromFN.scala 60:22]
  wire [7:0] _mux_data_rawIn_adjustedExp_T_8; // @[rawFloatFromFN.scala 60:22]
  wire [8:0] _GEN_32; // @[rawFloatFromFN.scala 59:15]
  wire [8:0] mux_data_rawIn_adjustedExp_1; // @[rawFloatFromFN.scala 59:15]
  wire  mux_data_rawIn_isZero_1; // @[rawFloatFromFN.scala 62:34]
  wire  mux_data_rawIn_isSpecial_1; // @[rawFloatFromFN.scala 63:62]
  wire  mux_data_rawIn_1_isNaN; // @[rawFloatFromFN.scala 66:33]
  wire [9:0] mux_data_rawIn_1_sExp; // @[rawFloatFromFN.scala 70:48]
  wire  mux_data_rawIn_out_sig_hi_lo_1; // @[rawFloatFromFN.scala 72:29]
  wire [22:0] mux_data_rawIn_out_sig_lo_1; // @[rawFloatFromFN.scala 72:42]
  wire [24:0] mux_data_rawIn_1_sig; // @[Cat.scala 30:58]
  wire [2:0] _mux_data_T_8; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_33; // @[recFNFromFN.scala 48:79]
  wire [2:0] mux_data_hi_lo_1; // @[recFNFromFN.scala 48:79]
  wire [5:0] mux_data_lo_hi_1; // @[recFNFromFN.scala 50:23]
  wire [22:0] mux_data_lo_lo_1; // @[recFNFromFN.scala 51:22]
  wire [32:0] _mux_data_T_10; // @[Cat.scala 30:58]
  wire [3:0] mux_data_swizzledNaN_hi_hi_hi; // @[FPU.scala 332:8]
  wire  mux_data_swizzledNaN_hi_hi_lo; // @[FPU.scala 333:42]
  wire [6:0] mux_data_swizzledNaN_hi_lo_hi; // @[FPU.scala 334:8]
  wire  mux_data_swizzledNaN_hi_lo_lo; // @[FPU.scala 335:8]
  wire  mux_data_swizzledNaN_lo_hi_lo; // @[FPU.scala 337:8]
  wire [30:0] mux_data_swizzledNaN_lo_lo; // @[FPU.scala 338:8]
  wire [64:0] mux_data_swizzledNaN; // @[Cat.scala 30:58]
  wire  _mux_data_T_12; // @[FPU.scala 243:56]
  wire [31:0] intValue_smallInt; // @[FPU.scala 539:33]
  wire [32:0] _intValue_res_T_1; // @[FPU.scala 541:45]
  wire [31:0] _intValue_res_T_2; // @[FPU.scala 541:60]
  wire [32:0] _intValue_res_T_3; // @[FPU.scala 541:19]
  wire [64:0] maskedNaN; // @[FPU.scala 408:25]
  wire  _T_1; // @[FPU.scala 243:56]
  wire [64:0] _T_2; // @[FPU.scala 409:10]
  wire [31:0] dataPadded_hi; // @[FPU.scala 560:55]
  wire [64:0] dataPadded_0; // @[Cat.scala 30:58]
  reg [64:0] io_out_b_data; // @[Reg.scala 15:16]
  reg [95:0] _RAND_6;
  reg [4:0] io_out_b_exc; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7;
  reg [3:0] IntToFP_state; // @[Register tracking IntToFP state]
  reg [31:0] _RAND_8;
  reg  IntToFP_cov [0:15]; // @[Coverage map for IntToFP]
  reg [31:0] _RAND_9;
  wire  IntToFP_cov_read_data; // @[Coverage map for IntToFP]
  wire [3:0] IntToFP_cov_read_addr; // @[Coverage map for IntToFP]
  wire  IntToFP_cov_write_data; // @[Coverage map for IntToFP]
  wire [3:0] IntToFP_cov_write_addr; // @[Coverage map for IntToFP]
  wire  IntToFP_cov_write_mask; // @[Coverage map for IntToFP]
  wire  IntToFP_cov_write_en; // @[Coverage map for IntToFP]
  reg [29:0] IntToFP_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_10;
  wire  inPipe_valid_shl;
  wire [3:0] inPipe_valid_pad;
  wire [1:0] inPipe_bits_wflags_shl;
  wire [3:0] inPipe_bits_wflags_pad;
  wire [3:0] inPipe_bits_typ_shl;
  wire [3:0] inPipe_bits_typ_pad;
  wire [3:0] IntToFP_xor2;
  wire [3:0] IntToFP_xor0;
  wire [29:0] i2f_sum;
  wire [29:0] i2f_1_sum;
  wire  i2f_metaAssert_wire;
  wire  i2f_1_metaAssert_wire;
  wire  IntToFP_or0;
  reg  IntToFP_metaAssert;
  reg [31:0] _RAND_11;
  INToRecFN i2f ( // @[FPU.scala 551:23]
    .io_signedIn(i2f_io_signedIn),
    .io_in(i2f_io_in),
    .io_roundingMode(i2f_io_roundingMode),
    .io_out(i2f_io_out),
    .io_exceptionFlags(i2f_io_exceptionFlags),
    .io_covSum(i2f_io_covSum),
    .metaAssert(i2f_metaAssert)
  );
  INToRecFN_1 i2f_1 ( // @[FPU.scala 551:23]
    .io_signedIn(i2f_1_io_signedIn),
    .io_in(i2f_1_io_in),
    .io_roundingMode(i2f_1_io_roundingMode),
    .io_out(i2f_1_io_out),
    .io_exceptionFlags(i2f_1_io_exceptionFlags),
    .io_covSum(i2f_1_io_covSum),
    .metaAssert(i2f_1_metaAssert)
  );
  assign mux_data_truncIdx = inPipe_bits_typeTagIn[0]; // @[package.scala 31:49]
  assign _mux_data_T_1 = mux_data_truncIdx ? 64'h0 : 64'hffffffff00000000; // @[package.scala 32:76]
  assign _mux_data_T_2 = _mux_data_T_1 | inPipe_bits_in1; // @[FPU.scala 426:23]
  assign mux_data_rawIn_sign = _mux_data_T_2[63]; // @[rawFloatFromFN.scala 46:22]
  assign mux_data_rawIn_expIn = _mux_data_T_2[62:52]; // @[rawFloatFromFN.scala 47:23]
  assign mux_data_rawIn_fractIn = _mux_data_T_2[51:0]; // @[rawFloatFromFN.scala 48:25]
  assign mux_data_rawIn_isZeroExpIn = mux_data_rawIn_expIn == 11'h0; // @[rawFloatFromFN.scala 50:34]
  assign mux_data_rawIn_isZeroFractIn = mux_data_rawIn_fractIn == 52'h0; // @[rawFloatFromFN.scala 51:38]
  assign _mux_data_rawIn_normDist_T_52 = mux_data_rawIn_fractIn[1] ? 6'h32 : 6'h33; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_53 = mux_data_rawIn_fractIn[2] ? 6'h31 : _mux_data_rawIn_normDist_T_52; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_54 = mux_data_rawIn_fractIn[3] ? 6'h30 : _mux_data_rawIn_normDist_T_53; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_55 = mux_data_rawIn_fractIn[4] ? 6'h2f : _mux_data_rawIn_normDist_T_54; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_56 = mux_data_rawIn_fractIn[5] ? 6'h2e : _mux_data_rawIn_normDist_T_55; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_57 = mux_data_rawIn_fractIn[6] ? 6'h2d : _mux_data_rawIn_normDist_T_56; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_58 = mux_data_rawIn_fractIn[7] ? 6'h2c : _mux_data_rawIn_normDist_T_57; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_59 = mux_data_rawIn_fractIn[8] ? 6'h2b : _mux_data_rawIn_normDist_T_58; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_60 = mux_data_rawIn_fractIn[9] ? 6'h2a : _mux_data_rawIn_normDist_T_59; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_61 = mux_data_rawIn_fractIn[10] ? 6'h29 : _mux_data_rawIn_normDist_T_60; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_62 = mux_data_rawIn_fractIn[11] ? 6'h28 : _mux_data_rawIn_normDist_T_61; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_63 = mux_data_rawIn_fractIn[12] ? 6'h27 : _mux_data_rawIn_normDist_T_62; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_64 = mux_data_rawIn_fractIn[13] ? 6'h26 : _mux_data_rawIn_normDist_T_63; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_65 = mux_data_rawIn_fractIn[14] ? 6'h25 : _mux_data_rawIn_normDist_T_64; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_66 = mux_data_rawIn_fractIn[15] ? 6'h24 : _mux_data_rawIn_normDist_T_65; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_67 = mux_data_rawIn_fractIn[16] ? 6'h23 : _mux_data_rawIn_normDist_T_66; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_68 = mux_data_rawIn_fractIn[17] ? 6'h22 : _mux_data_rawIn_normDist_T_67; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_69 = mux_data_rawIn_fractIn[18] ? 6'h21 : _mux_data_rawIn_normDist_T_68; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_70 = mux_data_rawIn_fractIn[19] ? 6'h20 : _mux_data_rawIn_normDist_T_69; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_71 = mux_data_rawIn_fractIn[20] ? 6'h1f : _mux_data_rawIn_normDist_T_70; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_72 = mux_data_rawIn_fractIn[21] ? 6'h1e : _mux_data_rawIn_normDist_T_71; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_73 = mux_data_rawIn_fractIn[22] ? 6'h1d : _mux_data_rawIn_normDist_T_72; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_74 = mux_data_rawIn_fractIn[23] ? 6'h1c : _mux_data_rawIn_normDist_T_73; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_75 = mux_data_rawIn_fractIn[24] ? 6'h1b : _mux_data_rawIn_normDist_T_74; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_76 = mux_data_rawIn_fractIn[25] ? 6'h1a : _mux_data_rawIn_normDist_T_75; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_77 = mux_data_rawIn_fractIn[26] ? 6'h19 : _mux_data_rawIn_normDist_T_76; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_78 = mux_data_rawIn_fractIn[27] ? 6'h18 : _mux_data_rawIn_normDist_T_77; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_79 = mux_data_rawIn_fractIn[28] ? 6'h17 : _mux_data_rawIn_normDist_T_78; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_80 = mux_data_rawIn_fractIn[29] ? 6'h16 : _mux_data_rawIn_normDist_T_79; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_81 = mux_data_rawIn_fractIn[30] ? 6'h15 : _mux_data_rawIn_normDist_T_80; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_82 = mux_data_rawIn_fractIn[31] ? 6'h14 : _mux_data_rawIn_normDist_T_81; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_83 = mux_data_rawIn_fractIn[32] ? 6'h13 : _mux_data_rawIn_normDist_T_82; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_84 = mux_data_rawIn_fractIn[33] ? 6'h12 : _mux_data_rawIn_normDist_T_83; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_85 = mux_data_rawIn_fractIn[34] ? 6'h11 : _mux_data_rawIn_normDist_T_84; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_86 = mux_data_rawIn_fractIn[35] ? 6'h10 : _mux_data_rawIn_normDist_T_85; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_87 = mux_data_rawIn_fractIn[36] ? 6'hf : _mux_data_rawIn_normDist_T_86; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_88 = mux_data_rawIn_fractIn[37] ? 6'he : _mux_data_rawIn_normDist_T_87; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_89 = mux_data_rawIn_fractIn[38] ? 6'hd : _mux_data_rawIn_normDist_T_88; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_90 = mux_data_rawIn_fractIn[39] ? 6'hc : _mux_data_rawIn_normDist_T_89; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_91 = mux_data_rawIn_fractIn[40] ? 6'hb : _mux_data_rawIn_normDist_T_90; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_92 = mux_data_rawIn_fractIn[41] ? 6'ha : _mux_data_rawIn_normDist_T_91; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_93 = mux_data_rawIn_fractIn[42] ? 6'h9 : _mux_data_rawIn_normDist_T_92; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_94 = mux_data_rawIn_fractIn[43] ? 6'h8 : _mux_data_rawIn_normDist_T_93; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_95 = mux_data_rawIn_fractIn[44] ? 6'h7 : _mux_data_rawIn_normDist_T_94; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_96 = mux_data_rawIn_fractIn[45] ? 6'h6 : _mux_data_rawIn_normDist_T_95; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_97 = mux_data_rawIn_fractIn[46] ? 6'h5 : _mux_data_rawIn_normDist_T_96; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_98 = mux_data_rawIn_fractIn[47] ? 6'h4 : _mux_data_rawIn_normDist_T_97; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_99 = mux_data_rawIn_fractIn[48] ? 6'h3 : _mux_data_rawIn_normDist_T_98; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_100 = mux_data_rawIn_fractIn[49] ? 6'h2 : _mux_data_rawIn_normDist_T_99; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_101 = mux_data_rawIn_fractIn[50] ? 6'h1 : _mux_data_rawIn_normDist_T_100; // @[Mux.scala 47:69]
  assign mux_data_rawIn_normDist = mux_data_rawIn_fractIn[51] ? 6'h0 : _mux_data_rawIn_normDist_T_101; // @[Mux.scala 47:69]
  assign _GEN_24 = {{63'd0}, mux_data_rawIn_fractIn}; // @[rawFloatFromFN.scala 54:36]
  assign _mux_data_rawIn_subnormFract_T = _GEN_24 << mux_data_rawIn_normDist; // @[rawFloatFromFN.scala 54:36]
  assign mux_data_rawIn_subnormFract = {_mux_data_rawIn_subnormFract_T[50:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  assign _GEN_25 = {{6'd0}, mux_data_rawIn_normDist}; // @[rawFloatFromFN.scala 57:26]
  assign _mux_data_rawIn_adjustedExp_T = _GEN_25 ^ 12'hfff; // @[rawFloatFromFN.scala 57:26]
  assign _mux_data_rawIn_adjustedExp_T_1 = mux_data_rawIn_isZeroExpIn ? _mux_data_rawIn_adjustedExp_T : {{1'd0}, mux_data_rawIn_expIn}; // @[rawFloatFromFN.scala 56:16]
  assign _mux_data_rawIn_adjustedExp_T_2 = mux_data_rawIn_isZeroExpIn ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  assign _GEN_26 = {{9'd0}, _mux_data_rawIn_adjustedExp_T_2}; // @[rawFloatFromFN.scala 60:22]
  assign _mux_data_rawIn_adjustedExp_T_3 = 11'h400 | _GEN_26; // @[rawFloatFromFN.scala 60:22]
  assign _GEN_27 = {{1'd0}, _mux_data_rawIn_adjustedExp_T_3}; // @[rawFloatFromFN.scala 59:15]
  assign mux_data_rawIn_adjustedExp = _mux_data_rawIn_adjustedExp_T_1 + _GEN_27; // @[rawFloatFromFN.scala 59:15]
  assign mux_data_rawIn_isZero = mux_data_rawIn_isZeroExpIn & mux_data_rawIn_isZeroFractIn; // @[rawFloatFromFN.scala 62:34]
  assign mux_data_rawIn_isSpecial = mux_data_rawIn_adjustedExp[11:10] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  assign mux_data_rawIn__isNaN = mux_data_rawIn_isSpecial & ~mux_data_rawIn_isZeroFractIn; // @[rawFloatFromFN.scala 66:33]
  assign mux_data_rawIn__sExp = {1'b0,$signed(mux_data_rawIn_adjustedExp)}; // @[rawFloatFromFN.scala 70:48]
  assign mux_data_rawIn_out_sig_hi_lo = ~mux_data_rawIn_isZero; // @[rawFloatFromFN.scala 72:29]
  assign mux_data_rawIn_out_sig_lo = mux_data_rawIn_isZeroExpIn ? mux_data_rawIn_subnormFract : mux_data_rawIn_fractIn; // @[rawFloatFromFN.scala 72:42]
  assign mux_data_rawIn__sig = {1'h0,mux_data_rawIn_out_sig_hi_lo,mux_data_rawIn_out_sig_lo}; // @[Cat.scala 30:58]
  assign _mux_data_T_4 = mux_data_rawIn_isZero ? 3'h0 : mux_data_rawIn__sExp[11:9]; // @[recFNFromFN.scala 48:16]
  assign _GEN_28 = {{2'd0}, mux_data_rawIn__isNaN}; // @[recFNFromFN.scala 48:79]
  assign mux_data_hi_lo = _mux_data_T_4 | _GEN_28; // @[recFNFromFN.scala 48:79]
  assign mux_data_lo_hi = mux_data_rawIn__sExp[8:0]; // @[recFNFromFN.scala 50:23]
  assign mux_data_lo_lo = mux_data_rawIn__sig[51:0]; // @[recFNFromFN.scala 51:22]
  assign _mux_data_T_6 = {mux_data_rawIn_sign,mux_data_hi_lo,mux_data_lo_hi,mux_data_lo_lo}; // @[Cat.scala 30:58]
  assign mux_data_rawIn_sign_1 = _mux_data_T_2[31]; // @[rawFloatFromFN.scala 46:22]
  assign mux_data_rawIn_expIn_1 = _mux_data_T_2[30:23]; // @[rawFloatFromFN.scala 47:23]
  assign mux_data_rawIn_fractIn_1 = _mux_data_T_2[22:0]; // @[rawFloatFromFN.scala 48:25]
  assign mux_data_rawIn_isZeroExpIn_1 = mux_data_rawIn_expIn_1 == 8'h0; // @[rawFloatFromFN.scala 50:34]
  assign mux_data_rawIn_isZeroFractIn_1 = mux_data_rawIn_fractIn_1 == 23'h0; // @[rawFloatFromFN.scala 51:38]
  assign _mux_data_rawIn_normDist_T_125 = mux_data_rawIn_fractIn_1[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_126 = mux_data_rawIn_fractIn_1[2] ? 5'h14 : _mux_data_rawIn_normDist_T_125; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_127 = mux_data_rawIn_fractIn_1[3] ? 5'h13 : _mux_data_rawIn_normDist_T_126; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_128 = mux_data_rawIn_fractIn_1[4] ? 5'h12 : _mux_data_rawIn_normDist_T_127; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_129 = mux_data_rawIn_fractIn_1[5] ? 5'h11 : _mux_data_rawIn_normDist_T_128; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_130 = mux_data_rawIn_fractIn_1[6] ? 5'h10 : _mux_data_rawIn_normDist_T_129; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_131 = mux_data_rawIn_fractIn_1[7] ? 5'hf : _mux_data_rawIn_normDist_T_130; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_132 = mux_data_rawIn_fractIn_1[8] ? 5'he : _mux_data_rawIn_normDist_T_131; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_133 = mux_data_rawIn_fractIn_1[9] ? 5'hd : _mux_data_rawIn_normDist_T_132; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_134 = mux_data_rawIn_fractIn_1[10] ? 5'hc : _mux_data_rawIn_normDist_T_133; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_135 = mux_data_rawIn_fractIn_1[11] ? 5'hb : _mux_data_rawIn_normDist_T_134; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_136 = mux_data_rawIn_fractIn_1[12] ? 5'ha : _mux_data_rawIn_normDist_T_135; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_137 = mux_data_rawIn_fractIn_1[13] ? 5'h9 : _mux_data_rawIn_normDist_T_136; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_138 = mux_data_rawIn_fractIn_1[14] ? 5'h8 : _mux_data_rawIn_normDist_T_137; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_139 = mux_data_rawIn_fractIn_1[15] ? 5'h7 : _mux_data_rawIn_normDist_T_138; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_140 = mux_data_rawIn_fractIn_1[16] ? 5'h6 : _mux_data_rawIn_normDist_T_139; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_141 = mux_data_rawIn_fractIn_1[17] ? 5'h5 : _mux_data_rawIn_normDist_T_140; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_142 = mux_data_rawIn_fractIn_1[18] ? 5'h4 : _mux_data_rawIn_normDist_T_141; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_143 = mux_data_rawIn_fractIn_1[19] ? 5'h3 : _mux_data_rawIn_normDist_T_142; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_144 = mux_data_rawIn_fractIn_1[20] ? 5'h2 : _mux_data_rawIn_normDist_T_143; // @[Mux.scala 47:69]
  assign _mux_data_rawIn_normDist_T_145 = mux_data_rawIn_fractIn_1[21] ? 5'h1 : _mux_data_rawIn_normDist_T_144; // @[Mux.scala 47:69]
  assign mux_data_rawIn_normDist_1 = mux_data_rawIn_fractIn_1[22] ? 5'h0 : _mux_data_rawIn_normDist_T_145; // @[Mux.scala 47:69]
  assign _GEN_29 = {{31'd0}, mux_data_rawIn_fractIn_1}; // @[rawFloatFromFN.scala 54:36]
  assign _mux_data_rawIn_subnormFract_T_2 = _GEN_29 << mux_data_rawIn_normDist_1; // @[rawFloatFromFN.scala 54:36]
  assign mux_data_rawIn_subnormFract_1 = {_mux_data_rawIn_subnormFract_T_2[21:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  assign _GEN_30 = {{4'd0}, mux_data_rawIn_normDist_1}; // @[rawFloatFromFN.scala 57:26]
  assign _mux_data_rawIn_adjustedExp_T_5 = _GEN_30 ^ 9'h1ff; // @[rawFloatFromFN.scala 57:26]
  assign _mux_data_rawIn_adjustedExp_T_6 = mux_data_rawIn_isZeroExpIn_1 ? _mux_data_rawIn_adjustedExp_T_5 : {{1'd0}, mux_data_rawIn_expIn_1}; // @[rawFloatFromFN.scala 56:16]
  assign _mux_data_rawIn_adjustedExp_T_7 = mux_data_rawIn_isZeroExpIn_1 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  assign _GEN_31 = {{6'd0}, _mux_data_rawIn_adjustedExp_T_7}; // @[rawFloatFromFN.scala 60:22]
  assign _mux_data_rawIn_adjustedExp_T_8 = 8'h80 | _GEN_31; // @[rawFloatFromFN.scala 60:22]
  assign _GEN_32 = {{1'd0}, _mux_data_rawIn_adjustedExp_T_8}; // @[rawFloatFromFN.scala 59:15]
  assign mux_data_rawIn_adjustedExp_1 = _mux_data_rawIn_adjustedExp_T_6 + _GEN_32; // @[rawFloatFromFN.scala 59:15]
  assign mux_data_rawIn_isZero_1 = mux_data_rawIn_isZeroExpIn_1 & mux_data_rawIn_isZeroFractIn_1; // @[rawFloatFromFN.scala 62:34]
  assign mux_data_rawIn_isSpecial_1 = mux_data_rawIn_adjustedExp_1[8:7] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  assign mux_data_rawIn_1_isNaN = mux_data_rawIn_isSpecial_1 & ~mux_data_rawIn_isZeroFractIn_1; // @[rawFloatFromFN.scala 66:33]
  assign mux_data_rawIn_1_sExp = {1'b0,$signed(mux_data_rawIn_adjustedExp_1)}; // @[rawFloatFromFN.scala 70:48]
  assign mux_data_rawIn_out_sig_hi_lo_1 = ~mux_data_rawIn_isZero_1; // @[rawFloatFromFN.scala 72:29]
  assign mux_data_rawIn_out_sig_lo_1 = mux_data_rawIn_isZeroExpIn_1 ? mux_data_rawIn_subnormFract_1 : mux_data_rawIn_fractIn_1; // @[rawFloatFromFN.scala 72:42]
  assign mux_data_rawIn_1_sig = {1'h0,mux_data_rawIn_out_sig_hi_lo_1,mux_data_rawIn_out_sig_lo_1}; // @[Cat.scala 30:58]
  assign _mux_data_T_8 = mux_data_rawIn_isZero_1 ? 3'h0 : mux_data_rawIn_1_sExp[8:6]; // @[recFNFromFN.scala 48:16]
  assign _GEN_33 = {{2'd0}, mux_data_rawIn_1_isNaN}; // @[recFNFromFN.scala 48:79]
  assign mux_data_hi_lo_1 = _mux_data_T_8 | _GEN_33; // @[recFNFromFN.scala 48:79]
  assign mux_data_lo_hi_1 = mux_data_rawIn_1_sExp[5:0]; // @[recFNFromFN.scala 50:23]
  assign mux_data_lo_lo_1 = mux_data_rawIn_1_sig[22:0]; // @[recFNFromFN.scala 51:22]
  assign _mux_data_T_10 = {mux_data_rawIn_sign_1,mux_data_hi_lo_1,mux_data_lo_hi_1,mux_data_lo_lo_1}; // @[Cat.scala 30:58]
  assign mux_data_swizzledNaN_hi_hi_hi = _mux_data_T_6[64:61]; // @[FPU.scala 332:8]
  assign mux_data_swizzledNaN_hi_hi_lo = &_mux_data_T_6[51:32]; // @[FPU.scala 333:42]
  assign mux_data_swizzledNaN_hi_lo_hi = _mux_data_T_6[59:53]; // @[FPU.scala 334:8]
  assign mux_data_swizzledNaN_hi_lo_lo = _mux_data_T_10[31]; // @[FPU.scala 335:8]
  assign mux_data_swizzledNaN_lo_hi_lo = _mux_data_T_10[32]; // @[FPU.scala 337:8]
  assign mux_data_swizzledNaN_lo_lo = _mux_data_T_10[30:0]; // @[FPU.scala 338:8]
  assign mux_data_swizzledNaN = {mux_data_swizzledNaN_hi_hi_hi,mux_data_swizzledNaN_hi_hi_lo,mux_data_swizzledNaN_hi_lo_hi,mux_data_swizzledNaN_hi_lo_lo,_mux_data_T_6[51:32],mux_data_swizzledNaN_lo_hi_lo,mux_data_swizzledNaN_lo_lo}; // @[Cat.scala 30:58]
  assign _mux_data_T_12 = &_mux_data_T_6[63:61]; // @[FPU.scala 243:56]
  assign intValue_smallInt = inPipe_bits_in1[31:0]; // @[FPU.scala 539:33]
  assign _intValue_res_T_1 = {1'b0,$signed(intValue_smallInt)}; // @[FPU.scala 541:45]
  assign _intValue_res_T_2 = inPipe_bits_in1[31:0]; // @[FPU.scala 541:60]
  assign _intValue_res_T_3 = inPipe_bits_typ[0] ? $signed(_intValue_res_T_1) : $signed({{1{_intValue_res_T_2[31]}},_intValue_res_T_2}); // @[FPU.scala 541:19]
  assign maskedNaN = i2f_1_io_out & 65'h1efefffffffffffff; // @[FPU.scala 408:25]
  assign _T_1 = &i2f_1_io_out[63:61]; // @[FPU.scala 243:56]
  assign _T_2 = _T_1 ? maskedNaN : i2f_1_io_out; // @[FPU.scala 409:10]
  assign dataPadded_hi = _T_2[64:33]; // @[FPU.scala 560:55]
  assign dataPadded_0 = {dataPadded_hi,i2f_io_out}; // @[Cat.scala 30:58]
  assign io_out_bits_data = io_out_b_data; // @[FPU.scala 565:10]
  assign io_out_bits_exc = io_out_b_exc; // @[FPU.scala 565:10]
  assign i2f_io_signedIn = ~inPipe_bits_typ[0]; // @[FPU.scala 552:23]
  assign i2f_io_in = inPipe_bits_typ[1] ? $signed(inPipe_bits_in1) : $signed({{31{_intValue_res_T_3[32]}},_intValue_res_T_3}); // @[FPU.scala 553:17]
  assign i2f_io_roundingMode = inPipe_bits_rm; // @[FPU.scala 554:27]
  assign i2f_1_io_signedIn = ~inPipe_bits_typ[0]; // @[FPU.scala 552:23]
  assign i2f_1_io_in = inPipe_bits_typ[1] ? $signed(inPipe_bits_in1) : $signed({{31{_intValue_res_T_3[32]}},_intValue_res_T_3}); // @[FPU.scala 553:17]
  assign i2f_1_io_roundingMode = inPipe_bits_rm; // @[FPU.scala 554:27]
  assign IntToFP_cov_read_addr = IntToFP_state;
  assign IntToFP_cov_read_data = IntToFP_cov[IntToFP_cov_read_addr]; // @[Coverage map for IntToFP]
  assign IntToFP_cov_write_data = 1'h1;
  assign IntToFP_cov_write_addr = IntToFP_state;
  assign IntToFP_cov_write_mask = 1'h1;
  assign IntToFP_cov_write_en = 1'h1;
  assign inPipe_valid_shl = inPipe_valid;
  assign inPipe_valid_pad = {3'h0,inPipe_valid_shl};
  assign inPipe_bits_wflags_shl = {inPipe_bits_wflags, 1'h0};
  assign inPipe_bits_wflags_pad = {2'h0,inPipe_bits_wflags_shl};
  assign inPipe_bits_typ_shl = {inPipe_bits_typ, 2'h0};
  assign inPipe_bits_typ_pad = inPipe_bits_typ_shl;
  assign IntToFP_xor2 = inPipe_bits_wflags_pad ^ inPipe_bits_typ_pad;
  assign IntToFP_xor0 = inPipe_valid_pad ^ IntToFP_xor2;
  assign i2f_sum = IntToFP_covSum + i2f_io_covSum;
  assign i2f_1_sum = i2f_sum + i2f_1_io_covSum;
  assign io_covSum = i2f_1_sum;
  assign i2f_metaAssert_wire = i2f_metaAssert;
  assign i2f_1_metaAssert_wire = i2f_1_metaAssert;
  assign IntToFP_or0 = i2f_metaAssert_wire | i2f_1_metaAssert_wire;
  assign metaAssert = IntToFP_metaAssert;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  inPipe_valid = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  inPipe_bits_typeTagIn = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  inPipe_bits_wflags = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  inPipe_bits_rm = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  inPipe_bits_typ = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {2{`RANDOM}};
  inPipe_bits_in1 = _RAND_5[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {3{`RANDOM}};
  io_out_b_data = _RAND_6[64:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  io_out_b_exc = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  IntToFP_state = _RAND_8[3:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    IntToFP_cov[initvar] = _RAND_9[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  IntToFP_covSum = _RAND_10[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  IntToFP_metaAssert = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      inPipe_valid <= 1'h0;
    end else if (reset) begin
      inPipe_valid <= 1'h0;
    end else begin
      inPipe_valid <= io_in_valid;
    end
    if (metaReset) begin
      inPipe_bits_typeTagIn <= 2'h0;
    end else if (io_in_valid) begin
      inPipe_bits_typeTagIn <= io_in_bits_typeTagIn;
    end
    if (metaReset) begin
      inPipe_bits_wflags <= 1'h0;
    end else if (io_in_valid) begin
      inPipe_bits_wflags <= io_in_bits_wflags;
    end
    if (metaReset) begin
      inPipe_bits_rm <= 3'h0;
    end else if (io_in_valid) begin
      inPipe_bits_rm <= io_in_bits_rm;
    end
    if (metaReset) begin
      inPipe_bits_typ <= 2'h0;
    end else if (io_in_valid) begin
      inPipe_bits_typ <= io_in_bits_typ;
    end
    if (metaReset) begin
      inPipe_bits_in1 <= 64'h0;
    end else if (io_in_valid) begin
      inPipe_bits_in1 <= io_in_bits_in1;
    end
    if (metaReset) begin
      io_out_b_data <= 65'h0;
    end else if (inPipe_valid) begin
      if (inPipe_bits_wflags) begin
        if (mux_data_truncIdx) begin
          if (_T_1) begin
            io_out_b_data <= maskedNaN;
          end else begin
            io_out_b_data <= i2f_1_io_out;
          end
        end else begin
          io_out_b_data <= dataPadded_0;
        end
      end else if (_mux_data_T_12) begin
        io_out_b_data <= mux_data_swizzledNaN;
      end else begin
        io_out_b_data <= _mux_data_T_6;
      end
    end
    if (metaReset) begin
      io_out_b_exc <= 5'h0;
    end else if (inPipe_valid) begin
      if (inPipe_bits_wflags) begin
        if (mux_data_truncIdx) begin
          io_out_b_exc <= i2f_1_io_exceptionFlags;
        end else begin
          io_out_b_exc <= i2f_io_exceptionFlags;
        end
      end else begin
        io_out_b_exc <= 5'h0;
      end
    end
    IntToFP_state <= IntToFP_xor0;
    if (!(IntToFP_cov_read_data)) begin
      IntToFP_covSum <= IntToFP_covSum + 1'h1;
    end
    if (metaReset) begin
      IntToFP_metaAssert <= 1'h0;
    end else begin
      IntToFP_metaAssert <= IntToFP_metaAssert | IntToFP_or0;
    end
  end
  always @(posedge clock) begin
    if(IntToFP_cov_write_en & IntToFP_cov_write_mask) begin
      IntToFP_cov[IntToFP_cov_write_addr] <= IntToFP_cov_write_data; // @[Coverage map for IntToFP]
    end
  end
endmodule
module FPToFP(
  input         clock,
  input         reset,
  input         io_in_valid,
  input         io_in_bits_ren2,
  input  [1:0]  io_in_bits_typeTagOut,
  input         io_in_bits_wflags,
  input  [2:0]  io_in_bits_rm,
  input  [64:0] io_in_bits_in1,
  input  [64:0] io_in_bits_in2,
  output [64:0] io_out_bits_data,
  output [4:0]  io_out_bits_exc,
  input         io_lt,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  wire [64:0] narrower_io_in; // @[FPU.scala 614:30]
  wire [2:0] narrower_io_roundingMode; // @[FPU.scala 614:30]
  wire [32:0] narrower_io_out; // @[FPU.scala 614:30]
  wire [4:0] narrower_io_exceptionFlags; // @[FPU.scala 614:30]
  wire [29:0] narrower_io_covSum; // @[FPU.scala 614:30]
  wire  narrower_metaAssert; // @[FPU.scala 614:30]
  reg  inPipe_valid; // @[Valid.scala 117:22]
  reg [31:0] _RAND_0;
  reg  inPipe_bits_ren2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  reg [1:0] inPipe_bits_typeTagOut; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg  inPipe_bits_wflags; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg [2:0] inPipe_bits_rm; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg [64:0] inPipe_bits_in1; // @[Reg.scala 15:16]
  reg [95:0] _RAND_5;
  reg [64:0] inPipe_bits_in2; // @[Reg.scala 15:16]
  reg [95:0] _RAND_6;
  wire [64:0] _signNum_T_1; // @[FPU.scala 577:48]
  wire [64:0] _signNum_T_4; // @[FPU.scala 577:66]
  wire [64:0] signNum; // @[FPU.scala 577:20]
  wire  fsgnj_hi; // @[FPU.scala 578:26]
  wire [63:0] fsgnj_lo; // @[FPU.scala 578:45]
  wire [64:0] fsgnj; // @[Cat.scala 30:58]
  wire  isnan1; // @[FPU.scala 243:56]
  wire  isnan2; // @[FPU.scala 243:56]
  wire  _isInvalid_T_4; // @[FPU.scala 244:34]
  wire  _isInvalid_T_9; // @[FPU.scala 244:34]
  wire  isInvalid; // @[FPU.scala 587:49]
  wire  isNaNOut; // @[FPU.scala 588:27]
  wire  _isLHS_T_1; // @[FPU.scala 589:41]
  wire  _isLHS_T_3; // @[FPU.scala 589:51]
  wire  isLHS; // @[FPU.scala 589:24]
  wire [4:0] _fsgnjMux_exc_T; // @[FPU.scala 590:31]
  wire [64:0] _fsgnjMux_data_T; // @[FPU.scala 591:53]
  wire [64:0] _fsgnjMux_data_T_1; // @[FPU.scala 591:25]
  wire [64:0] _GEN_24; // @[FPU.scala 584:25]
  wire  _T; // @[FPU.scala 598:18]
  wire  _T_2; // @[FPU.scala 603:24]
  wire [64:0] widened; // @[FPU.scala 606:24]
  wire [64:0] fsgnjMux_data; // @[FPU.scala 603:42]
  wire [31:0] mux_data_hi; // @[FPU.scala 599:37]
  wire  mux_data_hi_hi; // @[FPU.scala 268:17]
  wire [51:0] mux_data_fractIn; // @[FPU.scala 269:20]
  wire [11:0] mux_data_expIn; // @[FPU.scala 270:18]
  wire [75:0] _mux_data_fractOut_T; // @[FPU.scala 271:28]
  wire [22:0] mux_data_lo; // @[FPU.scala 271:38]
  wire [2:0] mux_data_expOut_hi; // @[FPU.scala 273:26]
  wire [11:0] _mux_data_expOut_commonCase_T_1; // @[FPU.scala 274:31]
  wire [11:0] mux_data_expOut_commonCase; // @[FPU.scala 274:48]
  wire  _mux_data_expOut_T; // @[FPU.scala 275:19]
  wire  _mux_data_expOut_T_1; // @[FPU.scala 275:36]
  wire  _mux_data_expOut_T_2; // @[FPU.scala 275:25]
  wire [5:0] mux_data_expOut_lo; // @[FPU.scala 275:65]
  wire [8:0] _mux_data_expOut_T_3; // @[Cat.scala 30:58]
  wire [8:0] mux_data_hi_lo; // @[FPU.scala 275:10]
  wire [64:0] _mux_data_T; // @[Cat.scala 30:58]
  wire [4:0] _fsgnjMux_exc_T_6; // @[FPU.scala 608:51]
  wire [64:0] _mux_data_T_1; // @[Cat.scala 30:58]
  reg [64:0] io_out_b_data; // @[Reg.scala 15:16]
  reg [95:0] _RAND_7;
  reg [4:0] io_out_b_exc; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8;
  reg [5:0] FPToFP_state; // @[Register tracking FPToFP state]
  reg [31:0] _RAND_9;
  reg  FPToFP_cov [0:63]; // @[Coverage map for FPToFP]
  reg [31:0] _RAND_10;
  wire  FPToFP_cov_read_data; // @[Coverage map for FPToFP]
  wire [5:0] FPToFP_cov_read_addr; // @[Coverage map for FPToFP]
  wire  FPToFP_cov_write_data; // @[Coverage map for FPToFP]
  wire [5:0] FPToFP_cov_write_addr; // @[Coverage map for FPToFP]
  wire  FPToFP_cov_write_mask; // @[Coverage map for FPToFP]
  wire  FPToFP_cov_write_en; // @[Coverage map for FPToFP]
  reg [29:0] FPToFP_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_11;
  wire  inPipe_valid_shl;
  wire [5:0] inPipe_valid_pad;
  wire [1:0] inPipe_bits_ren2_shl;
  wire [5:0] inPipe_bits_ren2_pad;
  wire [2:0] inPipe_bits_wflags_shl;
  wire [5:0] inPipe_bits_wflags_pad;
  wire [5:0] inPipe_bits_rm_shl;
  wire [5:0] inPipe_bits_rm_pad;
  wire [5:0] FPToFP_xor1;
  wire [5:0] FPToFP_xor2;
  wire [5:0] FPToFP_xor0;
  wire [29:0] narrower_sum;
  wire  narrower_metaAssert_wire;
  reg  FPToFP_metaAssert;
  reg [31:0] _RAND_12;
  RecFNToRecFN narrower ( // @[FPU.scala 614:30]
    .io_in(narrower_io_in),
    .io_roundingMode(narrower_io_roundingMode),
    .io_out(narrower_io_out),
    .io_exceptionFlags(narrower_io_exceptionFlags),
    .io_covSum(narrower_io_covSum),
    .metaAssert(narrower_metaAssert)
  );
  assign _signNum_T_1 = inPipe_bits_in1 ^ inPipe_bits_in2; // @[FPU.scala 577:48]
  assign _signNum_T_4 = inPipe_bits_rm[0] ? ~inPipe_bits_in2 : inPipe_bits_in2; // @[FPU.scala 577:66]
  assign signNum = inPipe_bits_rm[1] ? _signNum_T_1 : _signNum_T_4; // @[FPU.scala 577:20]
  assign fsgnj_hi = signNum[64]; // @[FPU.scala 578:26]
  assign fsgnj_lo = inPipe_bits_in1[63:0]; // @[FPU.scala 578:45]
  assign fsgnj = {fsgnj_hi,fsgnj_lo}; // @[Cat.scala 30:58]
  assign isnan1 = &inPipe_bits_in1[63:61]; // @[FPU.scala 243:56]
  assign isnan2 = &inPipe_bits_in2[63:61]; // @[FPU.scala 243:56]
  assign _isInvalid_T_4 = isnan1 & ~inPipe_bits_in1[51]; // @[FPU.scala 244:34]
  assign _isInvalid_T_9 = isnan2 & ~inPipe_bits_in2[51]; // @[FPU.scala 244:34]
  assign isInvalid = _isInvalid_T_4 | _isInvalid_T_9; // @[FPU.scala 587:49]
  assign isNaNOut = isnan1 & isnan2; // @[FPU.scala 588:27]
  assign _isLHS_T_1 = inPipe_bits_rm[0] != io_lt; // @[FPU.scala 589:41]
  assign _isLHS_T_3 = _isLHS_T_1 & ~isnan1; // @[FPU.scala 589:51]
  assign isLHS = isnan2 | _isLHS_T_3; // @[FPU.scala 589:24]
  assign _fsgnjMux_exc_T = {isInvalid, 4'h0}; // @[FPU.scala 590:31]
  assign _fsgnjMux_data_T = isLHS ? inPipe_bits_in1 : inPipe_bits_in2; // @[FPU.scala 591:53]
  assign _fsgnjMux_data_T_1 = isNaNOut ? 65'he008000000000000 : _fsgnjMux_data_T; // @[FPU.scala 591:25]
  assign _GEN_24 = inPipe_bits_wflags ? _fsgnjMux_data_T_1 : fsgnj; // @[FPU.scala 584:25]
  assign _T = inPipe_bits_typeTagOut == 2'h0; // @[FPU.scala 598:18]
  assign _T_2 = inPipe_bits_wflags & ~inPipe_bits_ren2; // @[FPU.scala 603:24]
  assign widened = isnan1 ? 65'he008000000000000 : inPipe_bits_in1; // @[FPU.scala 606:24]
  assign fsgnjMux_data = _T_2 ? widened : _GEN_24; // @[FPU.scala 603:42]
  assign mux_data_hi = fsgnjMux_data[64:33]; // @[FPU.scala 599:37]
  assign mux_data_hi_hi = fsgnjMux_data[64]; // @[FPU.scala 268:17]
  assign mux_data_fractIn = fsgnjMux_data[51:0]; // @[FPU.scala 269:20]
  assign mux_data_expIn = fsgnjMux_data[63:52]; // @[FPU.scala 270:18]
  assign _mux_data_fractOut_T = {mux_data_fractIn, 24'h0}; // @[FPU.scala 271:28]
  assign mux_data_lo = _mux_data_fractOut_T[75:53]; // @[FPU.scala 271:38]
  assign mux_data_expOut_hi = mux_data_expIn[11:9]; // @[FPU.scala 273:26]
  assign _mux_data_expOut_commonCase_T_1 = mux_data_expIn + 12'h100; // @[FPU.scala 274:31]
  assign mux_data_expOut_commonCase = _mux_data_expOut_commonCase_T_1 - 12'h800; // @[FPU.scala 274:48]
  assign _mux_data_expOut_T = mux_data_expOut_hi == 3'h0; // @[FPU.scala 275:19]
  assign _mux_data_expOut_T_1 = mux_data_expOut_hi >= 3'h6; // @[FPU.scala 275:36]
  assign _mux_data_expOut_T_2 = _mux_data_expOut_T | _mux_data_expOut_T_1; // @[FPU.scala 275:25]
  assign mux_data_expOut_lo = mux_data_expOut_commonCase[5:0]; // @[FPU.scala 275:65]
  assign _mux_data_expOut_T_3 = {mux_data_expOut_hi,mux_data_expOut_lo}; // @[Cat.scala 30:58]
  assign mux_data_hi_lo = _mux_data_expOut_T_2 ? _mux_data_expOut_T_3 : mux_data_expOut_commonCase[8:0]; // @[FPU.scala 275:10]
  assign _mux_data_T = {mux_data_hi,mux_data_hi_hi,mux_data_hi_lo,mux_data_lo}; // @[Cat.scala 30:58]
  assign _fsgnjMux_exc_T_6 = {_isInvalid_T_4, 4'h0}; // @[FPU.scala 608:51]
  assign _mux_data_T_1 = {mux_data_hi,narrower_io_out}; // @[Cat.scala 30:58]
  assign io_out_bits_data = io_out_b_data; // @[FPU.scala 625:10]
  assign io_out_bits_exc = io_out_b_exc; // @[FPU.scala 625:10]
  assign narrower_io_in = inPipe_bits_in1; // @[FPU.scala 615:24]
  assign narrower_io_roundingMode = inPipe_bits_rm; // @[FPU.scala 616:34]
  assign FPToFP_cov_read_addr = FPToFP_state;
  assign FPToFP_cov_read_data = FPToFP_cov[FPToFP_cov_read_addr]; // @[Coverage map for FPToFP]
  assign FPToFP_cov_write_data = 1'h1;
  assign FPToFP_cov_write_addr = FPToFP_state;
  assign FPToFP_cov_write_mask = 1'h1;
  assign FPToFP_cov_write_en = 1'h1;
  assign inPipe_valid_shl = inPipe_valid;
  assign inPipe_valid_pad = {5'h0,inPipe_valid_shl};
  assign inPipe_bits_ren2_shl = {inPipe_bits_ren2, 1'h0};
  assign inPipe_bits_ren2_pad = {4'h0,inPipe_bits_ren2_shl};
  assign inPipe_bits_wflags_shl = {inPipe_bits_wflags, 2'h0};
  assign inPipe_bits_wflags_pad = {3'h0,inPipe_bits_wflags_shl};
  assign inPipe_bits_rm_shl = {inPipe_bits_rm, 3'h0};
  assign inPipe_bits_rm_pad = inPipe_bits_rm_shl;
  assign FPToFP_xor1 = inPipe_valid_pad ^ inPipe_bits_ren2_pad;
  assign FPToFP_xor2 = inPipe_bits_wflags_pad ^ inPipe_bits_rm_pad;
  assign FPToFP_xor0 = FPToFP_xor1 ^ FPToFP_xor2;
  assign narrower_sum = FPToFP_covSum + narrower_io_covSum;
  assign io_covSum = narrower_sum;
  assign narrower_metaAssert_wire = narrower_metaAssert;
  assign metaAssert = FPToFP_metaAssert;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  inPipe_valid = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  inPipe_bits_ren2 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  inPipe_bits_typeTagOut = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  inPipe_bits_wflags = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  inPipe_bits_rm = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {3{`RANDOM}};
  inPipe_bits_in1 = _RAND_5[64:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {3{`RANDOM}};
  inPipe_bits_in2 = _RAND_6[64:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {3{`RANDOM}};
  io_out_b_data = _RAND_7[64:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  io_out_b_exc = _RAND_8[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  FPToFP_state = _RAND_9[5:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    FPToFP_cov[initvar] = _RAND_10[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  FPToFP_covSum = _RAND_11[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  FPToFP_metaAssert = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      inPipe_valid <= 1'h0;
    end else if (reset) begin
      inPipe_valid <= 1'h0;
    end else begin
      inPipe_valid <= io_in_valid;
    end
    if (metaReset) begin
      inPipe_bits_ren2 <= 1'h0;
    end else if (io_in_valid) begin
      inPipe_bits_ren2 <= io_in_bits_ren2;
    end
    if (metaReset) begin
      inPipe_bits_typeTagOut <= 2'h0;
    end else if (io_in_valid) begin
      inPipe_bits_typeTagOut <= io_in_bits_typeTagOut;
    end
    if (metaReset) begin
      inPipe_bits_wflags <= 1'h0;
    end else if (io_in_valid) begin
      inPipe_bits_wflags <= io_in_bits_wflags;
    end
    if (metaReset) begin
      inPipe_bits_rm <= 3'h0;
    end else if (io_in_valid) begin
      inPipe_bits_rm <= io_in_bits_rm;
    end
    if (metaReset) begin
      inPipe_bits_in1 <= 65'h0;
    end else if (io_in_valid) begin
      inPipe_bits_in1 <= io_in_bits_in1;
    end
    if (metaReset) begin
      inPipe_bits_in2 <= 65'h0;
    end else if (io_in_valid) begin
      inPipe_bits_in2 <= io_in_bits_in2;
    end
    if (metaReset) begin
      io_out_b_data <= 65'h0;
    end else if (inPipe_valid) begin
      if (_T_2) begin
        if (_T) begin
          io_out_b_data <= _mux_data_T_1;
        end else if (_T) begin
          io_out_b_data <= _mux_data_T;
        end else if (_T_2) begin
          if (isnan1) begin
            io_out_b_data <= 65'he008000000000000;
          end else begin
            io_out_b_data <= inPipe_bits_in1;
          end
        end else if (inPipe_bits_wflags) begin
          if (isNaNOut) begin
            io_out_b_data <= 65'he008000000000000;
          end else if (isLHS) begin
            io_out_b_data <= inPipe_bits_in1;
          end else begin
            io_out_b_data <= inPipe_bits_in2;
          end
        end else begin
          io_out_b_data <= fsgnj;
        end
      end else if (_T) begin
        io_out_b_data <= _mux_data_T;
      end else if (_T_2) begin
        if (isnan1) begin
          io_out_b_data <= 65'he008000000000000;
        end else begin
          io_out_b_data <= inPipe_bits_in1;
        end
      end else if (inPipe_bits_wflags) begin
        if (isNaNOut) begin
          io_out_b_data <= 65'he008000000000000;
        end else if (isLHS) begin
          io_out_b_data <= inPipe_bits_in1;
        end else begin
          io_out_b_data <= inPipe_bits_in2;
        end
      end else begin
        io_out_b_data <= fsgnj;
      end
    end
    if (metaReset) begin
      io_out_b_exc <= 5'h0;
    end else if (inPipe_valid) begin
      if (_T_2) begin
        if (_T) begin
          io_out_b_exc <= narrower_io_exceptionFlags;
        end else if (_T_2) begin
          io_out_b_exc <= _fsgnjMux_exc_T_6;
        end else if (inPipe_bits_wflags) begin
          io_out_b_exc <= _fsgnjMux_exc_T;
        end else begin
          io_out_b_exc <= 5'h0;
        end
      end else if (_T_2) begin
        io_out_b_exc <= _fsgnjMux_exc_T_6;
      end else if (inPipe_bits_wflags) begin
        io_out_b_exc <= _fsgnjMux_exc_T;
      end else begin
        io_out_b_exc <= 5'h0;
      end
    end
    FPToFP_state <= FPToFP_xor0;
    if (!(FPToFP_cov_read_data)) begin
      FPToFP_covSum <= FPToFP_covSum + 1'h1;
    end
    if (metaReset) begin
      FPToFP_metaAssert <= 1'h0;
    end else begin
      FPToFP_metaAssert <= FPToFP_metaAssert | narrower_metaAssert_wire;
    end
  end
  always @(posedge clock) begin
    if(FPToFP_cov_write_en & FPToFP_cov_write_mask) begin
      FPToFP_cov[FPToFP_cov_write_addr] <= FPToFP_cov_write_data; // @[Coverage map for FPToFP]
    end
  end
endmodule
module FPUFMAPipe_1(
  input         clock,
  input         reset,
  input         io_in_valid,
  input         io_in_bits_ren3,
  input         io_in_bits_swap23,
  input  [2:0]  io_in_bits_rm,
  input  [1:0]  io_in_bits_fmaCmd,
  input  [64:0] io_in_bits_in1,
  input  [64:0] io_in_bits_in2,
  input  [64:0] io_in_bits_in3,
  output [64:0] io_out_bits_data,
  output [4:0]  io_out_bits_exc,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset,
  input         fma_halt
);
  wire  fma_clock; // @[FPU.scala 712:19]
  wire  fma_reset; // @[FPU.scala 712:19]
  wire  fma_io_validin; // @[FPU.scala 712:19]
  wire [1:0] fma_io_op; // @[FPU.scala 712:19]
  wire [64:0] fma_io_a; // @[FPU.scala 712:19]
  wire [64:0] fma_io_b; // @[FPU.scala 712:19]
  wire [64:0] fma_io_c; // @[FPU.scala 712:19]
  wire [2:0] fma_io_roundingMode; // @[FPU.scala 712:19]
  wire [64:0] fma_io_out; // @[FPU.scala 712:19]
  wire [4:0] fma_io_exceptionFlags; // @[FPU.scala 712:19]
  wire  fma_io_validout; // @[FPU.scala 712:19]
  wire [29:0] fma_io_covSum; // @[FPU.scala 712:19]
  wire  fma_metaAssert; // @[FPU.scala 712:19]
  wire  fma_metaReset; // @[FPU.scala 712:19]
  reg  valid; // @[FPU.scala 700:18]
  reg [31:0] _RAND_0;
  reg [2:0] in_rm; // @[FPU.scala 701:15]
  reg [31:0] _RAND_1;
  reg [1:0] in_fmaCmd; // @[FPU.scala 701:15]
  reg [31:0] _RAND_2;
  reg [64:0] in_in1; // @[FPU.scala 701:15]
  reg [95:0] _RAND_3;
  reg [64:0] in_in2; // @[FPU.scala 701:15]
  reg [95:0] _RAND_4;
  reg [64:0] in_in3; // @[FPU.scala 701:15]
  reg [95:0] _RAND_5;
  wire [64:0] _zero_T; // @[FPU.scala 704:32]
  wire [64:0] zero; // @[FPU.scala 704:50]
  wire  _T; // @[FPU.scala 709:21]
  wire [64:0] res_data_maskedNaN; // @[FPU.scala 408:25]
  wire  _res_data_T_1; // @[FPU.scala 243:56]
  reg [64:0] io_out_b_data; // @[Reg.scala 15:16]
  reg [95:0] _RAND_6;
  reg [4:0] io_out_b_exc; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7;
  wire [4:0] res_exc; // @[FPU.scala 721:17 FPU.scala 723:11]
  wire [29:0] FPUFMAPipe_1_covSum;
  wire [29:0] fma_sum;
  wire  fma_metaAssert_wire;
  reg  FPUFMAPipe_1_metaAssert;
  reg [31:0] _RAND_8;
  MulAddRecFNPipe_1 fma ( // @[FPU.scala 712:19]
    .clock(fma_clock),
    .reset(fma_reset),
    .io_validin(fma_io_validin),
    .io_op(fma_io_op),
    .io_a(fma_io_a),
    .io_b(fma_io_b),
    .io_c(fma_io_c),
    .io_roundingMode(fma_io_roundingMode),
    .io_out(fma_io_out),
    .io_exceptionFlags(fma_io_exceptionFlags),
    .io_validout(fma_io_validout),
    .io_covSum(fma_io_covSum),
    .metaAssert(fma_metaAssert),
    .metaReset(fma_metaReset)
  );
  assign _zero_T = io_in_bits_in1 ^ io_in_bits_in2; // @[FPU.scala 704:32]
  assign zero = _zero_T & 65'h10000000000000000; // @[FPU.scala 704:50]
  assign _T = io_in_bits_ren3 | io_in_bits_swap23; // @[FPU.scala 709:21]
  assign res_data_maskedNaN = fma_io_out & 65'h1efefffffffffffff; // @[FPU.scala 408:25]
  assign _res_data_T_1 = &fma_io_out[63:61]; // @[FPU.scala 243:56]
  assign res_exc = fma_io_exceptionFlags; // @[FPU.scala 721:17 FPU.scala 723:11]
  assign io_out_bits_data = io_out_b_data; // @[FPU.scala 725:10]
  assign io_out_bits_exc = io_out_b_exc; // @[FPU.scala 725:10]
  assign fma_clock = clock;
  assign fma_reset = reset;
  assign fma_io_validin = valid; // @[FPU.scala 713:18]
  assign fma_io_op = in_fmaCmd; // @[FPU.scala 714:13]
  assign fma_io_a = in_in1; // @[FPU.scala 717:12]
  assign fma_io_b = in_in2; // @[FPU.scala 718:12]
  assign fma_io_c = in_in3; // @[FPU.scala 719:12]
  assign fma_io_roundingMode = in_rm; // @[FPU.scala 715:23]
  assign FPUFMAPipe_1_covSum = 30'h0;
  assign fma_sum = FPUFMAPipe_1_covSum + fma_io_covSum;
  assign io_covSum = fma_sum;
  assign fma_metaAssert_wire = fma_metaAssert;
  assign metaAssert = FPUFMAPipe_1_metaAssert;
  assign fma_metaReset = metaReset | fma_halt;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  valid = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  in_rm = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  in_fmaCmd = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {3{`RANDOM}};
  in_in1 = _RAND_3[64:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {3{`RANDOM}};
  in_in2 = _RAND_4[64:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {3{`RANDOM}};
  in_in3 = _RAND_5[64:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {3{`RANDOM}};
  io_out_b_data = _RAND_6[64:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  io_out_b_exc = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  FPUFMAPipe_1_metaAssert = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      valid <= 1'h0;
    end else begin
      valid <= io_in_valid;
    end
    if (metaReset) begin
      in_rm <= 3'h0;
    end else if (io_in_valid) begin
      in_rm <= io_in_bits_rm;
    end
    if (metaReset) begin
      in_fmaCmd <= 2'h0;
    end else if (io_in_valid) begin
      in_fmaCmd <= io_in_bits_fmaCmd;
    end
    if (metaReset) begin
      in_in1 <= 65'h0;
    end else if (io_in_valid) begin
      in_in1 <= io_in_bits_in1;
    end
    if (metaReset) begin
      in_in2 <= 65'h0;
    end else if (io_in_valid) begin
      if (io_in_bits_swap23) begin
        in_in2 <= 65'h8000000000000000;
      end else begin
        in_in2 <= io_in_bits_in2;
      end
    end
    if (metaReset) begin
      in_in3 <= 65'h0;
    end else if (io_in_valid) begin
      if (~_T) begin
        in_in3 <= zero;
      end else begin
        in_in3 <= io_in_bits_in3;
      end
    end
    if (metaReset) begin
      io_out_b_data <= 65'h0;
    end else if (fma_io_validout) begin
      if (_res_data_T_1) begin
        io_out_b_data <= res_data_maskedNaN;
      end else begin
        io_out_b_data <= fma_io_out;
      end
    end
    if (metaReset) begin
      io_out_b_exc <= 5'h0;
    end else if (fma_io_validout) begin
      io_out_b_exc <= res_exc;
    end
    if (metaReset) begin
      FPUFMAPipe_1_metaAssert <= 1'h0;
    end else begin
      FPUFMAPipe_1_metaAssert <= FPUFMAPipe_1_metaAssert | fma_metaAssert_wire;
    end
  end
endmodule
module DivSqrtRecFN_small(
  input         clock,
  input         reset,
  output        io_inReady,
  input         io_inValid,
  input         io_sqrtOp,
  input  [32:0] io_a,
  input  [32:0] io_b,
  input  [2:0]  io_roundingMode,
  output        io_outValid_div,
  output        io_outValid_sqrt,
  output [32:0] io_out,
  output [4:0]  io_exceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset,
  input         divSqrtRecFNToRaw_halt
);
  wire  divSqrtRecFNToRaw_clock; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_reset; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_io_inReady; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_io_inValid; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_io_sqrtOp; // @[DivSqrtRecFN_small.scala 462:15]
  wire [32:0] divSqrtRecFNToRaw_io_a; // @[DivSqrtRecFN_small.scala 462:15]
  wire [32:0] divSqrtRecFNToRaw_io_b; // @[DivSqrtRecFN_small.scala 462:15]
  wire [2:0] divSqrtRecFNToRaw_io_roundingMode; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_io_rawOutValid_div; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_io_rawOutValid_sqrt; // @[DivSqrtRecFN_small.scala 462:15]
  wire [2:0] divSqrtRecFNToRaw_io_roundingModeOut; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_io_invalidExc; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_io_infiniteExc; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_io_rawOut_isNaN; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_io_rawOut_isInf; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_io_rawOut_isZero; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_io_rawOut_sign; // @[DivSqrtRecFN_small.scala 462:15]
  wire [9:0] divSqrtRecFNToRaw_io_rawOut_sExp; // @[DivSqrtRecFN_small.scala 462:15]
  wire [26:0] divSqrtRecFNToRaw_io_rawOut_sig; // @[DivSqrtRecFN_small.scala 462:15]
  wire [29:0] divSqrtRecFNToRaw_io_covSum; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_metaAssert; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_metaReset; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_divSqrtRawFN__halt; // @[DivSqrtRecFN_small.scala 462:15]
  wire  roundRawFNToRecFN_io_invalidExc; // @[DivSqrtRecFN_small.scala 477:15]
  wire  roundRawFNToRecFN_io_infiniteExc; // @[DivSqrtRecFN_small.scala 477:15]
  wire  roundRawFNToRecFN_io_in_isNaN; // @[DivSqrtRecFN_small.scala 477:15]
  wire  roundRawFNToRecFN_io_in_isInf; // @[DivSqrtRecFN_small.scala 477:15]
  wire  roundRawFNToRecFN_io_in_isZero; // @[DivSqrtRecFN_small.scala 477:15]
  wire  roundRawFNToRecFN_io_in_sign; // @[DivSqrtRecFN_small.scala 477:15]
  wire [9:0] roundRawFNToRecFN_io_in_sExp; // @[DivSqrtRecFN_small.scala 477:15]
  wire [26:0] roundRawFNToRecFN_io_in_sig; // @[DivSqrtRecFN_small.scala 477:15]
  wire [2:0] roundRawFNToRecFN_io_roundingMode; // @[DivSqrtRecFN_small.scala 477:15]
  wire  roundRawFNToRecFN_io_detectTininess; // @[DivSqrtRecFN_small.scala 477:15]
  wire [32:0] roundRawFNToRecFN_io_out; // @[DivSqrtRecFN_small.scala 477:15]
  wire [4:0] roundRawFNToRecFN_io_exceptionFlags; // @[DivSqrtRecFN_small.scala 477:15]
  wire [29:0] roundRawFNToRecFN_io_covSum; // @[DivSqrtRecFN_small.scala 477:15]
  wire  roundRawFNToRecFN_metaAssert; // @[DivSqrtRecFN_small.scala 477:15]
  wire [29:0] DivSqrtRecFN_small_covSum;
  wire [29:0] divSqrtRecFNToRaw_sum;
  wire [29:0] roundRawFNToRecFN_sum;
  wire  divSqrtRecFNToRaw_metaAssert_wire;
  wire  roundRawFNToRecFN_metaAssert_wire;
  wire  DivSqrtRecFN_small_or0;
  reg  DivSqrtRecFN_small_metaAssert;
  reg [31:0] _RAND_0;
  DivSqrtRecFNToRaw_small divSqrtRecFNToRaw ( // @[DivSqrtRecFN_small.scala 462:15]
    .clock(divSqrtRecFNToRaw_clock),
    .reset(divSqrtRecFNToRaw_reset),
    .io_inReady(divSqrtRecFNToRaw_io_inReady),
    .io_inValid(divSqrtRecFNToRaw_io_inValid),
    .io_sqrtOp(divSqrtRecFNToRaw_io_sqrtOp),
    .io_a(divSqrtRecFNToRaw_io_a),
    .io_b(divSqrtRecFNToRaw_io_b),
    .io_roundingMode(divSqrtRecFNToRaw_io_roundingMode),
    .io_rawOutValid_div(divSqrtRecFNToRaw_io_rawOutValid_div),
    .io_rawOutValid_sqrt(divSqrtRecFNToRaw_io_rawOutValid_sqrt),
    .io_roundingModeOut(divSqrtRecFNToRaw_io_roundingModeOut),
    .io_invalidExc(divSqrtRecFNToRaw_io_invalidExc),
    .io_infiniteExc(divSqrtRecFNToRaw_io_infiniteExc),
    .io_rawOut_isNaN(divSqrtRecFNToRaw_io_rawOut_isNaN),
    .io_rawOut_isInf(divSqrtRecFNToRaw_io_rawOut_isInf),
    .io_rawOut_isZero(divSqrtRecFNToRaw_io_rawOut_isZero),
    .io_rawOut_sign(divSqrtRecFNToRaw_io_rawOut_sign),
    .io_rawOut_sExp(divSqrtRecFNToRaw_io_rawOut_sExp),
    .io_rawOut_sig(divSqrtRecFNToRaw_io_rawOut_sig),
    .io_covSum(divSqrtRecFNToRaw_io_covSum),
    .metaAssert(divSqrtRecFNToRaw_metaAssert),
    .metaReset(divSqrtRecFNToRaw_metaReset),
    .divSqrtRawFN__halt(divSqrtRecFNToRaw_divSqrtRawFN__halt)
  );
  RoundRawFNToRecFN_2 roundRawFNToRecFN ( // @[DivSqrtRecFN_small.scala 477:15]
    .io_invalidExc(roundRawFNToRecFN_io_invalidExc),
    .io_infiniteExc(roundRawFNToRecFN_io_infiniteExc),
    .io_in_isNaN(roundRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundRawFNToRecFN_io_in_sig),
    .io_roundingMode(roundRawFNToRecFN_io_roundingMode),
    .io_detectTininess(roundRawFNToRecFN_io_detectTininess),
    .io_out(roundRawFNToRecFN_io_out),
    .io_exceptionFlags(roundRawFNToRecFN_io_exceptionFlags),
    .io_covSum(roundRawFNToRecFN_io_covSum),
    .metaAssert(roundRawFNToRecFN_metaAssert)
  );
  assign io_inReady = divSqrtRecFNToRaw_io_inReady; // @[DivSqrtRecFN_small.scala 464:16]
  assign io_outValid_div = divSqrtRecFNToRaw_io_rawOutValid_div; // @[DivSqrtRecFN_small.scala 473:22]
  assign io_outValid_sqrt = divSqrtRecFNToRaw_io_rawOutValid_sqrt; // @[DivSqrtRecFN_small.scala 474:22]
  assign io_out = roundRawFNToRecFN_io_out; // @[DivSqrtRecFN_small.scala 483:23]
  assign io_exceptionFlags = roundRawFNToRecFN_io_exceptionFlags; // @[DivSqrtRecFN_small.scala 484:23]
  assign divSqrtRecFNToRaw_clock = clock;
  assign divSqrtRecFNToRaw_reset = reset;
  assign divSqrtRecFNToRaw_io_inValid = io_inValid; // @[DivSqrtRecFN_small.scala 465:39]
  assign divSqrtRecFNToRaw_io_sqrtOp = io_sqrtOp; // @[DivSqrtRecFN_small.scala 466:39]
  assign divSqrtRecFNToRaw_io_a = io_a; // @[DivSqrtRecFN_small.scala 467:39]
  assign divSqrtRecFNToRaw_io_b = io_b; // @[DivSqrtRecFN_small.scala 468:39]
  assign divSqrtRecFNToRaw_io_roundingMode = io_roundingMode; // @[DivSqrtRecFN_small.scala 469:39]
  assign roundRawFNToRecFN_io_invalidExc = divSqrtRecFNToRaw_io_invalidExc; // @[DivSqrtRecFN_small.scala 478:39]
  assign roundRawFNToRecFN_io_infiniteExc = divSqrtRecFNToRaw_io_infiniteExc; // @[DivSqrtRecFN_small.scala 479:39]
  assign roundRawFNToRecFN_io_in_isNaN = divSqrtRecFNToRaw_io_rawOut_isNaN; // @[DivSqrtRecFN_small.scala 480:39]
  assign roundRawFNToRecFN_io_in_isInf = divSqrtRecFNToRaw_io_rawOut_isInf; // @[DivSqrtRecFN_small.scala 480:39]
  assign roundRawFNToRecFN_io_in_isZero = divSqrtRecFNToRaw_io_rawOut_isZero; // @[DivSqrtRecFN_small.scala 480:39]
  assign roundRawFNToRecFN_io_in_sign = divSqrtRecFNToRaw_io_rawOut_sign; // @[DivSqrtRecFN_small.scala 480:39]
  assign roundRawFNToRecFN_io_in_sExp = divSqrtRecFNToRaw_io_rawOut_sExp; // @[DivSqrtRecFN_small.scala 480:39]
  assign roundRawFNToRecFN_io_in_sig = divSqrtRecFNToRaw_io_rawOut_sig; // @[DivSqrtRecFN_small.scala 480:39]
  assign roundRawFNToRecFN_io_roundingMode = divSqrtRecFNToRaw_io_roundingModeOut; // @[DivSqrtRecFN_small.scala 481:39]
  assign roundRawFNToRecFN_io_detectTininess = 1'h1; // @[DivSqrtRecFN_small.scala 482:41]
  assign DivSqrtRecFN_small_covSum = 30'h0;
  assign divSqrtRecFNToRaw_sum = DivSqrtRecFN_small_covSum + divSqrtRecFNToRaw_io_covSum;
  assign roundRawFNToRecFN_sum = divSqrtRecFNToRaw_sum + roundRawFNToRecFN_io_covSum;
  assign io_covSum = roundRawFNToRecFN_sum;
  assign divSqrtRecFNToRaw_metaAssert_wire = divSqrtRecFNToRaw_metaAssert;
  assign roundRawFNToRecFN_metaAssert_wire = roundRawFNToRecFN_metaAssert;
  assign DivSqrtRecFN_small_or0 = divSqrtRecFNToRaw_metaAssert_wire | roundRawFNToRecFN_metaAssert_wire;
  assign metaAssert = DivSqrtRecFN_small_metaAssert;
  assign divSqrtRecFNToRaw_metaReset = metaReset | divSqrtRecFNToRaw_halt;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  DivSqrtRecFN_small_metaAssert = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      DivSqrtRecFN_small_metaAssert <= 1'h0;
    end else begin
      DivSqrtRecFN_small_metaAssert <= DivSqrtRecFN_small_metaAssert | DivSqrtRecFN_small_or0;
    end
  end
endmodule
module DivSqrtRecFN_small_1(
  input         clock,
  input         reset,
  output        io_inReady,
  input         io_inValid,
  input         io_sqrtOp,
  input  [64:0] io_a,
  input  [64:0] io_b,
  input  [2:0]  io_roundingMode,
  output        io_outValid_div,
  output        io_outValid_sqrt,
  output [64:0] io_out,
  output [4:0]  io_exceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset,
  input         divSqrtRecFNToRaw_halt
);
  wire  divSqrtRecFNToRaw_clock; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_reset; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_io_inReady; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_io_inValid; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_io_sqrtOp; // @[DivSqrtRecFN_small.scala 462:15]
  wire [64:0] divSqrtRecFNToRaw_io_a; // @[DivSqrtRecFN_small.scala 462:15]
  wire [64:0] divSqrtRecFNToRaw_io_b; // @[DivSqrtRecFN_small.scala 462:15]
  wire [2:0] divSqrtRecFNToRaw_io_roundingMode; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_io_rawOutValid_div; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_io_rawOutValid_sqrt; // @[DivSqrtRecFN_small.scala 462:15]
  wire [2:0] divSqrtRecFNToRaw_io_roundingModeOut; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_io_invalidExc; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_io_infiniteExc; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_io_rawOut_isNaN; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_io_rawOut_isInf; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_io_rawOut_isZero; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_io_rawOut_sign; // @[DivSqrtRecFN_small.scala 462:15]
  wire [12:0] divSqrtRecFNToRaw_io_rawOut_sExp; // @[DivSqrtRecFN_small.scala 462:15]
  wire [55:0] divSqrtRecFNToRaw_io_rawOut_sig; // @[DivSqrtRecFN_small.scala 462:15]
  wire [29:0] divSqrtRecFNToRaw_io_covSum; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_metaAssert; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_metaReset; // @[DivSqrtRecFN_small.scala 462:15]
  wire  divSqrtRecFNToRaw_divSqrtRawFN__halt; // @[DivSqrtRecFN_small.scala 462:15]
  wire  roundRawFNToRecFN_io_invalidExc; // @[DivSqrtRecFN_small.scala 477:15]
  wire  roundRawFNToRecFN_io_infiniteExc; // @[DivSqrtRecFN_small.scala 477:15]
  wire  roundRawFNToRecFN_io_in_isNaN; // @[DivSqrtRecFN_small.scala 477:15]
  wire  roundRawFNToRecFN_io_in_isInf; // @[DivSqrtRecFN_small.scala 477:15]
  wire  roundRawFNToRecFN_io_in_isZero; // @[DivSqrtRecFN_small.scala 477:15]
  wire  roundRawFNToRecFN_io_in_sign; // @[DivSqrtRecFN_small.scala 477:15]
  wire [12:0] roundRawFNToRecFN_io_in_sExp; // @[DivSqrtRecFN_small.scala 477:15]
  wire [55:0] roundRawFNToRecFN_io_in_sig; // @[DivSqrtRecFN_small.scala 477:15]
  wire [2:0] roundRawFNToRecFN_io_roundingMode; // @[DivSqrtRecFN_small.scala 477:15]
  wire  roundRawFNToRecFN_io_detectTininess; // @[DivSqrtRecFN_small.scala 477:15]
  wire [64:0] roundRawFNToRecFN_io_out; // @[DivSqrtRecFN_small.scala 477:15]
  wire [4:0] roundRawFNToRecFN_io_exceptionFlags; // @[DivSqrtRecFN_small.scala 477:15]
  wire [29:0] roundRawFNToRecFN_io_covSum; // @[DivSqrtRecFN_small.scala 477:15]
  wire  roundRawFNToRecFN_metaAssert; // @[DivSqrtRecFN_small.scala 477:15]
  wire [29:0] DivSqrtRecFN_small_1_covSum;
  wire [29:0] divSqrtRecFNToRaw_sum;
  wire [29:0] roundRawFNToRecFN_sum;
  wire  divSqrtRecFNToRaw_metaAssert_wire;
  wire  roundRawFNToRecFN_metaAssert_wire;
  wire  DivSqrtRecFN_small_1_or0;
  reg  DivSqrtRecFN_small_1_metaAssert;
  reg [31:0] _RAND_0;
  DivSqrtRecFNToRaw_small_1 divSqrtRecFNToRaw ( // @[DivSqrtRecFN_small.scala 462:15]
    .clock(divSqrtRecFNToRaw_clock),
    .reset(divSqrtRecFNToRaw_reset),
    .io_inReady(divSqrtRecFNToRaw_io_inReady),
    .io_inValid(divSqrtRecFNToRaw_io_inValid),
    .io_sqrtOp(divSqrtRecFNToRaw_io_sqrtOp),
    .io_a(divSqrtRecFNToRaw_io_a),
    .io_b(divSqrtRecFNToRaw_io_b),
    .io_roundingMode(divSqrtRecFNToRaw_io_roundingMode),
    .io_rawOutValid_div(divSqrtRecFNToRaw_io_rawOutValid_div),
    .io_rawOutValid_sqrt(divSqrtRecFNToRaw_io_rawOutValid_sqrt),
    .io_roundingModeOut(divSqrtRecFNToRaw_io_roundingModeOut),
    .io_invalidExc(divSqrtRecFNToRaw_io_invalidExc),
    .io_infiniteExc(divSqrtRecFNToRaw_io_infiniteExc),
    .io_rawOut_isNaN(divSqrtRecFNToRaw_io_rawOut_isNaN),
    .io_rawOut_isInf(divSqrtRecFNToRaw_io_rawOut_isInf),
    .io_rawOut_isZero(divSqrtRecFNToRaw_io_rawOut_isZero),
    .io_rawOut_sign(divSqrtRecFNToRaw_io_rawOut_sign),
    .io_rawOut_sExp(divSqrtRecFNToRaw_io_rawOut_sExp),
    .io_rawOut_sig(divSqrtRecFNToRaw_io_rawOut_sig),
    .io_covSum(divSqrtRecFNToRaw_io_covSum),
    .metaAssert(divSqrtRecFNToRaw_metaAssert),
    .metaReset(divSqrtRecFNToRaw_metaReset),
    .divSqrtRawFN__halt(divSqrtRecFNToRaw_divSqrtRawFN__halt)
  );
  RoundRawFNToRecFN_3 roundRawFNToRecFN ( // @[DivSqrtRecFN_small.scala 477:15]
    .io_invalidExc(roundRawFNToRecFN_io_invalidExc),
    .io_infiniteExc(roundRawFNToRecFN_io_infiniteExc),
    .io_in_isNaN(roundRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundRawFNToRecFN_io_in_sig),
    .io_roundingMode(roundRawFNToRecFN_io_roundingMode),
    .io_detectTininess(roundRawFNToRecFN_io_detectTininess),
    .io_out(roundRawFNToRecFN_io_out),
    .io_exceptionFlags(roundRawFNToRecFN_io_exceptionFlags),
    .io_covSum(roundRawFNToRecFN_io_covSum),
    .metaAssert(roundRawFNToRecFN_metaAssert)
  );
  assign io_inReady = divSqrtRecFNToRaw_io_inReady; // @[DivSqrtRecFN_small.scala 464:16]
  assign io_outValid_div = divSqrtRecFNToRaw_io_rawOutValid_div; // @[DivSqrtRecFN_small.scala 473:22]
  assign io_outValid_sqrt = divSqrtRecFNToRaw_io_rawOutValid_sqrt; // @[DivSqrtRecFN_small.scala 474:22]
  assign io_out = roundRawFNToRecFN_io_out; // @[DivSqrtRecFN_small.scala 483:23]
  assign io_exceptionFlags = roundRawFNToRecFN_io_exceptionFlags; // @[DivSqrtRecFN_small.scala 484:23]
  assign divSqrtRecFNToRaw_clock = clock;
  assign divSqrtRecFNToRaw_reset = reset;
  assign divSqrtRecFNToRaw_io_inValid = io_inValid; // @[DivSqrtRecFN_small.scala 465:39]
  assign divSqrtRecFNToRaw_io_sqrtOp = io_sqrtOp; // @[DivSqrtRecFN_small.scala 466:39]
  assign divSqrtRecFNToRaw_io_a = io_a; // @[DivSqrtRecFN_small.scala 467:39]
  assign divSqrtRecFNToRaw_io_b = io_b; // @[DivSqrtRecFN_small.scala 468:39]
  assign divSqrtRecFNToRaw_io_roundingMode = io_roundingMode; // @[DivSqrtRecFN_small.scala 469:39]
  assign roundRawFNToRecFN_io_invalidExc = divSqrtRecFNToRaw_io_invalidExc; // @[DivSqrtRecFN_small.scala 478:39]
  assign roundRawFNToRecFN_io_infiniteExc = divSqrtRecFNToRaw_io_infiniteExc; // @[DivSqrtRecFN_small.scala 479:39]
  assign roundRawFNToRecFN_io_in_isNaN = divSqrtRecFNToRaw_io_rawOut_isNaN; // @[DivSqrtRecFN_small.scala 480:39]
  assign roundRawFNToRecFN_io_in_isInf = divSqrtRecFNToRaw_io_rawOut_isInf; // @[DivSqrtRecFN_small.scala 480:39]
  assign roundRawFNToRecFN_io_in_isZero = divSqrtRecFNToRaw_io_rawOut_isZero; // @[DivSqrtRecFN_small.scala 480:39]
  assign roundRawFNToRecFN_io_in_sign = divSqrtRecFNToRaw_io_rawOut_sign; // @[DivSqrtRecFN_small.scala 480:39]
  assign roundRawFNToRecFN_io_in_sExp = divSqrtRecFNToRaw_io_rawOut_sExp; // @[DivSqrtRecFN_small.scala 480:39]
  assign roundRawFNToRecFN_io_in_sig = divSqrtRecFNToRaw_io_rawOut_sig; // @[DivSqrtRecFN_small.scala 480:39]
  assign roundRawFNToRecFN_io_roundingMode = divSqrtRecFNToRaw_io_roundingModeOut; // @[DivSqrtRecFN_small.scala 481:39]
  assign roundRawFNToRecFN_io_detectTininess = 1'h1; // @[DivSqrtRecFN_small.scala 482:41]
  assign DivSqrtRecFN_small_1_covSum = 30'h0;
  assign divSqrtRecFNToRaw_sum = DivSqrtRecFN_small_1_covSum + divSqrtRecFNToRaw_io_covSum;
  assign roundRawFNToRecFN_sum = divSqrtRecFNToRaw_sum + roundRawFNToRecFN_io_covSum;
  assign io_covSum = roundRawFNToRecFN_sum;
  assign divSqrtRecFNToRaw_metaAssert_wire = divSqrtRecFNToRaw_metaAssert;
  assign roundRawFNToRecFN_metaAssert_wire = roundRawFNToRecFN_metaAssert;
  assign DivSqrtRecFN_small_1_or0 = divSqrtRecFNToRaw_metaAssert_wire | roundRawFNToRecFN_metaAssert_wire;
  assign metaAssert = DivSqrtRecFN_small_1_metaAssert;
  assign divSqrtRecFNToRaw_metaReset = metaReset | divSqrtRecFNToRaw_halt;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  DivSqrtRecFN_small_1_metaAssert = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      DivSqrtRecFN_small_1_metaAssert <= 1'h0;
    end else begin
      DivSqrtRecFN_small_1_metaAssert <= DivSqrtRecFN_small_1_metaAssert | DivSqrtRecFN_small_1_or0;
    end
  end
endmodule
module Arbiter(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [26:0] io_in_0_bits_bits_addr,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input         io_in_1_bits_valid,
  input  [26:0] io_in_1_bits_bits_addr,
  input         io_out_ready,
  output        io_out_valid,
  output        io_out_bits_valid,
  output [26:0] io_out_bits_bits_addr,
  output        io_chosen,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  grant_1; // @[Arbiter.scala 31:78]
  wire [29:0] Arbiter_covSum;
  assign grant_1 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:14]
  assign io_in_1_ready = grant_1 & io_out_ready; // @[Arbiter.scala 134:14]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[Arbiter.scala 135:16]
  assign io_out_bits_valid = io_in_0_valid | io_in_1_bits_valid; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_out_bits_bits_addr = io_in_0_valid ? io_in_0_bits_bits_addr : io_in_1_bits_bits_addr; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_chosen = io_in_0_valid ? 1'h0 : 1'h1; // @[Arbiter.scala 123:13 Arbiter.scala 127:17]
  assign Arbiter_covSum = 30'h0;
  assign io_covSum = Arbiter_covSum;
  assign metaAssert = 1'h0;
endmodule
module OptimizationBarrier_42(
  input  [2:0]  io_x,
  output [2:0]  io_y,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire [29:0] OptimizationBarrier_42_covSum;
  assign io_y = io_x; // @[package.scala 263:12]
  assign OptimizationBarrier_42_covSum = 30'h0;
  assign io_covSum = OptimizationBarrier_42_covSum;
  assign metaAssert = 1'h0;
endmodule
module OptimizationBarrier_43(
  input  [53:0] io_x_ppn,
  input         io_x_d,
  input         io_x_a,
  input         io_x_g,
  input         io_x_u,
  input         io_x_x,
  input         io_x_w,
  input         io_x_r,
  input         io_x_v,
  output [53:0] io_y_ppn,
  output        io_y_d,
  output        io_y_a,
  output        io_y_g,
  output        io_y_u,
  output        io_y_x,
  output        io_y_w,
  output        io_y_r,
  output        io_y_v,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire [29:0] OptimizationBarrier_43_covSum;
  assign io_y_ppn = io_x_ppn; // @[package.scala 263:12]
  assign io_y_d = io_x_d; // @[package.scala 263:12]
  assign io_y_a = io_x_a; // @[package.scala 263:12]
  assign io_y_g = io_x_g; // @[package.scala 263:12]
  assign io_y_u = io_x_u; // @[package.scala 263:12]
  assign io_y_x = io_x_x; // @[package.scala 263:12]
  assign io_y_w = io_x_w; // @[package.scala 263:12]
  assign io_y_r = io_x_r; // @[package.scala 263:12]
  assign io_y_v = io_x_v; // @[package.scala 263:12]
  assign OptimizationBarrier_43_covSum = 30'h0;
  assign io_covSum = OptimizationBarrier_43_covSum;
  assign metaAssert = 1'h0;
endmodule
module IBuf(
  input         clock,
  input         reset,
  output        io_imem_ready,
  input         io_imem_valid,
  input         io_imem_bits_btb_taken,
  input         io_imem_bits_btb_bridx,
  input  [4:0]  io_imem_bits_btb_entry,
  input  [7:0]  io_imem_bits_btb_bht_history,
  input  [39:0] io_imem_bits_pc,
  input  [31:0] io_imem_bits_data,
  input         io_imem_bits_xcpt_pf_inst,
  input         io_imem_bits_xcpt_ae_inst,
  input         io_imem_bits_replay,
  input         io_kill,
  output [39:0] io_pc,
  output [4:0]  io_btb_resp_entry,
  output [7:0]  io_btb_resp_bht_history,
  input         io_inst_0_ready,
  output        io_inst_0_valid,
  output        io_inst_0_bits_xcpt0_pf_inst,
  output        io_inst_0_bits_xcpt0_ae_inst,
  output        io_inst_0_bits_xcpt1_pf_inst,
  output        io_inst_0_bits_xcpt1_ae_inst,
  output        io_inst_0_bits_replay,
  output        io_inst_0_bits_rvc,
  output [31:0] io_inst_0_bits_inst_bits,
  output [4:0]  io_inst_0_bits_inst_rd,
  output [4:0]  io_inst_0_bits_inst_rs1,
  output [4:0]  io_inst_0_bits_inst_rs2,
  output [4:0]  io_inst_0_bits_inst_rs3,
  output [31:0] io_inst_0_bits_raw,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  wire [31:0] exp_io_in; // @[IBuf.scala 86:21]
  wire [31:0] exp_io_out_bits; // @[IBuf.scala 86:21]
  wire [4:0] exp_io_out_rd; // @[IBuf.scala 86:21]
  wire [4:0] exp_io_out_rs1; // @[IBuf.scala 86:21]
  wire [4:0] exp_io_out_rs2; // @[IBuf.scala 86:21]
  wire [4:0] exp_io_out_rs3; // @[IBuf.scala 86:21]
  wire  exp_io_rvc; // @[IBuf.scala 86:21]
  wire [29:0] exp_io_covSum; // @[IBuf.scala 86:21]
  wire  exp_metaAssert; // @[IBuf.scala 86:21]
  reg  nBufValid; // @[IBuf.scala 34:47]
  reg [31:0] _RAND_0;
  reg [39:0] buf__pc; // @[IBuf.scala 35:16]
  reg [63:0] _RAND_1;
  reg [31:0] buf__data; // @[IBuf.scala 35:16]
  reg [31:0] _RAND_2;
  reg  buf__xcpt_pf_inst; // @[IBuf.scala 35:16]
  reg [31:0] _RAND_3;
  reg  buf__xcpt_ae_inst; // @[IBuf.scala 35:16]
  reg [31:0] _RAND_4;
  reg  buf__replay; // @[IBuf.scala 35:16]
  reg [31:0] _RAND_5;
  reg [4:0] ibufBTBResp_entry; // @[IBuf.scala 36:24]
  reg [31:0] _RAND_6;
  reg [7:0] ibufBTBResp_bht_history; // @[IBuf.scala 36:24]
  reg [31:0] _RAND_7;
  wire  pcWordBits; // @[package.scala 154:13]
  wire [1:0] _nIC_T; // @[IBuf.scala 41:64]
  wire [1:0] _nIC_T_1; // @[IBuf.scala 41:16]
  wire [1:0] _GEN_56; // @[IBuf.scala 41:88]
  wire [1:0] nIC; // @[IBuf.scala 41:88]
  wire [1:0] _nValid_T; // @[IBuf.scala 43:19]
  wire [1:0] _GEN_57; // @[IBuf.scala 43:49]
  wire [1:0] nValid; // @[IBuf.scala 43:49]
  wire [3:0] _valid_T; // @[OneHot.scala 58:35]
  wire [3:0] _valid_T_2; // @[IBuf.scala 74:33]
  wire [1:0] valid; // @[IBuf.scala 74:37]
  wire [1:0] _full_insn_T_2; // @[IBuf.scala 93:42]
  wire  _full_insn_T_4; // @[IBuf.scala 93:34]
  wire [1:0] _bufMask_T; // @[OneHot.scala 58:35]
  wire [1:0] bufMask; // @[IBuf.scala 75:37]
  wire [1:0] buf_replay; // @[IBuf.scala 77:23]
  wire  full_insn; // @[IBuf.scala 93:48]
  wire [1:0] _nReady_T_4; // @[IBuf.scala 102:71]
  wire [1:0] nReady; // @[IBuf.scala 102:56]
  wire [1:0] nICReady; // @[IBuf.scala 42:25]
  wire  _io_imem_ready_T; // @[IBuf.scala 44:47]
  wire  _io_imem_ready_T_1; // @[IBuf.scala 44:37]
  wire  _io_imem_ready_T_2; // @[IBuf.scala 44:73]
  wire [1:0] _io_imem_ready_T_4; // @[IBuf.scala 44:92]
  wire  _io_imem_ready_T_5; // @[IBuf.scala 44:85]
  wire  _io_imem_ready_T_6; // @[IBuf.scala 44:80]
  wire  _nBufValid_T_2; // @[package.scala 209:38]
  wire [1:0] _nBufValid_T_4; // @[IBuf.scala 48:65]
  wire [1:0] _nBufValid_T_5; // @[IBuf.scala 48:23]
  wire  _T_1; // @[IBuf.scala 54:27]
  wire  _T_2; // @[IBuf.scala 54:62]
  wire  _T_3; // @[IBuf.scala 54:50]
  wire  _T_7; // @[IBuf.scala 54:68]
  wire [1:0] shamt; // @[IBuf.scala 55:32]
  wire [15:0] buf_data_data_hi; // @[IBuf.scala 127:58]
  wire [63:0] buf_data_data; // @[Cat.scala 30:58]
  wire [5:0] _buf_data_T; // @[IBuf.scala 128:19]
  wire [63:0] _buf_data_T_1; // @[IBuf.scala 128:10]
  wire [39:0] _buf_pc_T_1; // @[IBuf.scala 59:35]
  wire [2:0] _buf_pc_T_2; // @[IBuf.scala 59:80]
  wire [39:0] _GEN_65; // @[IBuf.scala 59:68]
  wire [39:0] _buf_pc_T_4; // @[IBuf.scala 59:68]
  wire [39:0] _buf_pc_T_5; // @[IBuf.scala 59:109]
  wire [39:0] _buf_pc_T_6; // @[IBuf.scala 59:49]
  wire [1:0] _GEN_0; // @[IBuf.scala 54:92]
  wire [1:0] _GEN_23; // @[IBuf.scala 47:29]
  wire [1:0] _GEN_46; // @[IBuf.scala 63:20]
  wire [1:0] _icShiftAmt_T_1; // @[IBuf.scala 68:32]
  wire [1:0] icShiftAmt; // @[IBuf.scala 68:44]
  wire [15:0] icData_hi; // @[IBuf.scala 69:87]
  wire [63:0] icData_data_lo; // @[Cat.scala 30:58]
  wire [15:0] icData_data_hi; // @[IBuf.scala 120:58]
  wire [127:0] icData_data; // @[Cat.scala 30:58]
  wire [5:0] _icData_T; // @[IBuf.scala 121:19]
  wire [190:0] _GEN_68; // @[IBuf.scala 121:10]
  wire [190:0] _icData_T_1; // @[IBuf.scala 121:10]
  wire [31:0] icData; // @[package.scala 154:13]
  wire [4:0] _icMask_T_1; // @[IBuf.scala 71:65]
  wire [62:0] _icMask_T_2; // @[IBuf.scala 71:51]
  wire [31:0] icMask; // @[IBuf.scala 71:92]
  wire [31:0] _inst_T; // @[IBuf.scala 72:21]
  wire [31:0] _inst_T_2; // @[IBuf.scala 72:41]
  wire  xcpt_1_pf_inst; // @[IBuf.scala 76:53]
  wire  xcpt_1_ae_inst; // @[IBuf.scala 76:53]
  wire [1:0] _ic_replay_T_1; // @[IBuf.scala 78:63]
  wire [1:0] _ic_replay_T_2; // @[IBuf.scala 78:35]
  wire [1:0] ic_replay; // @[IBuf.scala 78:30]
  wire  _T_10; // @[IBuf.scala 79:25]
  wire  _T_11; // @[IBuf.scala 79:78]
  wire  _T_12; // @[IBuf.scala 79:52]
  wire  _T_14; // @[IBuf.scala 79:9]
  wire  _io_pc_T; // @[IBuf.scala 82:26]
  wire [1:0] _replay_T_5; // @[IBuf.scala 92:61]
  wire  _replay_T_7; // @[IBuf.scala 92:49]
  wire [1:0] _io_inst_0_bits_xcpt1_T_4; // @[IBuf.scala 96:63]
  wire [1:0] _io_inst_0_bits_xcpt1_T_5; // @[IBuf.scala 96:35]
  wire  _T_18; // @[IBuf.scala 100:25]
  wire [1:0] _T_21; // @[IBuf.scala 100:50]
  wire  _T_23; // @[IBuf.scala 100:40]
  reg [1:0] IBuf_state; // @[Register tracking IBuf state]
  reg [31:0] _RAND_8;
  reg  IBuf_cov [0:3]; // @[Coverage map for IBuf]
  reg [31:0] _RAND_9;
  wire  IBuf_cov_read_data; // @[Coverage map for IBuf]
  wire [1:0] IBuf_cov_read_addr; // @[Coverage map for IBuf]
  wire  IBuf_cov_write_data; // @[Coverage map for IBuf]
  wire [1:0] IBuf_cov_write_addr; // @[Coverage map for IBuf]
  wire  IBuf_cov_write_mask; // @[Coverage map for IBuf]
  wire  IBuf_cov_write_en; // @[Coverage map for IBuf]
  reg [29:0] IBuf_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_10;
  wire  nBufValid_shl;
  wire [1:0] nBufValid_pad;
  wire [1:0] buf__replay_shl;
  wire [1:0] buf__replay_pad;
  wire [1:0] IBuf_xor0;
  wire [29:0] exp_sum;
  wire  stopEn0;
  wire  exp_metaAssert_wire;
  wire  IBuf_or0;
  reg  IBuf_metaAssert;
  reg [31:0] _RAND_11;
  RVCExpander exp ( // @[IBuf.scala 86:21]
    .io_in(exp_io_in),
    .io_out_bits(exp_io_out_bits),
    .io_out_rd(exp_io_out_rd),
    .io_out_rs1(exp_io_out_rs1),
    .io_out_rs2(exp_io_out_rs2),
    .io_out_rs3(exp_io_out_rs3),
    .io_rvc(exp_io_rvc),
    .io_covSum(exp_io_covSum),
    .metaAssert(exp_metaAssert)
  );
  assign pcWordBits = io_imem_bits_pc[1]; // @[package.scala 154:13]
  assign _nIC_T = io_imem_bits_btb_bridx + 1'h1; // @[IBuf.scala 41:64]
  assign _nIC_T_1 = io_imem_bits_btb_taken ? _nIC_T : 2'h2; // @[IBuf.scala 41:16]
  assign _GEN_56 = {{1'd0}, pcWordBits}; // @[IBuf.scala 41:88]
  assign nIC = _nIC_T_1 - _GEN_56; // @[IBuf.scala 41:88]
  assign _nValid_T = io_imem_valid ? nIC : 2'h0; // @[IBuf.scala 43:19]
  assign _GEN_57 = {{1'd0}, nBufValid}; // @[IBuf.scala 43:49]
  assign nValid = _nValid_T + _GEN_57; // @[IBuf.scala 43:49]
  assign _valid_T = 4'h1 << nValid; // @[OneHot.scala 58:35]
  assign _valid_T_2 = _valid_T - 4'h1; // @[IBuf.scala 74:33]
  assign valid = _valid_T_2[1:0]; // @[IBuf.scala 74:37]
  assign _full_insn_T_2 = {{1'd0}, valid[1]}; // @[IBuf.scala 93:42]
  assign _full_insn_T_4 = exp_io_rvc | _full_insn_T_2[0]; // @[IBuf.scala 93:34]
  assign _bufMask_T = 2'h1 << nBufValid; // @[OneHot.scala 58:35]
  assign bufMask = _bufMask_T - 2'h1; // @[IBuf.scala 75:37]
  assign buf_replay = buf__replay ? bufMask : 2'h0; // @[IBuf.scala 77:23]
  assign full_insn = _full_insn_T_4 | buf_replay[0]; // @[IBuf.scala 93:48]
  assign _nReady_T_4 = exp_io_rvc ? 2'h1 : 2'h2; // @[IBuf.scala 102:71]
  assign nReady = full_insn ? _nReady_T_4 : 2'h0; // @[IBuf.scala 102:56]
  assign nICReady = nReady - _GEN_57; // @[IBuf.scala 42:25]
  assign _io_imem_ready_T = nReady >= _GEN_57; // @[IBuf.scala 44:47]
  assign _io_imem_ready_T_1 = io_inst_0_ready & _io_imem_ready_T; // @[IBuf.scala 44:37]
  assign _io_imem_ready_T_2 = nICReady >= nIC; // @[IBuf.scala 44:73]
  assign _io_imem_ready_T_4 = nIC - nICReady; // @[IBuf.scala 44:92]
  assign _io_imem_ready_T_5 = 2'h1 >= _io_imem_ready_T_4; // @[IBuf.scala 44:85]
  assign _io_imem_ready_T_6 = _io_imem_ready_T_2 | _io_imem_ready_T_5; // @[IBuf.scala 44:80]
  assign _nBufValid_T_2 = _io_imem_ready_T | ~nBufValid; // @[package.scala 209:38]
  assign _nBufValid_T_4 = _GEN_57 - nReady; // @[IBuf.scala 48:65]
  assign _nBufValid_T_5 = _nBufValid_T_2 ? 2'h0 : _nBufValid_T_4; // @[IBuf.scala 48:23]
  assign _T_1 = io_imem_valid & _io_imem_ready_T; // @[IBuf.scala 54:27]
  assign _T_2 = nICReady < nIC; // @[IBuf.scala 54:62]
  assign _T_3 = _T_1 & _T_2; // @[IBuf.scala 54:50]
  assign _T_7 = _T_3 & _io_imem_ready_T_5; // @[IBuf.scala 54:68]
  assign shamt = _GEN_56 + nICReady; // @[IBuf.scala 55:32]
  assign buf_data_data_hi = io_imem_bits_data[31:16]; // @[IBuf.scala 127:58]
  assign buf_data_data = {buf_data_data_hi,buf_data_data_hi,io_imem_bits_data}; // @[Cat.scala 30:58]
  assign _buf_data_T = {shamt, 4'h0}; // @[IBuf.scala 128:19]
  assign _buf_data_T_1 = buf_data_data >> _buf_data_T; // @[IBuf.scala 128:10]
  assign _buf_pc_T_1 = io_imem_bits_pc & 40'hfffffffffc; // @[IBuf.scala 59:35]
  assign _buf_pc_T_2 = {nICReady, 1'h0}; // @[IBuf.scala 59:80]
  assign _GEN_65 = {{37'd0}, _buf_pc_T_2}; // @[IBuf.scala 59:68]
  assign _buf_pc_T_4 = io_imem_bits_pc + _GEN_65; // @[IBuf.scala 59:68]
  assign _buf_pc_T_5 = _buf_pc_T_4 & 40'h3; // @[IBuf.scala 59:109]
  assign _buf_pc_T_6 = _buf_pc_T_1 | _buf_pc_T_5; // @[IBuf.scala 59:49]
  assign _GEN_0 = _T_7 ? _io_imem_ready_T_4 : _nBufValid_T_5; // @[IBuf.scala 54:92]
  assign _GEN_23 = io_inst_0_ready ? _GEN_0 : {{1'd0}, nBufValid}; // @[IBuf.scala 47:29]
  assign _GEN_46 = io_kill ? 2'h0 : _GEN_23; // @[IBuf.scala 63:20]
  assign _icShiftAmt_T_1 = 2'h2 + _GEN_57; // @[IBuf.scala 68:32]
  assign icShiftAmt = _icShiftAmt_T_1 - _GEN_56; // @[IBuf.scala 68:44]
  assign icData_hi = io_imem_bits_data[15:0]; // @[IBuf.scala 69:87]
  assign icData_data_lo = {io_imem_bits_data,icData_hi,icData_hi}; // @[Cat.scala 30:58]
  assign icData_data_hi = icData_data_lo[63:48]; // @[IBuf.scala 120:58]
  assign icData_data = {icData_data_hi,icData_data_hi,icData_data_hi,icData_data_hi,io_imem_bits_data,icData_hi,icData_hi}; // @[Cat.scala 30:58]
  assign _icData_T = {icShiftAmt, 4'h0}; // @[IBuf.scala 121:19]
  assign _GEN_68 = {{63'd0}, icData_data}; // @[IBuf.scala 121:10]
  assign _icData_T_1 = _GEN_68 << _icData_T; // @[IBuf.scala 121:10]
  assign icData = _icData_T_1[95:64]; // @[package.scala 154:13]
  assign _icMask_T_1 = {nBufValid, 4'h0}; // @[IBuf.scala 71:65]
  assign _icMask_T_2 = 63'hffffffff << _icMask_T_1; // @[IBuf.scala 71:51]
  assign icMask = _icMask_T_2[31:0]; // @[IBuf.scala 71:92]
  assign _inst_T = icData & icMask; // @[IBuf.scala 72:21]
  assign _inst_T_2 = buf__data & ~icMask; // @[IBuf.scala 72:41]
  assign xcpt_1_pf_inst = bufMask[1] ? buf__xcpt_pf_inst : io_imem_bits_xcpt_pf_inst; // @[IBuf.scala 76:53]
  assign xcpt_1_ae_inst = bufMask[1] ? buf__xcpt_ae_inst : io_imem_bits_xcpt_ae_inst; // @[IBuf.scala 76:53]
  assign _ic_replay_T_1 = valid & ~bufMask; // @[IBuf.scala 78:63]
  assign _ic_replay_T_2 = io_imem_bits_replay ? _ic_replay_T_1 : 2'h0; // @[IBuf.scala 78:35]
  assign ic_replay = buf_replay | _ic_replay_T_2; // @[IBuf.scala 78:30]
  assign _T_10 = ~io_imem_valid | ~io_imem_bits_btb_taken; // @[IBuf.scala 79:25]
  assign _T_11 = io_imem_bits_btb_bridx >= pcWordBits; // @[IBuf.scala 79:78]
  assign _T_12 = _T_10 | _T_11; // @[IBuf.scala 79:52]
  assign _T_14 = _T_12 | reset; // @[IBuf.scala 79:9]
  assign _io_pc_T = nBufValid > 1'h0; // @[IBuf.scala 82:26]
  assign _replay_T_5 = {{1'd0}, ic_replay[1]}; // @[IBuf.scala 92:61]
  assign _replay_T_7 = ~exp_io_rvc & _replay_T_5[0]; // @[IBuf.scala 92:49]
  assign _io_inst_0_bits_xcpt1_T_4 = {xcpt_1_pf_inst,xcpt_1_ae_inst}; // @[IBuf.scala 96:63]
  assign _io_inst_0_bits_xcpt1_T_5 = exp_io_rvc ? 2'h0 : _io_inst_0_bits_xcpt1_T_4; // @[IBuf.scala 96:35]
  assign _T_18 = bufMask[0] & exp_io_rvc; // @[IBuf.scala 100:25]
  assign _T_21 = {{1'd0}, bufMask[1]}; // @[IBuf.scala 100:50]
  assign _T_23 = _T_18 | _T_21[0]; // @[IBuf.scala 100:40]
  assign io_imem_ready = _io_imem_ready_T_1 & _io_imem_ready_T_6; // @[IBuf.scala 44:17]
  assign io_pc = _io_pc_T ? buf__pc : io_imem_bits_pc; // @[IBuf.scala 82:9]
  assign io_btb_resp_entry = _T_23 ? ibufBTBResp_entry : io_imem_bits_btb_entry; // @[IBuf.scala 81:15 IBuf.scala 100:71]
  assign io_btb_resp_bht_history = _T_23 ? ibufBTBResp_bht_history : io_imem_bits_btb_bht_history; // @[IBuf.scala 81:15 IBuf.scala 100:71]
  assign io_inst_0_valid = valid[0] & full_insn; // @[IBuf.scala 94:24]
  assign io_inst_0_bits_xcpt0_pf_inst = bufMask[0] ? buf__xcpt_pf_inst : io_imem_bits_xcpt_pf_inst; // @[IBuf.scala 95:29]
  assign io_inst_0_bits_xcpt0_ae_inst = bufMask[0] ? buf__xcpt_ae_inst : io_imem_bits_xcpt_ae_inst; // @[IBuf.scala 95:29]
  assign io_inst_0_bits_xcpt1_pf_inst = _io_inst_0_bits_xcpt1_T_5[1]; // @[IBuf.scala 96:29]
  assign io_inst_0_bits_xcpt1_ae_inst = _io_inst_0_bits_xcpt1_T_5[0]; // @[IBuf.scala 96:29]
  assign io_inst_0_bits_replay = ic_replay[0] | _replay_T_7; // @[IBuf.scala 97:30]
  assign io_inst_0_bits_rvc = exp_io_rvc; // @[IBuf.scala 98:27]
  assign io_inst_0_bits_inst_bits = exp_io_out_bits; // @[IBuf.scala 88:26]
  assign io_inst_0_bits_inst_rd = exp_io_out_rd; // @[IBuf.scala 88:26]
  assign io_inst_0_bits_inst_rs1 = exp_io_out_rs1; // @[IBuf.scala 88:26]
  assign io_inst_0_bits_inst_rs2 = exp_io_out_rs2; // @[IBuf.scala 88:26]
  assign io_inst_0_bits_inst_rs3 = exp_io_out_rs3; // @[IBuf.scala 88:26]
  assign io_inst_0_bits_raw = _inst_T | _inst_T_2; // @[IBuf.scala 89:25]
  assign exp_io_in = _inst_T | _inst_T_2; // @[IBuf.scala 87:15]
  assign IBuf_cov_read_addr = IBuf_state;
  assign IBuf_cov_read_data = IBuf_cov[IBuf_cov_read_addr]; // @[Coverage map for IBuf]
  assign IBuf_cov_write_data = 1'h1;
  assign IBuf_cov_write_addr = IBuf_state;
  assign IBuf_cov_write_mask = 1'h1;
  assign IBuf_cov_write_en = 1'h1;
  assign nBufValid_shl = nBufValid;
  assign nBufValid_pad = {1'h0,nBufValid_shl};
  assign buf__replay_shl = {buf__replay, 1'h0};
  assign buf__replay_pad = buf__replay_shl;
  assign IBuf_xor0 = nBufValid_pad ^ buf__replay_pad;
  assign exp_sum = IBuf_covSum + exp_io_covSum;
  assign io_covSum = exp_sum;
  assign stopEn0 = ~_T_14;
  assign exp_metaAssert_wire = exp_metaAssert;
  assign IBuf_or0 = stopEn0 | exp_metaAssert_wire;
  assign metaAssert = IBuf_metaAssert;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  nBufValid = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {2{`RANDOM}};
  buf__pc = _RAND_1[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  buf__data = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  buf__xcpt_pf_inst = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  buf__xcpt_ae_inst = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  buf__replay = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  ibufBTBResp_entry = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  ibufBTBResp_bht_history = _RAND_7[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  IBuf_state = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    IBuf_cov[initvar] = _RAND_9[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  IBuf_covSum = _RAND_10[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  IBuf_metaAssert = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      nBufValid <= 1'h0;
    end else if (reset) begin
      nBufValid <= 1'h0;
    end else begin
      nBufValid <= _GEN_46[0];
    end
    if (metaReset) begin
      buf__pc <= 40'h0;
    end else if (io_inst_0_ready) begin
      if (_T_7) begin
        buf__pc <= _buf_pc_T_6;
      end
    end
    if (metaReset) begin
      buf__data <= 32'h0;
    end else if (io_inst_0_ready) begin
      if (_T_7) begin
        buf__data <= {{16'd0}, _buf_data_T_1[15:0]};
      end
    end
    if (metaReset) begin
      buf__xcpt_pf_inst <= 1'h0;
    end else if (io_inst_0_ready) begin
      if (_T_7) begin
        buf__xcpt_pf_inst <= io_imem_bits_xcpt_pf_inst;
      end
    end
    if (metaReset) begin
      buf__xcpt_ae_inst <= 1'h0;
    end else if (io_inst_0_ready) begin
      if (_T_7) begin
        buf__xcpt_ae_inst <= io_imem_bits_xcpt_ae_inst;
      end
    end
    if (metaReset) begin
      buf__replay <= 1'h0;
    end else if (io_inst_0_ready) begin
      if (_T_7) begin
        buf__replay <= io_imem_bits_replay;
      end
    end
    if (metaReset) begin
      ibufBTBResp_entry <= 5'h0;
    end else if (io_inst_0_ready) begin
      if (_T_7) begin
        ibufBTBResp_entry <= io_imem_bits_btb_entry;
      end
    end
    if (metaReset) begin
      ibufBTBResp_bht_history <= 8'h0;
    end else if (io_inst_0_ready) begin
      if (_T_7) begin
        ibufBTBResp_bht_history <= io_imem_bits_btb_bht_history;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_14) begin
          $fwrite(32'h80000002,"Assertion failed\n    at IBuf.scala:79 assert(!io.imem.valid || !io.imem.bits.btb.taken || io.imem.bits.btb.bridx >= pcWordBits)\n"); // @[IBuf.scala 79:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_14) begin
          $fatal; // @[IBuf.scala 79:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    IBuf_state <= IBuf_xor0;
    if (!(IBuf_cov_read_data)) begin
      IBuf_covSum <= IBuf_covSum + 1'h1;
    end
    if (metaReset) begin
      IBuf_metaAssert <= 1'h0;
    end else begin
      IBuf_metaAssert <= IBuf_metaAssert | IBuf_or0;
    end
  end
  always @(posedge clock) begin
    if(IBuf_cov_write_en & IBuf_cov_write_mask) begin
      IBuf_cov[IBuf_cov_write_addr] <= IBuf_cov_write_data; // @[Coverage map for IBuf]
    end
  end
endmodule
module CSRFile(
  input         clock,
  input         reset,
  input         io_ungated_clock,
  input         io_interrupts_debug,
  input         io_interrupts_mtip,
  input         io_interrupts_msip,
  input         io_interrupts_meip,
  input         io_interrupts_seip,
  input         io_hartid,
  input  [11:0] io_rw_addr,
  input  [2:0]  io_rw_cmd,
  output [63:0] io_rw_rdata,
  input  [63:0] io_rw_wdata,
  input  [11:0] io_decode_0_csr,
  output        io_decode_0_fp_illegal,
  output        io_decode_0_fp_csr,
  output        io_decode_0_read_illegal,
  output        io_decode_0_write_illegal,
  output        io_decode_0_write_flush,
  output        io_decode_0_system_illegal,
  output        io_csr_stall,
  output        io_eret,
  output        io_singleStep,
  output        io_status_debug,
  output        io_status_cease,
  output        io_status_wfi,
  output [31:0] io_status_isa,
  output [1:0]  io_status_dprv,
  output [1:0]  io_status_prv,
  output        io_status_sd,
  output [26:0] io_status_zero2,
  output [1:0]  io_status_sxl,
  output [1:0]  io_status_uxl,
  output        io_status_sd_rv32,
  output [7:0]  io_status_zero1,
  output        io_status_tsr,
  output        io_status_tw,
  output        io_status_tvm,
  output        io_status_mxr,
  output        io_status_sum,
  output        io_status_mprv,
  output [1:0]  io_status_xs,
  output [1:0]  io_status_fs,
  output [1:0]  io_status_mpp,
  output [1:0]  io_status_vs,
  output        io_status_spp,
  output        io_status_mpie,
  output        io_status_hpie,
  output        io_status_spie,
  output        io_status_upie,
  output        io_status_mie,
  output        io_status_hie,
  output        io_status_sie,
  output        io_status_uie,
  output [3:0]  io_ptbr_mode,
  output [43:0] io_ptbr_ppn,
  output [39:0] io_evec,
  input         io_exception,
  input         io_retire,
  input  [63:0] io_cause,
  input  [39:0] io_pc,
  input  [39:0] io_tval,
  output [63:0] io_time,
  output [2:0]  io_fcsr_rm,
  input         io_fcsr_flags_valid,
  input  [4:0]  io_fcsr_flags_bits,
  output        io_interrupt,
  output [63:0] io_interrupt_cause,
  output        io_bp_0_control_action,
  output [1:0]  io_bp_0_control_tmatch,
  output        io_bp_0_control_m,
  output        io_bp_0_control_s,
  output        io_bp_0_control_u,
  output        io_bp_0_control_x,
  output        io_bp_0_control_w,
  output        io_bp_0_control_r,
  output [38:0] io_bp_0_address,
  output        io_pmp_0_cfg_l,
  output [1:0]  io_pmp_0_cfg_a,
  output        io_pmp_0_cfg_x,
  output        io_pmp_0_cfg_w,
  output        io_pmp_0_cfg_r,
  output [29:0] io_pmp_0_addr,
  output [31:0] io_pmp_0_mask,
  output        io_pmp_1_cfg_l,
  output [1:0]  io_pmp_1_cfg_a,
  output        io_pmp_1_cfg_x,
  output        io_pmp_1_cfg_w,
  output        io_pmp_1_cfg_r,
  output [29:0] io_pmp_1_addr,
  output [31:0] io_pmp_1_mask,
  output        io_pmp_2_cfg_l,
  output [1:0]  io_pmp_2_cfg_a,
  output        io_pmp_2_cfg_x,
  output        io_pmp_2_cfg_w,
  output        io_pmp_2_cfg_r,
  output [29:0] io_pmp_2_addr,
  output [31:0] io_pmp_2_mask,
  output        io_pmp_3_cfg_l,
  output [1:0]  io_pmp_3_cfg_a,
  output        io_pmp_3_cfg_x,
  output        io_pmp_3_cfg_w,
  output        io_pmp_3_cfg_r,
  output [29:0] io_pmp_3_addr,
  output [31:0] io_pmp_3_mask,
  output        io_pmp_4_cfg_l,
  output [1:0]  io_pmp_4_cfg_a,
  output        io_pmp_4_cfg_x,
  output        io_pmp_4_cfg_w,
  output        io_pmp_4_cfg_r,
  output [29:0] io_pmp_4_addr,
  output [31:0] io_pmp_4_mask,
  output        io_pmp_5_cfg_l,
  output [1:0]  io_pmp_5_cfg_a,
  output        io_pmp_5_cfg_x,
  output        io_pmp_5_cfg_w,
  output        io_pmp_5_cfg_r,
  output [29:0] io_pmp_5_addr,
  output [31:0] io_pmp_5_mask,
  output        io_pmp_6_cfg_l,
  output [1:0]  io_pmp_6_cfg_a,
  output        io_pmp_6_cfg_x,
  output        io_pmp_6_cfg_w,
  output        io_pmp_6_cfg_r,
  output [29:0] io_pmp_6_addr,
  output [31:0] io_pmp_6_mask,
  output        io_pmp_7_cfg_l,
  output [1:0]  io_pmp_7_cfg_a,
  output        io_pmp_7_cfg_x,
  output        io_pmp_7_cfg_w,
  output        io_pmp_7_cfg_r,
  output [29:0] io_pmp_7_addr,
  output [31:0] io_pmp_7_mask,
  output        io_inhibit_cycle,
  input  [31:0] io_inst_0,
  output        io_trace_0_valid,
  output [39:0] io_trace_0_iaddr,
  output [31:0] io_trace_0_insn,
  output [2:0]  io_trace_0_priv,
  output        io_trace_0_exception,
  output        io_trace_0_interrupt,
  output [63:0] io_trace_0_cause,
  output [39:0] io_trace_0_tval,
  output [63:0] io_customCSRs_0_value,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  reg rv_dv; //SC_added to identify DV test and CP
  reg [1:0] reg_mstatus_prv; // @[CSR.scala 319:24]
  reg [31:0] _RAND_0;
  reg  reg_mstatus_tsr; // @[CSR.scala 319:24]
  reg [31:0] _RAND_1;
  reg  reg_mstatus_tw; // @[CSR.scala 319:24]
  reg [31:0] _RAND_2;
  reg  reg_mstatus_tvm; // @[CSR.scala 319:24]
  reg [31:0] _RAND_3;
  reg  reg_mstatus_mxr; // @[CSR.scala 319:24]
  reg [31:0] _RAND_4;
  reg  reg_mstatus_sum; // @[CSR.scala 319:24]
  reg [31:0] _RAND_5;
  reg  reg_mstatus_mprv; // @[CSR.scala 319:24]
  reg [31:0] _RAND_6;
  reg [1:0] reg_mstatus_fs; // @[CSR.scala 319:24]
  reg [31:0] _RAND_7;
  reg [1:0] reg_mstatus_mpp; // @[CSR.scala 319:24]
  reg [31:0] _RAND_8;
  reg  reg_mstatus_spp; // @[CSR.scala 319:24]
  reg [31:0] _RAND_9;
  reg  reg_mstatus_mpie; // @[CSR.scala 319:24]
  reg [31:0] _RAND_10;
  reg  reg_mstatus_spie; // @[CSR.scala 319:24]
  reg [31:0] _RAND_11;
  reg  reg_mstatus_mie; // @[CSR.scala 319:24]
  reg [31:0] _RAND_12;
  reg  reg_mstatus_sie; // @[CSR.scala 319:24]
  reg [31:0] _RAND_13;
  wire  system_insn; // @[CSR.scala 639:31]
  wire [31:0] _T_192; // @[CSR.scala 652:28]
  wire [31:0] _T_199; // @[Decode.scala 14:65]
  wire  _T_200; // @[Decode.scala 14:121]
  wire [31:0] _T_201; // @[Decode.scala 14:65]
  wire  _T_202; // @[Decode.scala 14:121]
  wire  _T_204; // @[Decode.scala 15:30]
  wire  insn_ret; // @[CSR.scala 652:95]
  wire  _T_406; // @[CSR.scala 821:52]
  reg [1:0] reg_dcsr_prv; // @[CSR.scala 327:21]
  reg [31:0] _RAND_14;
  wire [1:0] _GEN_149; // @[CSR.scala 821:70]
  wire [1:0] ret_prv; // @[CSR.scala 815:52]
  wire [31:0] _T_193; // @[Decode.scala 14:65]
  wire  _T_194; // @[Decode.scala 14:121]
  wire  insn_call; // @[CSR.scala 652:95]
  wire  _T_197; // @[Decode.scala 14:121]
  wire  insn_break; // @[CSR.scala 652:95]
  wire  _exception_T; // @[CSR.scala 738:29]
  wire  exception; // @[CSR.scala 738:43]
  reg  reg_singleStepped; // @[CSR.scala 372:30]
  reg [31:0] _RAND_15;
  wire [3:0] _GEN_20; // @[CSR.scala 688:36]
  wire [3:0] _cause_T_1; // @[CSR.scala 688:36]
  wire [63:0] _cause_T_2; // @[CSR.scala 689:14]
  wire [63:0] cause; // @[CSR.scala 688:8]
  wire [7:0] cause_lsbs; // @[CSR.scala 690:25]
  wire  _causeIsDebugInt_T_1; // @[CSR.scala 691:53]
  wire  causeIsDebugInt; // @[CSR.scala 691:39]
  wire  _trapToDebug_T; // @[CSR.scala 694:60]
  wire  causeIsDebugTrigger; // @[CSR.scala 692:44]
  wire  _trapToDebug_T_1; // @[CSR.scala 694:79]
  wire  _causeIsDebugBreak_T_2; // @[CSR.scala 693:42]
  reg  reg_dcsr_ebreakm; // @[CSR.scala 327:21]
  reg [31:0] _RAND_16;
  reg  reg_dcsr_ebreaks; // @[CSR.scala 327:21]
  reg [31:0] _RAND_17;
  reg  reg_dcsr_ebreaku; // @[CSR.scala 327:21]
  reg [31:0] _RAND_18;
  wire [3:0] _causeIsDebugBreak_T_3; // @[Cat.scala 30:58]
  wire [3:0] _causeIsDebugBreak_T_4; // @[CSR.scala 693:134]
  wire  causeIsDebugBreak; // @[CSR.scala 693:56]
  wire  _trapToDebug_T_2; // @[CSR.scala 694:102]
  reg  reg_debug; // @[CSR.scala 368:22]
  reg [31:0] _RAND_19;
  wire  trapToDebug; // @[CSR.scala 694:123]
  wire [1:0] _GEN_56; // @[CSR.scala 756:25]
  reg  reg_rnmie; // @[CSR.scala 407:26]
  reg [31:0] _RAND_20;
  reg  reg_unmie; // @[CSR.scala 408:26]
  reg [31:0] _RAND_21;
  wire  _delegate_T; // @[CSR.scala 698:59]
  reg [63:0] reg_mideleg; // @[CSR.scala 383:18]
  reg [63:0] _RAND_22;
  wire [63:0] read_mideleg; // @[CSR.scala 384:36]
  wire [63:0] _delegate_T_3; // @[CSR.scala 698:102]
  reg [63:0] reg_medeleg; // @[CSR.scala 387:18]
  reg [63:0] _RAND_23;
  wire [63:0] read_medeleg; // @[CSR.scala 388:36]
  wire [63:0] _delegate_T_5; // @[CSR.scala 698:128]
  wire  _delegate_T_7; // @[CSR.scala 698:74]
  wire  delegate; // @[CSR.scala 698:68]
  wire  nmie; // @[CSR.scala 409:24]
  wire  _T_279; // @[CSR.scala 772:26]
  wire [1:0] _GEN_70; // @[CSR.scala 772:35]
  wire [1:0] _GEN_100; // @[CSR.scala 755:24]
  wire [1:0] _GEN_123; // @[CSR.scala 754:20]
  wire [1:0] new_prv; // @[CSR.scala 813:19]
  wire  _reg_mstatus_prv_T; // @[CSR.scala 1190:35]
  reg [2:0] reg_dcsr_cause; // @[CSR.scala 327:21]
  reg [31:0] _RAND_24;
  reg  reg_dcsr_step; // @[CSR.scala 327:21]
  reg [31:0] _RAND_25;
  reg [39:0] reg_dpc; // @[CSR.scala 369:20]
  reg [63:0] _RAND_26;
  reg [63:0] reg_dscratch; // @[CSR.scala 370:25]
  reg [63:0] _RAND_27;
  reg  reg_bp_0_control_dmode; // @[CSR.scala 378:19]
  reg [31:0] _RAND_28;
  reg  reg_bp_0_control_action; // @[CSR.scala 378:19]
  reg [31:0] _RAND_29;
  reg [1:0] reg_bp_0_control_tmatch; // @[CSR.scala 378:19]
  reg [31:0] _RAND_30;
  reg  reg_bp_0_control_m; // @[CSR.scala 378:19]
  reg [31:0] _RAND_31;
  reg  reg_bp_0_control_s; // @[CSR.scala 378:19]
  reg [31:0] _RAND_32;
  reg  reg_bp_0_control_u; // @[CSR.scala 378:19]
  reg [31:0] _RAND_33;
  reg  reg_bp_0_control_x; // @[CSR.scala 378:19]
  reg [31:0] _RAND_34;
  reg  reg_bp_0_control_w; // @[CSR.scala 378:19]
  reg [31:0] _RAND_35;
  reg  reg_bp_0_control_r; // @[CSR.scala 378:19]
  reg [31:0] _RAND_36;
  reg [38:0] reg_bp_0_address; // @[CSR.scala 378:19]
  reg [63:0] _RAND_37;
  reg  reg_pmp_0_cfg_l; // @[CSR.scala 379:20]
  reg [31:0] _RAND_38;
  reg [1:0] reg_pmp_0_cfg_a; // @[CSR.scala 379:20]
  reg [31:0] _RAND_39;
  reg  reg_pmp_0_cfg_x; // @[CSR.scala 379:20]
  reg [31:0] _RAND_40;
  reg  reg_pmp_0_cfg_w; // @[CSR.scala 379:20]
  reg [31:0] _RAND_41;
  reg  reg_pmp_0_cfg_r; // @[CSR.scala 379:20]
  reg [31:0] _RAND_42;
  reg [29:0] reg_pmp_0_addr; // @[CSR.scala 379:20]
  reg [31:0] _RAND_43;
  reg  reg_pmp_1_cfg_l; // @[CSR.scala 379:20]
  reg [31:0] _RAND_44;
  reg [1:0] reg_pmp_1_cfg_a; // @[CSR.scala 379:20]
  reg [31:0] _RAND_45;
  reg  reg_pmp_1_cfg_x; // @[CSR.scala 379:20]
  reg [31:0] _RAND_46;
  reg  reg_pmp_1_cfg_w; // @[CSR.scala 379:20]
  reg [31:0] _RAND_47;
  reg  reg_pmp_1_cfg_r; // @[CSR.scala 379:20]
  reg [31:0] _RAND_48;
  reg [29:0] reg_pmp_1_addr; // @[CSR.scala 379:20]
  reg [31:0] _RAND_49;
  reg  reg_pmp_2_cfg_l; // @[CSR.scala 379:20]
  reg [31:0] _RAND_50;
  reg [1:0] reg_pmp_2_cfg_a; // @[CSR.scala 379:20]
  reg [31:0] _RAND_51;
  reg  reg_pmp_2_cfg_x; // @[CSR.scala 379:20]
  reg [31:0] _RAND_52;
  reg  reg_pmp_2_cfg_w; // @[CSR.scala 379:20]
  reg [31:0] _RAND_53;
  reg  reg_pmp_2_cfg_r; // @[CSR.scala 379:20]
  reg [31:0] _RAND_54;
  reg [29:0] reg_pmp_2_addr; // @[CSR.scala 379:20]
  reg [31:0] _RAND_55;
  reg  reg_pmp_3_cfg_l; // @[CSR.scala 379:20]
  reg [31:0] _RAND_56;
  reg [1:0] reg_pmp_3_cfg_a; // @[CSR.scala 379:20]
  reg [31:0] _RAND_57;
  reg  reg_pmp_3_cfg_x; // @[CSR.scala 379:20]
  reg [31:0] _RAND_58;
  reg  reg_pmp_3_cfg_w; // @[CSR.scala 379:20]
  reg [31:0] _RAND_59;
  reg  reg_pmp_3_cfg_r; // @[CSR.scala 379:20]
  reg [31:0] _RAND_60;
  reg [29:0] reg_pmp_3_addr; // @[CSR.scala 379:20]
  reg [31:0] _RAND_61;
  reg  reg_pmp_4_cfg_l; // @[CSR.scala 379:20]
  reg [31:0] _RAND_62;
  reg [1:0] reg_pmp_4_cfg_a; // @[CSR.scala 379:20]
  reg [31:0] _RAND_63;
  reg  reg_pmp_4_cfg_x; // @[CSR.scala 379:20]
  reg [31:0] _RAND_64;
  reg  reg_pmp_4_cfg_w; // @[CSR.scala 379:20]
  reg [31:0] _RAND_65;
  reg  reg_pmp_4_cfg_r; // @[CSR.scala 379:20]
  reg [31:0] _RAND_66;
  reg [29:0] reg_pmp_4_addr; // @[CSR.scala 379:20]
  reg [31:0] _RAND_67;
  reg  reg_pmp_5_cfg_l; // @[CSR.scala 379:20]
  reg [31:0] _RAND_68;
  reg [1:0] reg_pmp_5_cfg_a; // @[CSR.scala 379:20]
  reg [31:0] _RAND_69;
  reg  reg_pmp_5_cfg_x; // @[CSR.scala 379:20]
  reg [31:0] _RAND_70;
  reg  reg_pmp_5_cfg_w; // @[CSR.scala 379:20]
  reg [31:0] _RAND_71;
  reg  reg_pmp_5_cfg_r; // @[CSR.scala 379:20]
  reg [31:0] _RAND_72;
  reg [29:0] reg_pmp_5_addr; // @[CSR.scala 379:20]
  reg [31:0] _RAND_73;
  reg  reg_pmp_6_cfg_l; // @[CSR.scala 379:20]
  reg [31:0] _RAND_74;
  reg [1:0] reg_pmp_6_cfg_a; // @[CSR.scala 379:20]
  reg [31:0] _RAND_75;
  reg  reg_pmp_6_cfg_x; // @[CSR.scala 379:20]
  reg [31:0] _RAND_76;
  reg  reg_pmp_6_cfg_w; // @[CSR.scala 379:20]
  reg [31:0] _RAND_77;
  reg  reg_pmp_6_cfg_r; // @[CSR.scala 379:20]
  reg [31:0] _RAND_78;
  reg [29:0] reg_pmp_6_addr; // @[CSR.scala 379:20]
  reg [31:0] _RAND_79;
  reg  reg_pmp_7_cfg_l; // @[CSR.scala 379:20]
  reg [31:0] _RAND_80;
  reg [1:0] reg_pmp_7_cfg_a; // @[CSR.scala 379:20]
  reg [31:0] _RAND_81;
  reg  reg_pmp_7_cfg_x; // @[CSR.scala 379:20]
  reg [31:0] _RAND_82;
  reg  reg_pmp_7_cfg_w; // @[CSR.scala 379:20]
  reg [31:0] _RAND_83;
  reg  reg_pmp_7_cfg_r; // @[CSR.scala 379:20]
  reg [31:0] _RAND_84;
  reg [29:0] reg_pmp_7_addr; // @[CSR.scala 379:20]
  reg [31:0] _RAND_85;
  reg [63:0] reg_mie; // @[CSR.scala 381:20]
  reg [63:0] _RAND_86;
  reg  reg_mip_seip; // @[CSR.scala 390:20]
  reg [31:0] _RAND_87;
  reg  reg_mip_stip; // @[CSR.scala 390:20]
  reg [31:0] _RAND_88;
  reg  reg_mip_ssip; // @[CSR.scala 390:20]
  reg [31:0] _RAND_89;
  reg [39:0] reg_mepc; // @[CSR.scala 391:21]
  reg [63:0] _RAND_90;
  reg [63:0] reg_mcause; // @[CSR.scala 392:27]
  reg [63:0] _RAND_91;
  reg [39:0] reg_mtval; // @[CSR.scala 393:22]
  reg [63:0] _RAND_92;
  reg [63:0] reg_mscratch; // @[CSR.scala 394:25]
  reg [63:0] _RAND_93;
  reg [31:0] reg_mtvec; // @[CSR.scala 397:27]
  reg [31:0] _RAND_94;
  reg [31:0] reg_mcounteren; // @[CSR.scala 413:18]
  reg [31:0] _RAND_95;
  wire [31:0] read_mcounteren; // @[CSR.scala 414:30]
  reg [31:0] reg_scounteren; // @[CSR.scala 417:18]
  reg [31:0] _RAND_96;
  wire [31:0] read_scounteren; // @[CSR.scala 418:36]
  reg [39:0] reg_sepc; // @[CSR.scala 421:21]
  reg [63:0] _RAND_97;
  reg [63:0] reg_scause; // @[CSR.scala 422:23]
  reg [63:0] _RAND_98;
  reg [39:0] reg_stval; // @[CSR.scala 423:22]
  reg [63:0] _RAND_99;
  reg [63:0] reg_sscratch; // @[CSR.scala 424:25]
  reg [63:0] _RAND_100;
  reg [38:0] reg_stvec; // @[CSR.scala 425:22]
  reg [63:0] _RAND_101;
  reg [3:0] reg_satp_mode; // @[CSR.scala 426:21]
  reg [31:0] _RAND_102;
  reg [43:0] reg_satp_ppn; // @[CSR.scala 426:21]
  reg [63:0] _RAND_103;
  reg  reg_wfi; // @[CSR.scala 427:50]
  reg [31:0] _RAND_104;
  reg [4:0] reg_fflags; // @[CSR.scala 429:23]
  reg [31:0] _RAND_105;
  reg [2:0] reg_frm; // @[CSR.scala 430:20]
  reg [31:0] _RAND_106;
  reg [2:0] reg_mcountinhibit; // @[CSR.scala 436:34]
  reg [31:0] _RAND_107;
  wire  x67; // @[CSR.scala 438:75]
  reg [5:0] value_lo; // @[Counters.scala 45:37]
  reg [31:0] _RAND_108;
  wire [5:0] _GEN_23; // @[Counters.scala 46:33]
  wire [6:0] nextSmall; // @[Counters.scala 46:33]
  wire [6:0] _GEN_0; // @[Counters.scala 47:19]
  reg [57:0] value_hi; // @[Counters.scala 50:27]
  reg [63:0] _RAND_109;
  wire  _large_T_2; // @[Counters.scala 51:33]
  wire [57:0] _large_r_T_1; // @[Counters.scala 51:55]
  wire [63:0] value; // @[Cat.scala 30:58]
  reg [5:0] value_lo_1; // @[Counters.scala 45:37]
  reg [31:0] _RAND_110;
  wire [6:0] nextSmall_1; // @[Counters.scala 46:33]
  wire [6:0] _GEN_2; // @[Counters.scala 47:19]
  reg [57:0] value_hi_1; // @[Counters.scala 50:27]
  reg [63:0] _RAND_111;
  wire  _large_T_5; // @[Counters.scala 51:33]
  wire [57:0] _large_r_T_3; // @[Counters.scala 51:55]
  wire [63:0] value_1; // @[Cat.scala 30:58]
  wire  mip_seip; // @[CSR.scala 452:57]
  wire [7:0] read_mip_lo; // @[CSR.scala 454:22]
  wire [15:0] _read_mip_T; // @[CSR.scala 454:22]
  wire [15:0] read_mip; // @[CSR.scala 454:29]
  wire [63:0] _GEN_45; // @[CSR.scala 457:56]
  wire [63:0] pending_interrupts; // @[CSR.scala 457:56]
  wire [14:0] d_interrupts; // @[CSR.scala 458:42]
  wire  _m_interrupts_T_1; // @[CSR.scala 464:60]
  wire  _m_interrupts_T_2; // @[CSR.scala 464:31]
  wire [63:0] _m_interrupts_T_4; // @[CSR.scala 464:103]
  wire [63:0] m_interrupts; // @[CSR.scala 464:25]
  wire  _s_interrupts_T; // @[CSR.scala 465:51]
  wire  _s_interrupts_T_1; // @[CSR.scala 465:79]
  wire  _s_interrupts_T_2; // @[CSR.scala 465:89]
  wire  _s_interrupts_T_3; // @[CSR.scala 465:59]
  wire  _s_interrupts_T_4; // @[CSR.scala 465:31]
  wire [63:0] _s_interrupts_T_5; // @[CSR.scala 465:130]
  wire [63:0] s_interrupts; // @[CSR.scala 465:25]
  wire  _any_T_38; // @[CSR.scala 1180:90]
  wire  _any_T_39; // @[CSR.scala 1180:90]
  wire  _any_T_40; // @[CSR.scala 1180:90]
  wire  _any_T_41; // @[CSR.scala 1180:90]
  wire  _any_T_42; // @[CSR.scala 1180:90]
  wire  _any_T_43; // @[CSR.scala 1180:90]
  wire  _any_T_44; // @[CSR.scala 1180:90]
  wire  _any_T_45; // @[CSR.scala 1180:90]
  wire  _any_T_46; // @[CSR.scala 1180:90]
  wire  _any_T_47; // @[CSR.scala 1180:90]
  wire  _any_T_48; // @[CSR.scala 1180:90]
  wire  _any_T_50; // @[CSR.scala 1180:90]
  wire  _any_T_51; // @[CSR.scala 1180:90]
  wire  _any_T_52; // @[CSR.scala 1180:90]
  wire  _any_T_53; // @[CSR.scala 1180:90]
  wire  _any_T_54; // @[CSR.scala 1180:90]
  wire  _any_T_55; // @[CSR.scala 1180:90]
  wire  _any_T_56; // @[CSR.scala 1180:90]
  wire  _any_T_57; // @[CSR.scala 1180:90]
  wire  _any_T_58; // @[CSR.scala 1180:90]
  wire  _any_T_59; // @[CSR.scala 1180:90]
  wire  _any_T_60; // @[CSR.scala 1180:90]
  wire  _any_T_61; // @[CSR.scala 1180:90]
  wire  _any_T_62; // @[CSR.scala 1180:90]
  wire  _any_T_63; // @[CSR.scala 1180:90]
  wire  _any_T_64; // @[CSR.scala 1180:90]
  wire  _any_T_65; // @[CSR.scala 1180:90]
  wire  _any_T_66; // @[CSR.scala 1180:90]
  wire  _any_T_67; // @[CSR.scala 1180:90]
  wire  _any_T_68; // @[CSR.scala 1180:90]
  wire  _any_T_69; // @[CSR.scala 1180:90]
  wire  _any_T_70; // @[CSR.scala 1180:90]
  wire  _any_T_71; // @[CSR.scala 1180:90]
  wire  _any_T_72; // @[CSR.scala 1180:90]
  wire  _any_T_73; // @[CSR.scala 1180:90]
  wire  _any_T_74; // @[CSR.scala 1180:90]
  wire  anyInterrupt; // @[CSR.scala 1180:90]
  wire [2:0] _which_T_38; // @[Mux.scala 47:69]
  wire [3:0] _which_T_39; // @[Mux.scala 47:69]
  wire [3:0] _which_T_40; // @[Mux.scala 47:69]
  wire [3:0] _which_T_41; // @[Mux.scala 47:69]
  wire [3:0] _which_T_42; // @[Mux.scala 47:69]
  wire [3:0] _which_T_43; // @[Mux.scala 47:69]
  wire [3:0] _which_T_44; // @[Mux.scala 47:69]
  wire [3:0] _which_T_45; // @[Mux.scala 47:69]
  wire [3:0] _which_T_46; // @[Mux.scala 47:69]
  wire [3:0] _which_T_47; // @[Mux.scala 47:69]
  wire [3:0] _which_T_48; // @[Mux.scala 47:69]
  wire [3:0] _which_T_49; // @[Mux.scala 47:69]
  wire [3:0] _which_T_50; // @[Mux.scala 47:69]
  wire [3:0] _which_T_51; // @[Mux.scala 47:69]
  wire [3:0] _which_T_52; // @[Mux.scala 47:69]
  wire [3:0] _which_T_53; // @[Mux.scala 47:69]
  wire [3:0] _which_T_54; // @[Mux.scala 47:69]
  wire [3:0] _which_T_55; // @[Mux.scala 47:69]
  wire [3:0] _which_T_56; // @[Mux.scala 47:69]
  wire [3:0] _which_T_57; // @[Mux.scala 47:69]
  wire [3:0] _which_T_58; // @[Mux.scala 47:69]
  wire [3:0] _which_T_59; // @[Mux.scala 47:69]
  wire [3:0] _which_T_60; // @[Mux.scala 47:69]
  wire [3:0] _which_T_61; // @[Mux.scala 47:69]
  wire [3:0] _which_T_62; // @[Mux.scala 47:69]
  wire [3:0] _which_T_64; // @[Mux.scala 47:69]
  wire [3:0] _which_T_65; // @[Mux.scala 47:69]
  wire [3:0] _which_T_66; // @[Mux.scala 47:69]
  wire [3:0] _which_T_67; // @[Mux.scala 47:69]
  wire [3:0] _which_T_68; // @[Mux.scala 47:69]
  wire [3:0] _which_T_69; // @[Mux.scala 47:69]
  wire [3:0] _which_T_70; // @[Mux.scala 47:69]
  wire [3:0] _which_T_71; // @[Mux.scala 47:69]
  wire [3:0] _which_T_72; // @[Mux.scala 47:69]
  wire [3:0] _which_T_73; // @[Mux.scala 47:69]
  wire [3:0] _which_T_74; // @[Mux.scala 47:69]
  wire [3:0] whichInterrupt; // @[Mux.scala 47:69]
  wire [63:0] _GEN_556; // @[CSR.scala 468:67]
  wire  _io_interrupt_T_1; // @[CSR.scala 469:33]
  wire  _io_interrupt_T_2; // @[CSR.scala 469:51]
  wire  _io_interrupt_T_3; // @[CSR.scala 469:88]
  wire  pmp_mask_base_lo; // @[PMP.scala 59:31]
  wire [30:0] pmp_mask_base; // @[Cat.scala 30:58]
  wire [30:0] _pmp_mask_T_1; // @[PMP.scala 60:23]
  wire [30:0] pmp_mask_hi; // @[PMP.scala 60:14]
  wire [32:0] _pmp_mask_T_3; // @[Cat.scala 30:58]
  wire  pmp_mask_base_lo_1; // @[PMP.scala 59:31]
  wire [30:0] pmp_mask_base_1; // @[Cat.scala 30:58]
  wire [30:0] _pmp_mask_T_5; // @[PMP.scala 60:23]
  wire [30:0] pmp_mask_hi_1; // @[PMP.scala 60:14]
  wire [32:0] _pmp_mask_T_7; // @[Cat.scala 30:58]
  wire  pmp_mask_base_lo_2; // @[PMP.scala 59:31]
  wire [30:0] pmp_mask_base_2; // @[Cat.scala 30:58]
  wire [30:0] _pmp_mask_T_9; // @[PMP.scala 60:23]
  wire [30:0] pmp_mask_hi_2; // @[PMP.scala 60:14]
  wire [32:0] _pmp_mask_T_11; // @[Cat.scala 30:58]
  wire  pmp_mask_base_lo_3; // @[PMP.scala 59:31]
  wire [30:0] pmp_mask_base_3; // @[Cat.scala 30:58]
  wire [30:0] _pmp_mask_T_13; // @[PMP.scala 60:23]
  wire [30:0] pmp_mask_hi_3; // @[PMP.scala 60:14]
  wire [32:0] _pmp_mask_T_15; // @[Cat.scala 30:58]
  wire  pmp_mask_base_lo_4; // @[PMP.scala 59:31]
  wire [30:0] pmp_mask_base_4; // @[Cat.scala 30:58]
  wire [30:0] _pmp_mask_T_17; // @[PMP.scala 60:23]
  wire [30:0] pmp_mask_hi_4; // @[PMP.scala 60:14]
  wire [32:0] _pmp_mask_T_19; // @[Cat.scala 30:58]
  wire  pmp_mask_base_lo_5; // @[PMP.scala 59:31]
  wire [30:0] pmp_mask_base_5; // @[Cat.scala 30:58]
  wire [30:0] _pmp_mask_T_21; // @[PMP.scala 60:23]
  wire [30:0] pmp_mask_hi_5; // @[PMP.scala 60:14]
  wire [32:0] _pmp_mask_T_23; // @[Cat.scala 30:58]
  wire  pmp_mask_base_lo_6; // @[PMP.scala 59:31]
  wire [30:0] pmp_mask_base_6; // @[Cat.scala 30:58]
  wire [30:0] _pmp_mask_T_25; // @[PMP.scala 60:23]
  wire [30:0] pmp_mask_hi_6; // @[PMP.scala 60:14]
  wire [32:0] _pmp_mask_T_27; // @[Cat.scala 30:58]
  wire  pmp_mask_base_lo_7; // @[PMP.scala 59:31]
  wire [30:0] pmp_mask_base_7; // @[Cat.scala 30:58]
  wire [30:0] _pmp_mask_T_29; // @[PMP.scala 60:23]
  wire [30:0] pmp_mask_hi_7; // @[PMP.scala 60:14]
  wire [32:0] _pmp_mask_T_31; // @[Cat.scala 30:58]
  reg [63:0] reg_misa; // @[CSR.scala 490:21]
  reg [63:0] _RAND_112;
  wire [6:0] read_mstatus_lo_lo; // @[CSR.scala 491:38]
  wire [18:0] read_mstatus_lo; // @[CSR.scala 491:38]
  wire [16:0] read_mstatus_hi_lo; // @[CSR.scala 491:38]
  wire [102:0] _read_mstatus_T; // @[CSR.scala 491:38]
  wire [63:0] read_mstatus; // @[CSR.scala 491:40]
  wire [7:0] _read_mtvec_T_1; // @[CSR.scala 1209:39]
  wire [31:0] _read_mtvec_T_3; // @[package.scala 165:41]
  wire [31:0] read_mtvec_lo; // @[package.scala 165:35]
  wire [63:0] read_mtvec; // @[Cat.scala 30:58]
  wire [7:0] _read_stvec_T_1; // @[CSR.scala 1209:39]
  wire [38:0] _read_stvec_T_3; // @[package.scala 165:41]
  wire [38:0] read_stvec_lo; // @[package.scala 165:35]
  wire [24:0] read_stvec_hi; // @[Bitwise.scala 72:12]
  wire [63:0] read_stvec; // @[Cat.scala 30:58]
  wire [6:0] lo_2; // @[CSR.scala 497:48]
  wire [63:0] _T_7; // @[CSR.scala 497:48]
  wire [24:0] hi_3; // @[Bitwise.scala 72:12]
  wire [63:0] _T_10; // @[Cat.scala 30:58]
  wire [1:0] _T_14; // @[CSR.scala 1208:36]
  wire [39:0] _GEN_557; // @[CSR.scala 1208:31]
  wire [39:0] _T_15; // @[CSR.scala 1208:31]
  wire [39:0] lo_4; // @[CSR.scala 1208:26]
  wire [23:0] hi_5; // @[Bitwise.scala 72:12]
  wire [63:0] _T_18; // @[Cat.scala 30:58]
  wire [23:0] hi_6; // @[Bitwise.scala 72:12]
  wire [63:0] _T_21; // @[Cat.scala 30:58]
  wire [11:0] lo_5; // @[CSR.scala 512:27]
  wire [31:0] _T_22; // @[CSR.scala 512:27]
  wire [39:0] _T_26; // @[CSR.scala 1208:31]
  wire [39:0] lo_6; // @[CSR.scala 1208:26]
  wire [23:0] hi_8; // @[Bitwise.scala 72:12]
  wire [63:0] _T_29; // @[Cat.scala 30:58]
  wire [7:0] read_fcsr; // @[Cat.scala 30:58]
  wire [63:0] read_sie; // @[CSR.scala 584:28]
  wire [63:0] read_sip; // @[CSR.scala 585:29]
  wire [6:0] lo_lo_4; // @[CSR.scala 599:57]
  wire [18:0] lo_7; // @[CSR.scala 599:57]
  wire [16:0] hi_lo_4; // @[CSR.scala 599:57]
  wire [102:0] _T_30; // @[CSR.scala 599:57]
  wire [23:0] hi_10; // @[Bitwise.scala 72:12]
  wire [63:0] _T_34; // @[Cat.scala 30:58]
  wire [63:0] _T_35; // @[CSR.scala 605:43]
  wire [39:0] _T_39; // @[CSR.scala 1208:31]
  wire [39:0] lo_8; // @[CSR.scala 1208:26]
  wire [23:0] hi_12; // @[Bitwise.scala 72:12]
  wire [63:0] _T_42; // @[Cat.scala 30:58]
  wire [7:0] lo_lo_lo_3; // @[package.scala 36:38]
  wire [7:0] lo_hi_lo_5; // @[package.scala 36:38]
  wire [7:0] hi_lo_lo_4; // @[package.scala 36:38]
  wire [7:0] hi_hi_lo_5; // @[package.scala 36:38]
  wire [15:0] lo_lo_5; // @[Cat.scala 30:58]
  wire [31:0] lo_17; // @[Cat.scala 30:58]
  wire [15:0] hi_lo_5; // @[Cat.scala 30:58]
  wire [63:0] _T_43; // @[Cat.scala 30:58]
  reg [63:0] reg_custom_0; // @[CSR.scala 628:43]
  reg [63:0] _RAND_113;
  wire  _T_46; // @[CSR.scala 636:73]
  wire  _T_47; // @[CSR.scala 636:73]
  wire  _T_49; // @[CSR.scala 636:73]
  wire  _T_50; // @[CSR.scala 636:73]
  wire  _T_51; // @[CSR.scala 636:73]
  wire  _T_52; // @[CSR.scala 636:73]
  wire  _T_53; // @[CSR.scala 636:73]
  wire  _T_54; // @[CSR.scala 636:73]
  wire  _T_55; // @[CSR.scala 636:73]
  wire  _T_56; // @[CSR.scala 636:73]
  wire  _T_57; // @[CSR.scala 636:73]
  wire  _T_58; // @[CSR.scala 636:73]
  wire  _T_59; // @[CSR.scala 636:73]
  wire  _T_60; // @[CSR.scala 636:73]
  wire  _T_61; // @[CSR.scala 636:73]
  wire  _T_62; // @[CSR.scala 636:73]
  wire  _T_63; // @[CSR.scala 636:73]
  wire  _T_64; // @[CSR.scala 636:73]
  wire  _T_65; // @[CSR.scala 636:73]
  wire  _T_66; // @[CSR.scala 636:73]
  wire  _T_67; // @[CSR.scala 636:73]
  wire  _T_155; // @[CSR.scala 636:73]
  wire  _T_156; // @[CSR.scala 636:73]
  wire  _T_157; // @[CSR.scala 636:73]
  wire  _T_158; // @[CSR.scala 636:73]
  wire  _T_159; // @[CSR.scala 636:73]
  wire  _T_160; // @[CSR.scala 636:73]
  wire  _T_161; // @[CSR.scala 636:73]
  wire  _T_162; // @[CSR.scala 636:73]
  wire  _T_163; // @[CSR.scala 636:73]
  wire  _T_164; // @[CSR.scala 636:73]
  wire  _T_165; // @[CSR.scala 636:73]
  wire  _T_166; // @[CSR.scala 636:73]
  wire  _T_167; // @[CSR.scala 636:73]
  wire  _T_168; // @[CSR.scala 636:73]
  wire  _T_169; // @[CSR.scala 636:73]
  wire  _T_170; // @[CSR.scala 636:73]
  wire  _T_172; // @[CSR.scala 636:73]
  wire  _T_173; // @[CSR.scala 636:73]
  wire  _T_174; // @[CSR.scala 636:73]
  wire  _T_175; // @[CSR.scala 636:73]
  wire  _T_176; // @[CSR.scala 636:73]
  wire  _T_177; // @[CSR.scala 636:73]
  wire  _T_178; // @[CSR.scala 636:73]
  wire  _T_179; // @[CSR.scala 636:73]
  wire  _T_188; // @[CSR.scala 636:73]
  wire  _T_189; // @[CSR.scala 636:73]
  wire  _T_191; // @[CSR.scala 636:73]
  wire [63:0] _wdata_T_1; // @[CSR.scala 1186:9]
  wire [63:0] _wdata_T_2; // @[CSR.scala 1186:34]
  wire  _wdata_T_4; // @[CSR.scala 1186:59]
  wire [63:0] _wdata_T_5; // @[CSR.scala 1186:49]
  wire [63:0] wdata; // @[CSR.scala 1186:43]
  wire [31:0] _T_205; // @[Decode.scala 14:65]
  wire  _T_206; // @[Decode.scala 14:121]
  wire [31:0] _T_208; // @[Decode.scala 14:65]
  wire  _T_209; // @[Decode.scala 14:121]
  wire  insn_cease; // @[CSR.scala 652:95]
  wire  insn_wfi; // @[CSR.scala 652:95]
  wire [31:0] _T_220; // @[CSR.scala 659:30]
  wire [31:0] _T_227; // @[Decode.scala 14:65]
  wire  _T_228; // @[Decode.scala 14:121]
  wire [31:0] _T_229; // @[Decode.scala 14:65]
  wire  _T_230; // @[Decode.scala 14:121]
  wire  is_ret; // @[Decode.scala 15:30]
  wire [31:0] _T_236; // @[Decode.scala 14:65]
  wire  is_wfi; // @[Decode.scala 14:121]
  wire [31:0] _T_239; // @[Decode.scala 14:65]
  wire  is_sfence; // @[Decode.scala 14:121]
  wire  _allow_wfi_T; // @[CSR.scala 661:63]
  wire  allow_wfi; // @[CSR.scala 661:71]
  wire  allow_sfence_vma; // @[CSR.scala 662:70]
  wire  allow_sret; // @[CSR.scala 663:72]
  wire [4:0] counter_addr; // @[CSR.scala 664:34]
  wire [31:0] _allow_counter_T_1; // @[CSR.scala 665:68]
  wire  _allow_counter_T_3; // @[CSR.scala 665:50]
  wire  _allow_counter_T_4; // @[CSR.scala 666:44]
  wire [31:0] _allow_counter_T_6; // @[CSR.scala 666:71]
  wire  _allow_counter_T_8; // @[CSR.scala 666:53]
  wire  allow_counter; // @[CSR.scala 665:84]
  wire  _io_decode_0_fp_illegal_T; // @[CSR.scala 667:39]
  wire [11:0] _io_decode_0_fp_csr_T; // @[Decode.scala 14:65]
  wire  _io_decode_0_read_illegal_T_1; // @[CSR.scala 671:44]
  wire  _io_decode_0_read_illegal_T_2; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_3; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_4; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_5; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_6; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_7; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_8; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_9; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_10; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_11; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_12; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_13; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_14; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_15; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_16; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_17; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_18; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_19; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_20; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_21; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_22; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_23; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_24; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_25; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_26; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_27; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_28; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_29; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_30; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_31; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_32; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_33; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_34; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_35; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_36; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_37; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_38; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_39; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_40; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_41; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_42; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_43; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_44; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_45; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_46; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_47; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_48; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_49; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_50; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_51; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_52; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_53; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_54; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_55; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_56; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_57; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_58; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_59; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_60; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_61; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_62; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_63; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_64; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_65; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_66; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_67; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_68; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_69; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_70; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_71; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_72; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_73; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_74; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_75; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_76; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_77; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_78; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_79; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_80; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_81; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_82; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_83; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_84; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_85; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_86; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_87; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_88; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_89; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_90; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_91; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_92; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_93; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_94; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_95; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_96; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_97; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_98; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_99; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_100; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_101; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_102; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_103; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_104; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_105; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_106; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_107; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_108; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_109; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_110; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_111; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_112; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_113; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_114; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_115; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_116; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_117; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_118; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_119; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_120; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_121; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_122; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_123; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_124; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_125; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_126; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_127; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_128; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_129; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_130; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_131; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_132; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_133; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_134; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_135; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_136; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_137; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_138; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_139; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_140; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_141; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_142; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_143; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_144; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_145; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_146; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_147; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_148; // @[CSR.scala 655:99]
  wire  _io_decode_0_read_illegal_T_149; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_150; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_151; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_152; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_153; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_154; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_155; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_156; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_157; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_158; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_159; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_160; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_161; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_162; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_163; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_164; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_165; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_166; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_167; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_168; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_169; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_170; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_171; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_172; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_173; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_174; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_175; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_176; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_177; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_178; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_179; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_180; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_181; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_182; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_183; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_184; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_185; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_186; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_187; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_188; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_189; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_190; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_191; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_192; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_193; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_194; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_195; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_196; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_197; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_198; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_199; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_200; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_201; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_202; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_203; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_204; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_205; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_206; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_207; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_208; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_209; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_210; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_211; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_212; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_213; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_214; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_215; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_216; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_217; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_218; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_219; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_220; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_221; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_222; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_223; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_224; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_225; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_226; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_227; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_228; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_229; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_230; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_231; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_232; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_233; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_234; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_235; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_236; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_237; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_238; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_239; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_240; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_241; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_242; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_243; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_244; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_245; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_246; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_247; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_248; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_249; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_250; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_251; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_252; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_253; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_254; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_255; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_256; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_257; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_258; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_259; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_260; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_261; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_262; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_263; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_264; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_265; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_266; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_267; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_268; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_269; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_270; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_271; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_272; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_273; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_274; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_275; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_276; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_277; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_278; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_279; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_280; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_281; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_282; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_283; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_284; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_285; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_286; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_287; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_288; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_289; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_290; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_291; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_292; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_293; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_294; // @[CSR.scala 655:115]
  wire  _io_decode_0_read_illegal_T_296; // @[CSR.scala 671:62]
  wire  _io_decode_0_read_illegal_T_299; // @[CSR.scala 673:32]
  wire  _io_decode_0_read_illegal_T_300; // @[CSR.scala 672:32]
  wire  _io_decode_0_read_illegal_T_301; // @[package.scala 204:47]
  wire  _io_decode_0_read_illegal_T_302; // @[package.scala 204:60]
  wire  _io_decode_0_read_illegal_T_303; // @[package.scala 204:55]
  wire  _io_decode_0_read_illegal_T_304; // @[package.scala 204:47]
  wire  _io_decode_0_read_illegal_T_305; // @[package.scala 204:60]
  wire  _io_decode_0_read_illegal_T_306; // @[package.scala 204:55]
  wire  _io_decode_0_read_illegal_T_307; // @[CSR.scala 674:66]
  wire  _io_decode_0_read_illegal_T_309; // @[CSR.scala 674:130]
  wire  _io_decode_0_read_illegal_T_310; // @[CSR.scala 673:53]
  wire [11:0] _io_decode_0_read_illegal_T_311; // @[Decode.scala 14:65]
  wire  _io_decode_0_read_illegal_T_312; // @[Decode.scala 14:121]
  wire  _io_decode_0_read_illegal_T_316; // @[CSR.scala 675:42]
  wire  _io_decode_0_read_illegal_T_317; // @[CSR.scala 674:148]
  wire  _io_decode_0_read_illegal_T_320; // @[CSR.scala 677:21]
  wire  _io_decode_0_write_flush_T; // @[CSR.scala 679:40]
  wire  _io_decode_0_write_flush_T_1; // @[CSR.scala 679:71]
  wire  _io_decode_0_write_flush_T_2; // @[CSR.scala 679:57]
  wire  _io_decode_0_write_flush_T_3; // @[CSR.scala 679:99]
  wire  _io_decode_0_write_flush_T_4; // @[CSR.scala 679:130]
  wire  _io_decode_0_write_flush_T_5; // @[CSR.scala 679:116]
  wire  _io_decode_0_write_flush_T_6; // @[CSR.scala 679:85]
  wire  _io_decode_0_system_illegal_T_3; // @[CSR.scala 681:14]
  wire  _io_decode_0_system_illegal_T_4; // @[CSR.scala 680:64]
  wire  _io_decode_0_system_illegal_T_6; // @[CSR.scala 682:14]
  wire  _io_decode_0_system_illegal_T_7; // @[CSR.scala 681:28]
  wire  _io_decode_0_system_illegal_T_9; // @[CSR.scala 683:14]
  wire  _io_decode_0_system_illegal_T_11; // @[CSR.scala 683:32]
  wire  _io_decode_0_system_illegal_T_13; // @[CSR.scala 683:49]
  wire  _io_decode_0_system_illegal_T_14; // @[CSR.scala 682:29]
  wire  _io_decode_0_system_illegal_T_16; // @[CSR.scala 684:17]
  wire [11:0] _debugTVec_T; // @[CSR.scala 697:37]
  wire [11:0] debugTVec; // @[CSR.scala 697:22]
  wire [63:0] notDebugTVec_base; // @[CSR.scala 705:19]
  wire [7:0] notDebugTVec_interruptVec_lo; // @[CSR.scala 706:59]
  wire [55:0] notDebugTVec_interruptVec_hi; // @[CSR.scala 707:33]
  wire [63:0] notDebugTVec_interruptVec; // @[Cat.scala 30:58]
  wire  _notDebugTVec_doVector_T_2; // @[CSR.scala 708:28]
  wire  _notDebugTVec_doVector_T_4; // @[CSR.scala 708:94]
  wire  notDebugTVec_doVector; // @[CSR.scala 708:55]
  wire [63:0] _notDebugTVec_T_1; // @[CSR.scala 709:56]
  wire [63:0] notDebugTVec; // @[CSR.scala 709:8]
  wire [63:0] tvec; // @[CSR.scala 723:17]
  wire  _io_status_sd_T; // @[CSR.scala 729:32]
  wire  _io_status_sd_T_1; // @[CSR.scala 729:53]
  wire  _io_status_sd_T_2; // @[CSR.scala 729:37]
  wire  _io_status_sd_T_3; // @[CSR.scala 729:74]
  wire  _io_status_dprv_x87_T_1; // @[CSR.scala 734:53]
  reg [1:0] io_status_dprv_REG; // @[CSR.scala 734:24]
  reg [31:0] _RAND_114;
  wire [1:0] _T_244; // @[Bitwise.scala 47:55]
  wire [1:0] _T_246; // @[Bitwise.scala 47:55]
  wire [2:0] _T_248; // @[Bitwise.scala 47:55]
  wire  _T_250; // @[CSR.scala 739:79]
  wire  _T_252; // @[CSR.scala 739:9]
  wire  _T_255; // @[CSR.scala 741:18]
  wire  _T_257; // @[CSR.scala 741:36]
  wire  _GEN_48; // @[CSR.scala 741:51]
  wire  _T_258; // @[CSR.scala 742:28]
  wire  _T_259; // @[CSR.scala 742:32]
  wire  _T_260; // @[CSR.scala 742:55]
  wire  _T_262; // @[CSR.scala 745:22]
  wire  _GEN_50; // @[CSR.scala 745:36]
  wire  _T_272; // @[CSR.scala 748:29]
  wire  _T_274; // @[CSR.scala 748:9]
  wire [39:0] _epc_T_1; // @[CSR.scala 1207:31]
  wire [39:0] epc; // @[CSR.scala 1207:26]
  wire [1:0] _reg_dcsr_cause_T; // @[CSR.scala 759:86]
  wire [1:0] _reg_dcsr_cause_T_1; // @[CSR.scala 759:56]
  wire  _GEN_52; // @[CSR.scala 756:25]
  wire [39:0] _GEN_53; // @[CSR.scala 756:25]
  wire [39:0] _GEN_63; // @[CSR.scala 772:35]
  wire  _GEN_67; // @[CSR.scala 772:35]
  wire [1:0] _GEN_68; // @[CSR.scala 772:35]
  wire [39:0] _GEN_71; // @[CSR.scala 772:35]
  wire  _GEN_74; // @[CSR.scala 772:35]
  wire [1:0] _GEN_75; // @[CSR.scala 772:35]
  wire  _GEN_76; // @[CSR.scala 772:35]
  wire [39:0] _GEN_97; // @[CSR.scala 755:24]
  wire [39:0] _GEN_106; // @[CSR.scala 755:24]
  wire  _GEN_110; // @[CSR.scala 755:24]
  wire [1:0] _GEN_111; // @[CSR.scala 755:24]
  wire [39:0] _GEN_113; // @[CSR.scala 755:24]
  wire  _GEN_116; // @[CSR.scala 755:24]
  wire [1:0] _GEN_117; // @[CSR.scala 755:24]
  wire  _GEN_118; // @[CSR.scala 755:24]
  wire [39:0] _GEN_120; // @[CSR.scala 754:20]
  wire [39:0] _GEN_129; // @[CSR.scala 754:20]
  wire  _GEN_133; // @[CSR.scala 754:20]
  wire [1:0] _GEN_134; // @[CSR.scala 754:20]
  wire [39:0] _GEN_136; // @[CSR.scala 754:20]
  wire  _GEN_139; // @[CSR.scala 754:20]
  wire [1:0] _GEN_140; // @[CSR.scala 754:20]
  wire  _GEN_141; // @[CSR.scala 754:20]
  wire [39:0] _GEN_151; // @[CSR.scala 821:70]
  wire  _GEN_158; // @[CSR.scala 815:52]
  wire [1:0] _GEN_159; // @[CSR.scala 815:52]
  wire [39:0] _GEN_161; // @[CSR.scala 815:52]
  wire  _T_412; // @[CSR.scala 839:32]
  wire [1:0] _GEN_171; // @[CSR.scala 813:19]
  wire [63:0] _GEN_172; // @[CSR.scala 813:19]
  reg  io_status_cease_r; // @[Reg.scala 27:20]
  reg [31:0] _RAND_115;
  wire  _GEN_181; // @[Reg.scala 28:19]
  wire [63:0] _io_rw_rdata_T_1; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_2; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_4; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_5; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_6; // @[Mux.scala 27:72]
  wire [15:0] _io_rw_rdata_T_7; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_8; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_9; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_10; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_11; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_12; // @[Mux.scala 27:72]
  wire  _io_rw_rdata_T_13; // @[Mux.scala 27:72]
  wire [31:0] _io_rw_rdata_T_14; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_15; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_16; // @[Mux.scala 27:72]
  wire [4:0] _io_rw_rdata_T_17; // @[Mux.scala 27:72]
  wire [2:0] _io_rw_rdata_T_18; // @[Mux.scala 27:72]
  wire [7:0] _io_rw_rdata_T_19; // @[Mux.scala 27:72]
  wire [2:0] _io_rw_rdata_T_20; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_21; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_22; // @[Mux.scala 27:72]
  wire [31:0] _io_rw_rdata_T_110; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_111; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_112; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_113; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_114; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_115; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_116; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_117; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_118; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_119; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_120; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_121; // @[Mux.scala 27:72]
  wire [31:0] _io_rw_rdata_T_122; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_123; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_124; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_125; // @[Mux.scala 27:72]
  wire [29:0] _io_rw_rdata_T_127; // @[Mux.scala 27:72]
  wire [29:0] _io_rw_rdata_T_128; // @[Mux.scala 27:72]
  wire [29:0] _io_rw_rdata_T_129; // @[Mux.scala 27:72]
  wire [29:0] _io_rw_rdata_T_130; // @[Mux.scala 27:72]
  wire [29:0] _io_rw_rdata_T_131; // @[Mux.scala 27:72]
  wire [29:0] _io_rw_rdata_T_132; // @[Mux.scala 27:72]
  wire [29:0] _io_rw_rdata_T_133; // @[Mux.scala 27:72]
  wire [29:0] _io_rw_rdata_T_134; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_143; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_144; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_146; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_148; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_150; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_151; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_152; // @[Mux.scala 27:72]
  wire [63:0] _GEN_565; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_153; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_154; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_155; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_156; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_157; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_158; // @[Mux.scala 27:72]
  wire [63:0] _GEN_566; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_159; // @[Mux.scala 27:72]
  wire [63:0] _GEN_567; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_160; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_161; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_162; // @[Mux.scala 27:72]
  wire [63:0] _GEN_568; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_163; // @[Mux.scala 27:72]
  wire [63:0] _GEN_569; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_164; // @[Mux.scala 27:72]
  wire [63:0] _GEN_570; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_165; // @[Mux.scala 27:72]
  wire [63:0] _GEN_571; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_166; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_167; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_168; // @[Mux.scala 27:72]
  wire [63:0] _GEN_572; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_256; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_257; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_258; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_259; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_260; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_261; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_262; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_263; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_264; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_265; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_266; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_267; // @[Mux.scala 27:72]
  wire [63:0] _GEN_573; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_268; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_269; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_270; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_271; // @[Mux.scala 27:72]
  wire [63:0] _GEN_574; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_273; // @[Mux.scala 27:72]
  wire [63:0] _GEN_575; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_274; // @[Mux.scala 27:72]
  wire [63:0] _GEN_576; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_275; // @[Mux.scala 27:72]
  wire [63:0] _GEN_577; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_276; // @[Mux.scala 27:72]
  wire [63:0] _GEN_578; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_277; // @[Mux.scala 27:72]
  wire [63:0] _GEN_579; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_278; // @[Mux.scala 27:72]
  wire [63:0] _GEN_580; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_279; // @[Mux.scala 27:72]
  wire [63:0] _GEN_581; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_280; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_289; // @[Mux.scala 27:72]
  wire [63:0] _io_rw_rdata_T_290; // @[Mux.scala 27:72]
  wire  _T_416; // @[package.scala 15:47]
  wire  _T_417; // @[package.scala 15:47]
  wire  _T_418; // @[package.scala 15:47]
  wire [4:0] _lo_T; // @[CSR.scala 887:30]
  wire [4:0] _GEN_182; // @[CSR.scala 886:30]
  wire  _csr_wen_T_3; // @[package.scala 72:59]
  wire  csr_wen; // @[package.scala 72:59]
  wire [102:0] _new_mstatus_WIRE;
  wire  new_mstatus_sie; // @[CSR.scala 902:47]
  wire  new_mstatus_mie; // @[CSR.scala 902:47]
  wire  new_mstatus_spie; // @[CSR.scala 902:47]
  wire  new_mstatus_mpie; // @[CSR.scala 902:47]
  wire  new_mstatus_spp; // @[CSR.scala 902:47]
  wire [1:0] new_mstatus_mpp; // @[CSR.scala 902:47]
  wire [1:0] new_mstatus_fs; // @[CSR.scala 902:47]
  wire  new_mstatus_mprv; // @[CSR.scala 902:47]
  wire  new_mstatus_sum; // @[CSR.scala 902:47]
  wire  new_mstatus_mxr; // @[CSR.scala 902:47]
  wire  new_mstatus_tvm; // @[CSR.scala 902:47]
  wire  new_mstatus_tw; // @[CSR.scala 902:47]
  wire  new_mstatus_tsr; // @[CSR.scala 902:47]
  wire  _reg_mstatus_mpp_T_2; // @[CSR.scala 1190:35]
  wire  _reg_mstatus_fs_T; // @[CSR.scala 1211:73]
  wire [1:0] _GEN_188; // @[CSR.scala 901:39]
  wire  f; // @[CSR.scala 928:20]
  wire  _T_1834; // @[CSR.scala 930:43]
  wire [3:0] _reg_misa_T_2; // @[CSR.scala 932:38]
  wire [63:0] _GEN_582; // @[CSR.scala 932:32]
  wire [63:0] _reg_misa_T_3; // @[CSR.scala 932:32]
  wire [63:0] _reg_misa_T_5; // @[CSR.scala 932:55]
  wire [63:0] _reg_misa_T_7; // @[CSR.scala 932:73]
  wire [63:0] _reg_misa_T_8; // @[CSR.scala 932:62]
  wire [15:0] _new_mip_T; // @[CSR.scala 940:59]
  wire [15:0] _new_mip_T_2; // @[CSR.scala 1186:9]
  wire [63:0] _GEN_583; // @[CSR.scala 1186:34]
  wire [63:0] _new_mip_T_3; // @[CSR.scala 1186:34]
  wire [63:0] _new_mip_T_8; // @[CSR.scala 1186:43]
  wire  new_mip_ssip; // @[CSR.scala 940:88]
  wire  new_mip_stip; // @[CSR.scala 940:88]
  wire  new_mip_seip; // @[CSR.scala 940:88]
  wire [63:0] _reg_mie_T; // @[CSR.scala 947:59]
  wire [63:0] _reg_mepc_T_1; // @[CSR.scala 1207:31]
  wire [63:0] _GEN_204; // @[CSR.scala 948:40]
  wire [63:0] _GEN_206; // @[CSR.scala 951:40]
  wire [63:0] _reg_mcause_T; // @[CSR.scala 952:62]
  wire [63:0] _reg_mcountinhibit_T_1; // @[CSR.scala 968:76]
  wire [63:0] _GEN_209; // @[CSR.scala 968:47]
  wire [63:0] _GEN_210; // @[CSR.scala 1204:31]
  wire [63:0] _GEN_212; // @[CSR.scala 1204:31]
  wire [63:0] _GEN_215; // @[CSR.scala 974:40]
  wire [63:0] _GEN_217; // @[CSR.scala 975:40]
  wire [63:0] _GEN_219; // @[CSR.scala 976:38]
  wire [63:0] _GEN_220; // @[CSR.scala 976:38]
  wire [1:0] new_dcsr_prv; // @[CSR.scala 984:43]
  wire  new_dcsr_step; // @[CSR.scala 984:43]
  wire  new_dcsr_ebreaku; // @[CSR.scala 984:43]
  wire  new_dcsr_ebreaks; // @[CSR.scala 984:43]
  wire  new_dcsr_ebreakm; // @[CSR.scala 984:43]
  wire  _reg_dcsr_prv_T; // @[CSR.scala 1190:35]
  wire [63:0] _GEN_226; // @[CSR.scala 991:42]
  wire [1:0] _GEN_230; // @[CSR.scala 998:41]
  wire [63:0] _new_sip_T_1; // @[CSR.scala 1011:52]
  wire [63:0] _new_sip_T_2; // @[CSR.scala 1011:78]
  wire [63:0] _new_sip_T_3; // @[CSR.scala 1011:69]
  wire  new_sip_ssip; // @[CSR.scala 1011:41]
  wire [43:0] new_satp_ppn; // @[CSR.scala 1016:45]
  wire [3:0] new_satp_mode; // @[CSR.scala 1016:45]
  wire  _T_1837; // @[package.scala 15:47]
  wire  _T_1838; // @[package.scala 15:47]
  wire  _T_1839; // @[package.scala 72:59]
  wire [3:0] _reg_satp_mode_T; // @[CSR.scala 1019:44]
  wire [63:0] _reg_mie_T_2; // @[CSR.scala 1025:64]
  wire [63:0] _reg_mie_T_4; // @[CSR.scala 1025:81]
  wire [63:0] _GEN_242; // @[CSR.scala 1027:42]
  wire [63:0] _GEN_243; // @[CSR.scala 1028:42]
  wire [63:0] _reg_scause_T; // @[CSR.scala 1029:64]
  wire [63:0] _GEN_248; // @[CSR.scala 1033:44]
  wire [63:0] _GEN_249; // @[CSR.scala 1036:44]
  wire  _T_1842; // @[CSR.scala 1042:55]
  wire [63:0] _GEN_251; // @[CSR.scala 1043:44]
  wire [63:0] _newBPC_T_2; // @[CSR.scala 1186:9]
  wire [63:0] _newBPC_T_3; // @[CSR.scala 1186:34]
  wire [63:0] _newBPC_T_8; // @[CSR.scala 1186:43]
  wire  newBPC_action; // @[CSR.scala 1061:96]
  wire  newBPC_dmode; // @[CSR.scala 1061:96]
  wire  dMode; // @[CSR.scala 1062:38]
  wire  _GEN_252; // @[CSR.scala 1064:51]
  wire [63:0] _GEN_268; // @[CSR.scala 1042:70]
  wire  _T_1853; // @[CSR.scala 1074:57]
  wire  newCfg_r; // @[CSR.scala 1075:46]
  wire  newCfg_w; // @[CSR.scala 1075:46]
  wire  newCfg_x; // @[CSR.scala 1075:46]
  wire [1:0] newCfg_a; // @[CSR.scala 1075:46]
  wire  newCfg_l; // @[CSR.scala 1075:46]
  wire  _reg_pmp_0_cfg_w_T; // @[CSR.scala 1078:31]
  wire  _T_1857; // @[PMP.scala 49:20]
  wire  _T_1858; // @[PMP.scala 51:62]
  wire  _T_1859; // @[PMP.scala 51:44]
  wire  _T_1861; // @[CSR.scala 1083:45]
  wire [63:0] _GEN_323; // @[CSR.scala 1083:71]
  wire  _T_1863; // @[CSR.scala 1074:57]
  wire  newCfg_1_r; // @[CSR.scala 1075:46]
  wire  newCfg_1_w; // @[CSR.scala 1075:46]
  wire  newCfg_1_x; // @[CSR.scala 1075:46]
  wire [1:0] newCfg_1_a; // @[CSR.scala 1075:46]
  wire  newCfg_1_l; // @[CSR.scala 1075:46]
  wire  _reg_pmp_1_cfg_w_T; // @[CSR.scala 1078:31]
  wire  _T_1867; // @[PMP.scala 49:20]
  wire  _T_1868; // @[PMP.scala 51:62]
  wire  _T_1869; // @[PMP.scala 51:44]
  wire  _T_1871; // @[CSR.scala 1083:45]
  wire [63:0] _GEN_330; // @[CSR.scala 1083:71]
  wire  _T_1873; // @[CSR.scala 1074:57]
  wire  newCfg_2_r; // @[CSR.scala 1075:46]
  wire  newCfg_2_w; // @[CSR.scala 1075:46]
  wire  newCfg_2_x; // @[CSR.scala 1075:46]
  wire [1:0] newCfg_2_a; // @[CSR.scala 1075:46]
  wire  newCfg_2_l; // @[CSR.scala 1075:46]
  wire  _reg_pmp_2_cfg_w_T; // @[CSR.scala 1078:31]
  wire  _T_1877; // @[PMP.scala 49:20]
  wire  _T_1878; // @[PMP.scala 51:62]
  wire  _T_1879; // @[PMP.scala 51:44]
  wire  _T_1881; // @[CSR.scala 1083:45]
  wire [63:0] _GEN_337; // @[CSR.scala 1083:71]
  wire  _T_1883; // @[CSR.scala 1074:57]
  wire  newCfg_3_r; // @[CSR.scala 1075:46]
  wire  newCfg_3_w; // @[CSR.scala 1075:46]
  wire  newCfg_3_x; // @[CSR.scala 1075:46]
  wire [1:0] newCfg_3_a; // @[CSR.scala 1075:46]
  wire  newCfg_3_l; // @[CSR.scala 1075:46]
  wire  _reg_pmp_3_cfg_w_T; // @[CSR.scala 1078:31]
  wire  _T_1887; // @[PMP.scala 49:20]
  wire  _T_1888; // @[PMP.scala 51:62]
  wire  _T_1889; // @[PMP.scala 51:44]
  wire  _T_1891; // @[CSR.scala 1083:45]
  wire [63:0] _GEN_344; // @[CSR.scala 1083:71]
  wire  _T_1893; // @[CSR.scala 1074:57]
  wire  newCfg_4_r; // @[CSR.scala 1075:46]
  wire  newCfg_4_w; // @[CSR.scala 1075:46]
  wire  newCfg_4_x; // @[CSR.scala 1075:46]
  wire [1:0] newCfg_4_a; // @[CSR.scala 1075:46]
  wire  newCfg_4_l; // @[CSR.scala 1075:46]
  wire  _reg_pmp_4_cfg_w_T; // @[CSR.scala 1078:31]
  wire  _T_1897; // @[PMP.scala 49:20]
  wire  _T_1898; // @[PMP.scala 51:62]
  wire  _T_1899; // @[PMP.scala 51:44]
  wire  _T_1901; // @[CSR.scala 1083:45]
  wire [63:0] _GEN_351; // @[CSR.scala 1083:71]
  wire  _T_1903; // @[CSR.scala 1074:57]
  wire  newCfg_5_r; // @[CSR.scala 1075:46]
  wire  newCfg_5_w; // @[CSR.scala 1075:46]
  wire  newCfg_5_x; // @[CSR.scala 1075:46]
  wire [1:0] newCfg_5_a; // @[CSR.scala 1075:46]
  wire  newCfg_5_l; // @[CSR.scala 1075:46]
  wire  _reg_pmp_5_cfg_w_T; // @[CSR.scala 1078:31]
  wire  _T_1907; // @[PMP.scala 49:20]
  wire  _T_1908; // @[PMP.scala 51:62]
  wire  _T_1909; // @[PMP.scala 51:44]
  wire  _T_1911; // @[CSR.scala 1083:45]
  wire [63:0] _GEN_358; // @[CSR.scala 1083:71]
  wire  _T_1913; // @[CSR.scala 1074:57]
  wire  newCfg_6_r; // @[CSR.scala 1075:46]
  wire  newCfg_6_w; // @[CSR.scala 1075:46]
  wire  newCfg_6_x; // @[CSR.scala 1075:46]
  wire [1:0] newCfg_6_a; // @[CSR.scala 1075:46]
  wire  newCfg_6_l; // @[CSR.scala 1075:46]
  wire  _reg_pmp_6_cfg_w_T; // @[CSR.scala 1078:31]
  wire  _T_1917; // @[PMP.scala 49:20]
  wire  _T_1918; // @[PMP.scala 51:62]
  wire  _T_1919; // @[PMP.scala 51:44]
  wire  _T_1921; // @[CSR.scala 1083:45]
  wire [63:0] _GEN_365; // @[CSR.scala 1083:71]
  wire  _T_1923; // @[CSR.scala 1074:57]
  wire  newCfg_7_r; // @[CSR.scala 1075:46]
  wire  newCfg_7_w; // @[CSR.scala 1075:46]
  wire  newCfg_7_x; // @[CSR.scala 1075:46]
  wire [1:0] newCfg_7_a; // @[CSR.scala 1075:46]
  wire  newCfg_7_l; // @[CSR.scala 1075:46]
  wire  _reg_pmp_7_cfg_w_T; // @[CSR.scala 1078:31]
  wire  _T_1929; // @[PMP.scala 51:44]
  wire  _T_1931; // @[CSR.scala 1083:45]
  wire [63:0] _GEN_372; // @[CSR.scala 1083:71]
  wire [63:0] _reg_custom_0_T; // @[CSR.scala 1090:23]
  wire [63:0] _reg_custom_0_T_2; // @[CSR.scala 1090:38]
  wire [63:0] _reg_custom_0_T_3; // @[CSR.scala 1090:31]
  wire [1:0] _GEN_385; // @[CSR.scala 900:18]
  wire [63:0] _GEN_400; // @[CSR.scala 900:18]
  wire [63:0] _GEN_402; // @[CSR.scala 900:18]
  wire [63:0] _GEN_405; // @[CSR.scala 900:18]
  wire [63:0] _GEN_406; // @[CSR.scala 900:18]
  wire [63:0] _GEN_408; // @[CSR.scala 900:18]
  wire [63:0] _GEN_411; // @[CSR.scala 900:18]
  wire [63:0] _GEN_412; // @[CSR.scala 900:18]
  wire [63:0] _GEN_418; // @[CSR.scala 900:18]
  wire [63:0] _GEN_423; // @[CSR.scala 900:18]
  wire [63:0] _GEN_424; // @[CSR.scala 900:18]
  wire [63:0] _GEN_429; // @[CSR.scala 900:18]
  wire [63:0] _GEN_430; // @[CSR.scala 900:18]
  wire [63:0] _GEN_432; // @[CSR.scala 900:18]
  wire [63:0] _GEN_470; // @[CSR.scala 900:18]
  wire [63:0] _GEN_477; // @[CSR.scala 900:18]
  wire [63:0] _GEN_484; // @[CSR.scala 900:18]
  wire [63:0] _GEN_491; // @[CSR.scala 900:18]
  wire [63:0] _GEN_498; // @[CSR.scala 900:18]
  wire [63:0] _GEN_505; // @[CSR.scala 900:18]
  wire [63:0] _GEN_512; // @[CSR.scala 900:18]
  wire [63:0] _GEN_519; // @[CSR.scala 900:18]
  wire  _io_trace_0_valid_T; // @[CSR.scala 1165:26]
  reg [19:0] CSRFile_state; // @[Register tracking CSRFile state]
  reg [31:0] _RAND_116;
  reg  CSRFile_cov [0:1048575]; // @[Coverage map for CSRFile]
  reg [31:0] _RAND_117;
  wire  CSRFile_cov_read_data; // @[Coverage map for CSRFile]
  wire [19:0] CSRFile_cov_read_addr; // @[Coverage map for CSRFile]
  wire  CSRFile_cov_write_data; // @[Coverage map for CSRFile]
  wire [19:0] CSRFile_cov_write_addr; // @[Coverage map for CSRFile]
  wire  CSRFile_cov_write_mask; // @[Coverage map for CSRFile]
  wire  CSRFile_cov_write_en; // @[Coverage map for CSRFile]
  reg [29:0] CSRFile_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_118;
  wire [19:0] reg_pmp_5_cfg_l_shl;
  wire [19:0] reg_pmp_5_cfg_l_pad;
  wire [1:0] reg_debug_shl;
  wire [19:0] reg_debug_pad;
  wire [16:0] reg_mstatus_sie_shl;
  wire [19:0] reg_mstatus_sie_pad;
  wire [14:0] reg_dcsr_prv_shl;
  wire [19:0] reg_dcsr_prv_pad;
  wire [17:0] reg_mcountinhibit_shl;
  wire [19:0] reg_mcountinhibit_pad;
  wire [2:0] reg_unmie_shl;
  wire [19:0] reg_unmie_pad;
  wire [14:0] reg_pmp_7_cfg_a_shl;
  wire [19:0] reg_pmp_7_cfg_a_pad;
  wire [1:0] reg_mstatus_mpp_shl;
  wire [19:0] reg_mstatus_mpp_pad;
  wire [6:0] reg_pmp_2_cfg_l_shl;
  wire [19:0] reg_pmp_2_cfg_l_pad;
  wire [18:0] reg_pmp_1_cfg_l_shl;
  wire [19:0] reg_pmp_1_cfg_l_pad;
  wire [9:0] reg_mip_seip_shl;
  wire [19:0] reg_mip_seip_pad;
  wire [1:0] reg_rnmie_shl;
  wire [19:0] reg_rnmie_pad;
  wire [10:0] reg_mip_ssip_shl;
  wire [19:0] reg_mip_ssip_pad;
  wire [2:0] reg_bp_0_control_dmode_shl;
  wire [19:0] reg_bp_0_control_dmode_pad;
  wire [11:0] reg_pmp_4_cfg_l_shl;
  wire [19:0] reg_pmp_4_cfg_l_pad;
  wire [1:0] reg_dcsr_ebreaks_shl;
  wire [19:0] reg_dcsr_ebreaks_pad;
  wire [13:0] reg_pmp_6_cfg_l_shl;
  wire [19:0] reg_pmp_6_cfg_l_pad;
  wire [3:0] reg_mstatus_prv_shl;
  wire [19:0] reg_mstatus_prv_pad;
  wire [8:0] reg_dcsr_ebreakm_shl;
  wire [19:0] reg_dcsr_ebreakm_pad;
  wire  reg_pmp_7_cfg_l_shl;
  wire [19:0] reg_pmp_7_cfg_l_pad;
  wire [18:0] reg_pmp_0_cfg_l_shl;
  wire [19:0] reg_pmp_0_cfg_l_pad;
  wire [1:0] reg_pmp_3_cfg_l_shl;
  wire [19:0] reg_pmp_3_cfg_l_pad;
  wire [13:0] reg_mstatus_spp_shl;
  wire [19:0] reg_mstatus_spp_pad;
  wire [12:0] reg_mip_stip_shl;
  wire [19:0] reg_mip_stip_pad;
  wire [13:0] reg_dcsr_ebreaku_shl;
  wire [19:0] reg_dcsr_ebreaku_pad;
  wire  reg_mstatus_mprv_shl;
  wire [19:0] reg_mstatus_mprv_pad;
  wire [13:0] reg_singleStepped_shl;
  wire [19:0] reg_singleStepped_pad;
  wire [11:0] reg_mstatus_mie_shl;
  wire [19:0] reg_mstatus_mie_pad;
  wire [19:0] CSRFile_xor16;
  wire [19:0] CSRFile_xor7;
  wire [19:0] CSRFile_xor17;
  wire [19:0] CSRFile_xor18;
  wire [19:0] CSRFile_xor8;
  wire [19:0] CSRFile_xor3;
  wire [19:0] CSRFile_xor20;
  wire [19:0] CSRFile_xor9;
  wire [19:0] CSRFile_xor21;
  wire [19:0] CSRFile_xor22;
  wire [19:0] CSRFile_xor10;
  wire [19:0] CSRFile_xor4;
  wire [19:0] CSRFile_xor1;
  wire [19:0] CSRFile_xor24;
  wire [19:0] CSRFile_xor11;
  wire [19:0] CSRFile_xor25;
  wire [19:0] CSRFile_xor26;
  wire [19:0] CSRFile_xor12;
  wire [19:0] CSRFile_xor5;
  wire [19:0] CSRFile_xor28;
  wire [19:0] CSRFile_xor13;
  wire [19:0] CSRFile_xor29;
  wire [19:0] CSRFile_xor30;
  wire [19:0] CSRFile_xor14;
  wire [19:0] CSRFile_xor6;
  wire [19:0] CSRFile_xor2;
  wire [19:0] CSRFile_xor0;
  wire  stopEn0;
  wire  stopEn1;
  wire  CSRFile_or0;
  reg  CSRFile_metaAssert;
  reg [31:0] _RAND_119;
  assign system_insn = io_rw_cmd == 3'h4; // @[CSR.scala 639:31]
  assign _T_192 = {io_rw_addr, 20'h0}; // @[CSR.scala 652:28]
  assign _T_199 = _T_192 & 32'h12400000; // @[Decode.scala 14:65]
  assign _T_200 = _T_199 == 32'h10000000; // @[Decode.scala 14:121]
  assign _T_201 = _T_192 & 32'h40000000; // @[Decode.scala 14:65]
  assign _T_202 = _T_201 == 32'h40000000; // @[Decode.scala 14:121]
  assign _T_204 = _T_200 | _T_202; // @[Decode.scala 15:30]
  assign insn_ret = system_insn & _T_204; // @[CSR.scala 652:95]
  assign _T_406 = io_rw_addr[10] & io_rw_addr[7]; // @[CSR.scala 821:52]
  assign _GEN_149 = _T_406 ? reg_dcsr_prv : reg_mstatus_mpp; // @[CSR.scala 821:70]
  assign ret_prv = io_rw_addr[9] ? _GEN_149 : {{1'd0}, reg_mstatus_spp}; // @[CSR.scala 815:52]
  assign _T_193 = _T_192 & 32'h10100000; // @[Decode.scala 14:65]
  assign _T_194 = _T_193 == 32'h0; // @[Decode.scala 14:121]
  assign insn_call = system_insn & _T_194; // @[CSR.scala 652:95]
  assign _T_197 = _T_193 == 32'h100000; // @[Decode.scala 14:121]
  assign insn_break = system_insn & _T_197; // @[CSR.scala 652:95]
  assign _exception_T = insn_call | insn_break; // @[CSR.scala 738:29]
  assign exception = _exception_T | io_exception; // @[CSR.scala 738:43]
  assign _GEN_20 = {{2'd0}, reg_mstatus_prv}; // @[CSR.scala 688:36]
  assign _cause_T_1 = _GEN_20 + 4'h8; // @[CSR.scala 688:36]
  assign _cause_T_2 = insn_break ? 64'h3 : io_cause; // @[CSR.scala 689:14]
  assign cause = insn_call ? {{60'd0}, _cause_T_1} : _cause_T_2; // @[CSR.scala 688:8]
  assign cause_lsbs = cause[7:0]; // @[CSR.scala 690:25]
  assign _causeIsDebugInt_T_1 = cause_lsbs == 8'he; // @[CSR.scala 691:53]
  assign causeIsDebugInt = cause[63] & _causeIsDebugInt_T_1; // @[CSR.scala 691:39]
  assign _trapToDebug_T = reg_singleStepped | causeIsDebugInt; // @[CSR.scala 694:60]
  assign causeIsDebugTrigger = ~cause[63] & _causeIsDebugInt_T_1; // @[CSR.scala 692:44]
  assign _trapToDebug_T_1 = _trapToDebug_T | causeIsDebugTrigger; // @[CSR.scala 694:79]
  assign _causeIsDebugBreak_T_2 = ~cause[63] & insn_break; // @[CSR.scala 693:42]
  assign _causeIsDebugBreak_T_3 = {reg_dcsr_ebreakm,1'h0,reg_dcsr_ebreaks,reg_dcsr_ebreaku}; // @[Cat.scala 30:58]
  assign _causeIsDebugBreak_T_4 = _causeIsDebugBreak_T_3 >> reg_mstatus_prv; // @[CSR.scala 693:134]
  assign causeIsDebugBreak = _causeIsDebugBreak_T_2 & _causeIsDebugBreak_T_4[0]; // @[CSR.scala 693:56]
  assign _trapToDebug_T_2 = _trapToDebug_T_1 | causeIsDebugBreak; // @[CSR.scala 694:102]
  assign trapToDebug = _trapToDebug_T_2 | reg_debug; // @[CSR.scala 694:123]
  assign _GEN_56 = reg_debug ? reg_mstatus_prv : 2'h3; // @[CSR.scala 756:25]
  assign _delegate_T = reg_mstatus_prv <= 2'h1; // @[CSR.scala 698:59]
  assign read_mideleg = reg_mideleg & 64'h222; // @[CSR.scala 384:36]
  assign _delegate_T_3 = read_mideleg >> cause_lsbs; // @[CSR.scala 698:102]
  assign read_medeleg = reg_medeleg & 64'hb15d; // @[CSR.scala 388:36]
  assign _delegate_T_5 = read_medeleg >> cause_lsbs; // @[CSR.scala 698:128]
  assign _delegate_T_7 = cause[63] ? _delegate_T_3[0] : _delegate_T_5[0]; // @[CSR.scala 698:74]
  assign delegate = _delegate_T & _delegate_T_7; // @[CSR.scala 698:68]
  assign nmie = reg_rnmie & reg_unmie; // @[CSR.scala 409:24]
  assign _T_279 = delegate & nmie; // @[CSR.scala 772:26]
  assign _GEN_70 = _T_279 ? 2'h1 : 2'h3; // @[CSR.scala 772:35]
  assign _GEN_100 = trapToDebug ? _GEN_56 : _GEN_70; // @[CSR.scala 755:24]
  assign _GEN_123 = exception ? _GEN_100 : reg_mstatus_prv; // @[CSR.scala 754:20]
  assign new_prv = insn_ret ? ret_prv : _GEN_123; // @[CSR.scala 813:19]
  assign _reg_mstatus_prv_T = new_prv == 2'h2; // @[CSR.scala 1190:35]
  assign read_mcounteren = reg_mcounteren & 32'h7; // @[CSR.scala 414:30]
  assign read_scounteren = reg_scounteren & 32'h7; // @[CSR.scala 418:36]
  assign x67 = reg_mcountinhibit[2]; // @[CSR.scala 438:75]
  assign _GEN_23 = {{5'd0}, io_retire}; // @[Counters.scala 46:33]
  assign nextSmall = value_lo + _GEN_23; // @[Counters.scala 46:33]
  assign _GEN_0 = x67 ? {{1'd0}, value_lo} : nextSmall; // @[Counters.scala 47:19]
  assign _large_T_2 = nextSmall[6] & ~x67; // @[Counters.scala 51:33]
  assign _large_r_T_1 = value_hi + 58'h1; // @[Counters.scala 51:55]
  assign value = {value_hi,value_lo}; // @[Cat.scala 30:58]
  assign nextSmall_1 = value_lo_1 + _GEN_23; // @[Counters.scala 46:33]
  assign _GEN_2 = reg_mcountinhibit[0] ? {{1'd0}, value_lo_1} : nextSmall_1; // @[Counters.scala 47:19]
  assign _large_T_5 = nextSmall_1[6] & ~reg_mcountinhibit[0]; // @[Counters.scala 51:33]
  assign _large_r_T_3 = value_hi_1 + 58'h1; // @[Counters.scala 51:55]
  assign value_1 = {value_hi_1,value_lo_1}; // @[Cat.scala 30:58]
  assign mip_seip = reg_mip_seip | io_interrupts_seip; // @[CSR.scala 452:57]
  assign read_mip_lo = {io_interrupts_mtip,1'h0,reg_mip_stip,1'h0,io_interrupts_msip,1'h0,reg_mip_ssip,1'h0}; // @[CSR.scala 454:22]
  assign _read_mip_T = {4'h0,io_interrupts_meip,1'h0,mip_seip,1'h0,read_mip_lo}; // @[CSR.scala 454:22]
  assign read_mip = _read_mip_T & 16'haaa; // @[CSR.scala 454:29]
  reg [15:0] reg_mip; //SC
  assign reg_mip = read_mip;

  assign _GEN_45 = {{48'd0}, read_mip}; // @[CSR.scala 457:56]
  assign pending_interrupts = _GEN_45 & reg_mie; // @[CSR.scala 457:56]
  assign d_interrupts = {io_interrupts_debug, 14'h0}; // @[CSR.scala 458:42]
  assign _m_interrupts_T_1 = _delegate_T | reg_mstatus_mie; // @[CSR.scala 464:60]
  assign _m_interrupts_T_2 = nmie & _m_interrupts_T_1; // @[CSR.scala 464:31]
  assign _m_interrupts_T_4 = ~pending_interrupts | read_mideleg; // @[CSR.scala 464:103]
  assign m_interrupts = _m_interrupts_T_2 ? ~_m_interrupts_T_4 : 64'h0; // @[CSR.scala 464:25]
  assign _s_interrupts_T = reg_mstatus_prv < 2'h1; // @[CSR.scala 465:51]
  assign _s_interrupts_T_1 = reg_mstatus_prv == 2'h1; // @[CSR.scala 465:79]
  assign _s_interrupts_T_2 = _s_interrupts_T_1 & reg_mstatus_sie; // @[CSR.scala 465:89]
  assign _s_interrupts_T_3 = _s_interrupts_T | _s_interrupts_T_2; // @[CSR.scala 465:59]
  assign _s_interrupts_T_4 = nmie & _s_interrupts_T_3; // @[CSR.scala 465:31]
  assign _s_interrupts_T_5 = pending_interrupts & read_mideleg; // @[CSR.scala 465:130]
  assign s_interrupts = _s_interrupts_T_4 ? _s_interrupts_T_5 : 64'h0; // @[CSR.scala 465:25]
  assign _any_T_38 = d_interrupts[14] | d_interrupts[13]; // @[CSR.scala 1180:90]
  assign _any_T_39 = _any_T_38 | d_interrupts[12]; // @[CSR.scala 1180:90]
  assign _any_T_40 = _any_T_39 | d_interrupts[11]; // @[CSR.scala 1180:90]
  assign _any_T_41 = _any_T_40 | d_interrupts[3]; // @[CSR.scala 1180:90]
  assign _any_T_42 = _any_T_41 | d_interrupts[7]; // @[CSR.scala 1180:90]
  assign _any_T_43 = _any_T_42 | d_interrupts[9]; // @[CSR.scala 1180:90]
  assign _any_T_44 = _any_T_43 | d_interrupts[1]; // @[CSR.scala 1180:90]
  assign _any_T_45 = _any_T_44 | d_interrupts[5]; // @[CSR.scala 1180:90]
  assign _any_T_46 = _any_T_45 | d_interrupts[8]; // @[CSR.scala 1180:90]
  assign _any_T_47 = _any_T_46 | d_interrupts[0]; // @[CSR.scala 1180:90]
  assign _any_T_48 = _any_T_47 | d_interrupts[4]; // @[CSR.scala 1180:90]
  assign _any_T_50 = _any_T_48 | m_interrupts[15]; // @[CSR.scala 1180:90]
  assign _any_T_51 = _any_T_50 | m_interrupts[14]; // @[CSR.scala 1180:90]
  assign _any_T_52 = _any_T_51 | m_interrupts[13]; // @[CSR.scala 1180:90]
  assign _any_T_53 = _any_T_52 | m_interrupts[12]; // @[CSR.scala 1180:90]
  assign _any_T_54 = _any_T_53 | m_interrupts[11]; // @[CSR.scala 1180:90]
  assign _any_T_55 = _any_T_54 | m_interrupts[3]; // @[CSR.scala 1180:90]
  assign _any_T_56 = _any_T_55 | m_interrupts[7]; // @[CSR.scala 1180:90]
  assign _any_T_57 = _any_T_56 | m_interrupts[9]; // @[CSR.scala 1180:90]
  assign _any_T_58 = _any_T_57 | m_interrupts[1]; // @[CSR.scala 1180:90]
  assign _any_T_59 = _any_T_58 | m_interrupts[5]; // @[CSR.scala 1180:90]
  assign _any_T_60 = _any_T_59 | m_interrupts[8]; // @[CSR.scala 1180:90]
  assign _any_T_61 = _any_T_60 | m_interrupts[0]; // @[CSR.scala 1180:90]
  assign _any_T_62 = _any_T_61 | m_interrupts[4]; // @[CSR.scala 1180:90]
  assign _any_T_63 = _any_T_62 | s_interrupts[15]; // @[CSR.scala 1180:90]
  assign _any_T_64 = _any_T_63 | s_interrupts[14]; // @[CSR.scala 1180:90]
  assign _any_T_65 = _any_T_64 | s_interrupts[13]; // @[CSR.scala 1180:90]
  assign _any_T_66 = _any_T_65 | s_interrupts[12]; // @[CSR.scala 1180:90]
  assign _any_T_67 = _any_T_66 | s_interrupts[11]; // @[CSR.scala 1180:90]
  assign _any_T_68 = _any_T_67 | s_interrupts[3]; // @[CSR.scala 1180:90]
  assign _any_T_69 = _any_T_68 | s_interrupts[7]; // @[CSR.scala 1180:90]
  assign _any_T_70 = _any_T_69 | s_interrupts[9]; // @[CSR.scala 1180:90]
  assign _any_T_71 = _any_T_70 | s_interrupts[1]; // @[CSR.scala 1180:90]
  assign _any_T_72 = _any_T_71 | s_interrupts[5]; // @[CSR.scala 1180:90]
  assign _any_T_73 = _any_T_72 | s_interrupts[8]; // @[CSR.scala 1180:90]
  assign _any_T_74 = _any_T_73 | s_interrupts[0]; // @[CSR.scala 1180:90]
  assign anyInterrupt = _any_T_74 | s_interrupts[4]; // @[CSR.scala 1180:90]
  assign _which_T_38 = s_interrupts[0] ? 3'h0 : 3'h4; // @[Mux.scala 47:69]
  assign _which_T_39 = s_interrupts[8] ? 4'h8 : {{1'd0}, _which_T_38}; // @[Mux.scala 47:69]
  assign _which_T_40 = s_interrupts[5] ? 4'h5 : _which_T_39; // @[Mux.scala 47:69]
  assign _which_T_41 = s_interrupts[1] ? 4'h1 : _which_T_40; // @[Mux.scala 47:69]
  assign _which_T_42 = s_interrupts[9] ? 4'h9 : _which_T_41; // @[Mux.scala 47:69]
  assign _which_T_43 = s_interrupts[7] ? 4'h7 : _which_T_42; // @[Mux.scala 47:69]
  assign _which_T_44 = s_interrupts[3] ? 4'h3 : _which_T_43; // @[Mux.scala 47:69]
  assign _which_T_45 = s_interrupts[11] ? 4'hb : _which_T_44; // @[Mux.scala 47:69]
  assign _which_T_46 = s_interrupts[12] ? 4'hc : _which_T_45; // @[Mux.scala 47:69]
  assign _which_T_47 = s_interrupts[13] ? 4'hd : _which_T_46; // @[Mux.scala 47:69]
  assign _which_T_48 = s_interrupts[14] ? 4'he : _which_T_47; // @[Mux.scala 47:69]
  assign _which_T_49 = s_interrupts[15] ? 4'hf : _which_T_48; // @[Mux.scala 47:69]
  assign _which_T_50 = m_interrupts[4] ? 4'h4 : _which_T_49; // @[Mux.scala 47:69]
  assign _which_T_51 = m_interrupts[0] ? 4'h0 : _which_T_50; // @[Mux.scala 47:69]
  assign _which_T_52 = m_interrupts[8] ? 4'h8 : _which_T_51; // @[Mux.scala 47:69]
  assign _which_T_53 = m_interrupts[5] ? 4'h5 : _which_T_52; // @[Mux.scala 47:69]
  assign _which_T_54 = m_interrupts[1] ? 4'h1 : _which_T_53; // @[Mux.scala 47:69]
  assign _which_T_55 = m_interrupts[9] ? 4'h9 : _which_T_54; // @[Mux.scala 47:69]
  assign _which_T_56 = m_interrupts[7] ? 4'h7 : _which_T_55; // @[Mux.scala 47:69]
  assign _which_T_57 = m_interrupts[3] ? 4'h3 : _which_T_56; // @[Mux.scala 47:69]
  assign _which_T_58 = m_interrupts[11] ? 4'hb : _which_T_57; // @[Mux.scala 47:69]
  assign _which_T_59 = m_interrupts[12] ? 4'hc : _which_T_58; // @[Mux.scala 47:69]
  assign _which_T_60 = m_interrupts[13] ? 4'hd : _which_T_59; // @[Mux.scala 47:69]
  assign _which_T_61 = m_interrupts[14] ? 4'he : _which_T_60; // @[Mux.scala 47:69]
  assign _which_T_62 = m_interrupts[15] ? 4'hf : _which_T_61; // @[Mux.scala 47:69]
  assign _which_T_64 = d_interrupts[4] ? 4'h4 : _which_T_62; // @[Mux.scala 47:69]
  assign _which_T_65 = d_interrupts[0] ? 4'h0 : _which_T_64; // @[Mux.scala 47:69]
  assign _which_T_66 = d_interrupts[8] ? 4'h8 : _which_T_65; // @[Mux.scala 47:69]
  assign _which_T_67 = d_interrupts[5] ? 4'h5 : _which_T_66; // @[Mux.scala 47:69]
  assign _which_T_68 = d_interrupts[1] ? 4'h1 : _which_T_67; // @[Mux.scala 47:69]
  assign _which_T_69 = d_interrupts[9] ? 4'h9 : _which_T_68; // @[Mux.scala 47:69]
  assign _which_T_70 = d_interrupts[7] ? 4'h7 : _which_T_69; // @[Mux.scala 47:69]
  assign _which_T_71 = d_interrupts[3] ? 4'h3 : _which_T_70; // @[Mux.scala 47:69]
  assign _which_T_72 = d_interrupts[11] ? 4'hb : _which_T_71; // @[Mux.scala 47:69]
  assign _which_T_73 = d_interrupts[12] ? 4'hc : _which_T_72; // @[Mux.scala 47:69]
  assign _which_T_74 = d_interrupts[13] ? 4'hd : _which_T_73; // @[Mux.scala 47:69]
  assign whichInterrupt = d_interrupts[14] ? 4'he : _which_T_74; // @[Mux.scala 47:69]
  assign _GEN_556 = {{60'd0}, whichInterrupt}; // @[CSR.scala 468:67]
  assign _io_interrupt_T_1 = anyInterrupt & ~io_singleStep; // @[CSR.scala 469:33]
  assign _io_interrupt_T_2 = _io_interrupt_T_1 | reg_singleStepped; // @[CSR.scala 469:51]
  assign _io_interrupt_T_3 = reg_debug | io_status_cease; // @[CSR.scala 469:88]
  assign pmp_mask_base_lo = reg_pmp_0_cfg_a[0]; // @[PMP.scala 59:31]
  assign pmp_mask_base = {reg_pmp_0_addr,pmp_mask_base_lo}; // @[Cat.scala 30:58]
  assign _pmp_mask_T_1 = pmp_mask_base + 31'h1; // @[PMP.scala 60:23]
  assign pmp_mask_hi = pmp_mask_base & ~_pmp_mask_T_1; // @[PMP.scala 60:14]
  assign _pmp_mask_T_3 = {pmp_mask_hi,2'h3}; // @[Cat.scala 30:58]
  assign pmp_mask_base_lo_1 = reg_pmp_1_cfg_a[0]; // @[PMP.scala 59:31]
  assign pmp_mask_base_1 = {reg_pmp_1_addr,pmp_mask_base_lo_1}; // @[Cat.scala 30:58]
  assign _pmp_mask_T_5 = pmp_mask_base_1 + 31'h1; // @[PMP.scala 60:23]
  assign pmp_mask_hi_1 = pmp_mask_base_1 & ~_pmp_mask_T_5; // @[PMP.scala 60:14]
  assign _pmp_mask_T_7 = {pmp_mask_hi_1,2'h3}; // @[Cat.scala 30:58]
  assign pmp_mask_base_lo_2 = reg_pmp_2_cfg_a[0]; // @[PMP.scala 59:31]
  assign pmp_mask_base_2 = {reg_pmp_2_addr,pmp_mask_base_lo_2}; // @[Cat.scala 30:58]
  assign _pmp_mask_T_9 = pmp_mask_base_2 + 31'h1; // @[PMP.scala 60:23]
  assign pmp_mask_hi_2 = pmp_mask_base_2 & ~_pmp_mask_T_9; // @[PMP.scala 60:14]
  assign _pmp_mask_T_11 = {pmp_mask_hi_2,2'h3}; // @[Cat.scala 30:58]
  assign pmp_mask_base_lo_3 = reg_pmp_3_cfg_a[0]; // @[PMP.scala 59:31]
  assign pmp_mask_base_3 = {reg_pmp_3_addr,pmp_mask_base_lo_3}; // @[Cat.scala 30:58]
  assign _pmp_mask_T_13 = pmp_mask_base_3 + 31'h1; // @[PMP.scala 60:23]
  assign pmp_mask_hi_3 = pmp_mask_base_3 & ~_pmp_mask_T_13; // @[PMP.scala 60:14]
  assign _pmp_mask_T_15 = {pmp_mask_hi_3,2'h3}; // @[Cat.scala 30:58]
  assign pmp_mask_base_lo_4 = reg_pmp_4_cfg_a[0]; // @[PMP.scala 59:31]
  assign pmp_mask_base_4 = {reg_pmp_4_addr,pmp_mask_base_lo_4}; // @[Cat.scala 30:58]
  assign _pmp_mask_T_17 = pmp_mask_base_4 + 31'h1; // @[PMP.scala 60:23]
  assign pmp_mask_hi_4 = pmp_mask_base_4 & ~_pmp_mask_T_17; // @[PMP.scala 60:14]
  assign _pmp_mask_T_19 = {pmp_mask_hi_4,2'h3}; // @[Cat.scala 30:58]
  assign pmp_mask_base_lo_5 = reg_pmp_5_cfg_a[0]; // @[PMP.scala 59:31]
  assign pmp_mask_base_5 = {reg_pmp_5_addr,pmp_mask_base_lo_5}; // @[Cat.scala 30:58]
  assign _pmp_mask_T_21 = pmp_mask_base_5 + 31'h1; // @[PMP.scala 60:23]
  assign pmp_mask_hi_5 = pmp_mask_base_5 & ~_pmp_mask_T_21; // @[PMP.scala 60:14]
  assign _pmp_mask_T_23 = {pmp_mask_hi_5,2'h3}; // @[Cat.scala 30:58]
  assign pmp_mask_base_lo_6 = reg_pmp_6_cfg_a[0]; // @[PMP.scala 59:31]
  assign pmp_mask_base_6 = {reg_pmp_6_addr,pmp_mask_base_lo_6}; // @[Cat.scala 30:58]
  assign _pmp_mask_T_25 = pmp_mask_base_6 + 31'h1; // @[PMP.scala 60:23]
  assign pmp_mask_hi_6 = pmp_mask_base_6 & ~_pmp_mask_T_25; // @[PMP.scala 60:14]
  assign _pmp_mask_T_27 = {pmp_mask_hi_6,2'h3}; // @[Cat.scala 30:58]
  assign pmp_mask_base_lo_7 = reg_pmp_7_cfg_a[0]; // @[PMP.scala 59:31]
  assign pmp_mask_base_7 = {reg_pmp_7_addr,pmp_mask_base_lo_7}; // @[Cat.scala 30:58]
  assign _pmp_mask_T_29 = pmp_mask_base_7 + 31'h1; // @[PMP.scala 60:23]
  assign pmp_mask_hi_7 = pmp_mask_base_7 & ~_pmp_mask_T_29; // @[PMP.scala 60:14]
  assign _pmp_mask_T_31 = {pmp_mask_hi_7,2'h3}; // @[Cat.scala 30:58]
  assign read_mstatus_lo_lo = {io_status_hpie,io_status_spie,io_status_upie,io_status_mie,io_status_hie,io_status_sie,io_status_uie}; // @[CSR.scala 491:38]
  assign read_mstatus_lo = {io_status_sum,io_status_mprv,io_status_xs,io_status_fs,io_status_mpp,io_status_vs,io_status_spp,io_status_mpie,read_mstatus_lo_lo}; // @[CSR.scala 491:38]
  assign read_mstatus_hi_lo = {io_status_sxl,io_status_uxl,io_status_sd_rv32,io_status_zero1,io_status_tsr,io_status_tw,io_status_tvm,io_status_mxr}; // @[CSR.scala 491:38]
  assign _read_mstatus_T = {io_status_debug,io_status_cease,io_status_wfi,io_status_isa,io_status_dprv,io_status_prv,io_status_sd,io_status_zero2,read_mstatus_hi_lo,read_mstatus_lo}; // @[CSR.scala 491:38]
  reg [63:0] reg_mstatus;
  assign reg_mstatus = read_mstatus; //SC
  assign read_mstatus = _read_mstatus_T[63:0]; // @[CSR.scala 491:40]
  assign _read_mtvec_T_1 = reg_mtvec[0] ? 8'hfe : 8'h2; // @[CSR.scala 1209:39]
  assign _read_mtvec_T_3 = {{24'd0}, _read_mtvec_T_1}; // @[package.scala 165:41]
  assign read_mtvec_lo = reg_mtvec & ~_read_mtvec_T_3; // @[package.scala 165:35]
  assign read_mtvec = {32'h0,read_mtvec_lo}; // @[Cat.scala 30:58]
  assign _read_stvec_T_1 = reg_stvec[0] ? 8'hfe : 8'h2; // @[CSR.scala 1209:39]
  assign _read_stvec_T_3 = {{31'd0}, _read_stvec_T_1}; // @[package.scala 165:41]
  assign read_stvec_lo = reg_stvec & ~_read_stvec_T_3; // @[package.scala 165:35]
  assign read_stvec_hi = read_stvec_lo[38] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  assign read_stvec = {read_stvec_hi,read_stvec_lo}; // @[Cat.scala 30:58]
  assign lo_2 = {reg_bp_0_control_m,1'h0,reg_bp_0_control_s,reg_bp_0_control_u,reg_bp_0_control_x,reg_bp_0_control_w,reg_bp_0_control_r}; // @[CSR.scala 497:48]
  assign _T_7 = {4'h2,reg_bp_0_control_dmode,46'h40000000000,reg_bp_0_control_action,1'h0,2'h0,reg_bp_0_control_tmatch,lo_2}; // @[CSR.scala 497:48]
  assign hi_3 = reg_bp_0_address[38] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  assign _T_10 = {hi_3,reg_bp_0_address}; // @[Cat.scala 30:58]
  assign _T_14 = reg_misa[2] ? 2'h1 : 2'h3; // @[CSR.scala 1208:36]
  assign _GEN_557 = {{38'd0}, _T_14}; // @[CSR.scala 1208:31]
  assign _T_15 = ~reg_mepc | _GEN_557; // @[CSR.scala 1208:31]
  assign lo_4 = ~_T_15; // @[CSR.scala 1208:26]
  assign hi_5 = lo_4[39] ? 24'hffffff : 24'h0; // @[Bitwise.scala 72:12]
  assign _T_18 = {hi_5,lo_4}; // @[Cat.scala 30:58]
  assign hi_6 = reg_mtval[39] ? 24'hffffff : 24'h0; // @[Bitwise.scala 72:12]
  assign _T_21 = {hi_6,reg_mtval}; // @[Cat.scala 30:58]
  assign lo_5 = {2'h0,1'h0,reg_dcsr_cause,3'h0,reg_dcsr_step,reg_dcsr_prv}; // @[CSR.scala 512:27]
  assign _T_22 = {4'h4,12'h0,reg_dcsr_ebreakm,1'h0,reg_dcsr_ebreaks,reg_dcsr_ebreaku,lo_5}; // @[CSR.scala 512:27]
  reg [31:0] reg_dcsr; //SC
  assign reg_dcsr = _T_22;
  assign _T_26 = ~reg_dpc | _GEN_557; // @[CSR.scala 1208:31]
  assign lo_6 = ~_T_26; // @[CSR.scala 1208:26]
  assign hi_8 = lo_6[39] ? 24'hffffff : 24'h0; // @[Bitwise.scala 72:12]
  assign _T_29 = {hi_8,lo_6}; // @[Cat.scala 30:58]
  reg [7:0] reg_fcsr ; //SC
  assign reg_fcsr = read_fcsr;
  assign read_fcsr = {reg_frm,reg_fflags}; // @[Cat.scala 30:58]
  assign read_sie = reg_mie & read_mideleg; // @[CSR.scala 584:28]
  assign read_sip = _GEN_45 & read_mideleg; // @[CSR.scala 585:29]
  assign lo_lo_4 = {1'h0,io_status_spie,2'h0,1'h0,io_status_sie,1'h0}; // @[CSR.scala 599:57]
  assign lo_7 = {io_status_sum,1'h0,io_status_xs,io_status_fs,2'h0,io_status_vs,io_status_spp,1'h0,lo_lo_4}; // @[CSR.scala 599:57]
  assign hi_lo_4 = {2'h0,io_status_uxl,io_status_sd_rv32,8'h0,2'h0,1'h0,io_status_mxr}; // @[CSR.scala 599:57]
  assign _T_30 = {35'h0,4'h0,io_status_sd,27'h0,hi_lo_4,lo_7}; // @[CSR.scala 599:57]
  assign hi_10 = reg_stval[39] ? 24'hffffff : 24'h0; // @[Bitwise.scala 72:12]
  assign _T_34 = {hi_10,reg_stval}; // @[Cat.scala 30:58]
  reg [63:0] reg_satp;
  assign reg_satp = _T_35;
  assign _T_35 = {reg_satp_mode,16'h0,reg_satp_ppn}; // @[CSR.scala 605:43]
  
  assign _T_39 = ~reg_sepc | _GEN_557; // @[CSR.scala 1208:31]
  assign lo_8 = ~_T_39; // @[CSR.scala 1208:26]
  assign hi_12 = lo_8[39] ? 24'hffffff : 24'h0; // @[Bitwise.scala 72:12]
  assign _T_42 = {hi_12,lo_8}; // @[Cat.scala 30:58]
  assign lo_lo_lo_3 = {reg_pmp_0_cfg_l,2'h0,reg_pmp_0_cfg_a,reg_pmp_0_cfg_x,reg_pmp_0_cfg_w,reg_pmp_0_cfg_r}; // @[package.scala 36:38]
  assign lo_hi_lo_5 = {reg_pmp_2_cfg_l,2'h0,reg_pmp_2_cfg_a,reg_pmp_2_cfg_x,reg_pmp_2_cfg_w,reg_pmp_2_cfg_r}; // @[package.scala 36:38]
  assign hi_lo_lo_4 = {reg_pmp_4_cfg_l,2'h0,reg_pmp_4_cfg_a,reg_pmp_4_cfg_x,reg_pmp_4_cfg_w,reg_pmp_4_cfg_r}; // @[package.scala 36:38]
  assign hi_hi_lo_5 = {reg_pmp_6_cfg_l,2'h0,reg_pmp_6_cfg_a,reg_pmp_6_cfg_x,reg_pmp_6_cfg_w,reg_pmp_6_cfg_r}; // @[package.scala 36:38]
  assign lo_lo_5 = {reg_pmp_1_cfg_l,2'h0,reg_pmp_1_cfg_a,reg_pmp_1_cfg_x,reg_pmp_1_cfg_w,reg_pmp_1_cfg_r,lo_lo_lo_3}; // @[Cat.scala 30:58]
  assign lo_17 = {reg_pmp_3_cfg_l,2'h0,reg_pmp_3_cfg_a,reg_pmp_3_cfg_x,reg_pmp_3_cfg_w,reg_pmp_3_cfg_r,lo_hi_lo_5,lo_lo_5}; // @[Cat.scala 30:58]
  assign hi_lo_5 = {reg_pmp_5_cfg_l,2'h0,reg_pmp_5_cfg_a,reg_pmp_5_cfg_x,reg_pmp_5_cfg_w,reg_pmp_5_cfg_r,hi_lo_lo_4}; // @[Cat.scala 30:58]
  assign _T_43 = {reg_pmp_7_cfg_l,2'h0,reg_pmp_7_cfg_a,reg_pmp_7_cfg_x,reg_pmp_7_cfg_w,reg_pmp_7_cfg_r,hi_hi_lo_5,hi_lo_5,lo_17}; // @[Cat.scala 30:58]
  reg [63:0] pmpcfg0; //SC
  assign pmpcfg0 = _T_43;
  assign _T_46 = io_rw_addr == 12'h7a1; // @[CSR.scala 636:73]
  assign _T_47 = io_rw_addr == 12'h7a2; // @[CSR.scala 636:73]
  assign _T_49 = io_rw_addr == 12'h301; // @[CSR.scala 636:73]
  assign _T_50 = io_rw_addr == 12'h300; // @[CSR.scala 636:73]
  assign _T_51 = io_rw_addr == 12'h305; // @[CSR.scala 636:73]
  assign _T_52 = io_rw_addr == 12'h344; // @[CSR.scala 636:73]
  assign _T_53 = io_rw_addr == 12'h304; // @[CSR.scala 636:73]
  assign _T_54 = io_rw_addr == 12'h340; // @[CSR.scala 636:73]
  assign _T_55 = io_rw_addr == 12'h341; // @[CSR.scala 636:73]
  assign _T_56 = io_rw_addr == 12'h343; // @[CSR.scala 636:73]
  assign _T_57 = io_rw_addr == 12'h342; // @[CSR.scala 636:73]
  assign _T_58 = io_rw_addr == 12'hf14; // @[CSR.scala 636:73]
  assign _T_59 = io_rw_addr == 12'h7b0; // @[CSR.scala 636:73]
  assign _T_60 = io_rw_addr == 12'h7b1; // @[CSR.scala 636:73]
  assign _T_61 = io_rw_addr == 12'h7b2; // @[CSR.scala 636:73]
  assign _T_62 = io_rw_addr == 12'h1; // @[CSR.scala 636:73]
  assign _T_63 = io_rw_addr == 12'h2; // @[CSR.scala 636:73]
  assign _T_64 = io_rw_addr == 12'h3; // @[CSR.scala 636:73]
  assign _T_65 = io_rw_addr == 12'h320; // @[CSR.scala 636:73]
  assign _T_66 = io_rw_addr == 12'hb00; // @[CSR.scala 636:73]
  assign _T_67 = io_rw_addr == 12'hb02; // @[CSR.scala 636:73]
  assign _T_155 = io_rw_addr == 12'h306; // @[CSR.scala 636:73]
  assign _T_156 = io_rw_addr == 12'hc00; // @[CSR.scala 636:73]
  assign _T_157 = io_rw_addr == 12'hc02; // @[CSR.scala 636:73]
  assign _T_158 = io_rw_addr == 12'h100; // @[CSR.scala 636:73]
  assign _T_159 = io_rw_addr == 12'h144; // @[CSR.scala 636:73]
  assign _T_160 = io_rw_addr == 12'h104; // @[CSR.scala 636:73]
  assign _T_161 = io_rw_addr == 12'h140; // @[CSR.scala 636:73]
  assign _T_162 = io_rw_addr == 12'h142; // @[CSR.scala 636:73]
  assign _T_163 = io_rw_addr == 12'h143; // @[CSR.scala 636:73]
  assign _T_164 = io_rw_addr == 12'h180; // @[CSR.scala 636:73]
  assign _T_165 = io_rw_addr == 12'h141; // @[CSR.scala 636:73]
  assign _T_166 = io_rw_addr == 12'h105; // @[CSR.scala 636:73]
  assign _T_167 = io_rw_addr == 12'h106; // @[CSR.scala 636:73]
  assign _T_168 = io_rw_addr == 12'h303; // @[CSR.scala 636:73]
  assign _T_169 = io_rw_addr == 12'h302; // @[CSR.scala 636:73]
  assign _T_170 = io_rw_addr == 12'h3a0; // @[CSR.scala 636:73]
  assign _T_172 = io_rw_addr == 12'h3b0; // @[CSR.scala 636:73]
  assign _T_173 = io_rw_addr == 12'h3b1; // @[CSR.scala 636:73]
  assign _T_174 = io_rw_addr == 12'h3b2; // @[CSR.scala 636:73]
  assign _T_175 = io_rw_addr == 12'h3b3; // @[CSR.scala 636:73]
  assign _T_176 = io_rw_addr == 12'h3b4; // @[CSR.scala 636:73]
  assign _T_177 = io_rw_addr == 12'h3b5; // @[CSR.scala 636:73]
  assign _T_178 = io_rw_addr == 12'h3b6; // @[CSR.scala 636:73]
  assign _T_179 = io_rw_addr == 12'h3b7; // @[CSR.scala 636:73]
  assign _T_188 = io_rw_addr == 12'h7c1; // @[CSR.scala 636:73]
  assign _T_189 = io_rw_addr == 12'hf12; // @[CSR.scala 636:73]
  assign _T_191 = io_rw_addr == 12'hf13; // @[CSR.scala 636:73]
  assign _wdata_T_1 = io_rw_cmd[1] ? io_rw_rdata : 64'h0; // @[CSR.scala 1186:9]
  assign _wdata_T_2 = _wdata_T_1 | io_rw_wdata; // @[CSR.scala 1186:34]
  assign _wdata_T_4 = &io_rw_cmd[1:0]; // @[CSR.scala 1186:59]
  assign _wdata_T_5 = _wdata_T_4 ? io_rw_wdata : 64'h0; // @[CSR.scala 1186:49]
  assign wdata = _wdata_T_2 & ~_wdata_T_5; // @[CSR.scala 1186:43]
  assign _T_205 = _T_192 & 32'h20200000; // @[Decode.scala 14:65]
  assign _T_206 = _T_205 == 32'h20000000; // @[Decode.scala 14:121]
  assign _T_208 = _T_192 & 32'h32200000; // @[Decode.scala 14:65]
  assign _T_209 = _T_208 == 32'h10000000; // @[Decode.scala 14:121]
  assign insn_cease = system_insn & _T_206; // @[CSR.scala 652:95]
  assign insn_wfi = system_insn & _T_209; // @[CSR.scala 652:95]
  assign _T_220 = {io_decode_0_csr, 20'h0}; // @[CSR.scala 659:30]
  assign _T_227 = _T_220 & 32'h12400000; // @[Decode.scala 14:65]
  assign _T_228 = _T_227 == 32'h10000000; // @[Decode.scala 14:121]
  assign _T_229 = _T_220 & 32'h40000000; // @[Decode.scala 14:65]
  assign _T_230 = _T_229 == 32'h40000000; // @[Decode.scala 14:121]
  assign is_ret = _T_228 | _T_230; // @[Decode.scala 15:30]
  assign _T_236 = _T_220 & 32'h32200000; // @[Decode.scala 14:65]
  assign is_wfi = _T_236 == 32'h10000000; // @[Decode.scala 14:121]
  assign _T_239 = _T_220 & 32'h42000000; // @[Decode.scala 14:65]
  assign is_sfence = _T_239 == 32'h2000000; // @[Decode.scala 14:121]
  assign _allow_wfi_T = reg_mstatus_prv > 2'h1; // @[CSR.scala 661:63]
  assign allow_wfi = _allow_wfi_T | ~reg_mstatus_tw; // @[CSR.scala 661:71]
  assign allow_sfence_vma = _allow_wfi_T | ~reg_mstatus_tvm; // @[CSR.scala 662:70]
  assign allow_sret = _allow_wfi_T | ~reg_mstatus_tsr; // @[CSR.scala 663:72]
  assign counter_addr = io_decode_0_csr[4:0]; // @[CSR.scala 664:34]
  assign _allow_counter_T_1 = read_mcounteren >> counter_addr; // @[CSR.scala 665:68]
  assign _allow_counter_T_3 = _allow_wfi_T | _allow_counter_T_1[0]; // @[CSR.scala 665:50]
  assign _allow_counter_T_4 = reg_mstatus_prv >= 2'h1; // @[CSR.scala 666:44]
  assign _allow_counter_T_6 = read_scounteren >> counter_addr; // @[CSR.scala 666:71]
  assign _allow_counter_T_8 = _allow_counter_T_4 | _allow_counter_T_6[0]; // @[CSR.scala 666:53]
  assign allow_counter = _allow_counter_T_3 & _allow_counter_T_8; // @[CSR.scala 665:84]
  assign _io_decode_0_fp_illegal_T = io_status_fs == 2'h0; // @[CSR.scala 667:39]
  assign _io_decode_0_fp_csr_T = io_decode_0_csr & 12'h900; // @[Decode.scala 14:65]
  assign _io_decode_0_read_illegal_T_1 = reg_mstatus_prv < io_decode_0_csr[9:8]; // @[CSR.scala 671:44]
  assign _io_decode_0_read_illegal_T_2 = io_decode_0_csr == 12'h7a0; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_3 = io_decode_0_csr == 12'h7a1; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_4 = io_decode_0_csr == 12'h7a2; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_5 = io_decode_0_csr == 12'h7a3; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_6 = io_decode_0_csr == 12'h301; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_7 = io_decode_0_csr == 12'h300; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_8 = io_decode_0_csr == 12'h305; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_9 = io_decode_0_csr == 12'h344; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_10 = io_decode_0_csr == 12'h304; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_11 = io_decode_0_csr == 12'h340; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_12 = io_decode_0_csr == 12'h341; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_13 = io_decode_0_csr == 12'h343; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_14 = io_decode_0_csr == 12'h342; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_15 = io_decode_0_csr == 12'hf14; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_16 = io_decode_0_csr == 12'h7b0; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_17 = io_decode_0_csr == 12'h7b1; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_18 = io_decode_0_csr == 12'h7b2; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_19 = io_decode_0_csr == 12'h1; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_20 = io_decode_0_csr == 12'h2; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_21 = io_decode_0_csr == 12'h3; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_22 = io_decode_0_csr == 12'h320; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_23 = io_decode_0_csr == 12'hb00; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_24 = io_decode_0_csr == 12'hb02; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_25 = io_decode_0_csr == 12'h323; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_26 = io_decode_0_csr == 12'hb03; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_27 = io_decode_0_csr == 12'hc03; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_28 = io_decode_0_csr == 12'h324; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_29 = io_decode_0_csr == 12'hb04; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_30 = io_decode_0_csr == 12'hc04; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_31 = io_decode_0_csr == 12'h325; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_32 = io_decode_0_csr == 12'hb05; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_33 = io_decode_0_csr == 12'hc05; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_34 = io_decode_0_csr == 12'h326; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_35 = io_decode_0_csr == 12'hb06; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_36 = io_decode_0_csr == 12'hc06; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_37 = io_decode_0_csr == 12'h327; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_38 = io_decode_0_csr == 12'hb07; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_39 = io_decode_0_csr == 12'hc07; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_40 = io_decode_0_csr == 12'h328; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_41 = io_decode_0_csr == 12'hb08; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_42 = io_decode_0_csr == 12'hc08; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_43 = io_decode_0_csr == 12'h329; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_44 = io_decode_0_csr == 12'hb09; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_45 = io_decode_0_csr == 12'hc09; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_46 = io_decode_0_csr == 12'h32a; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_47 = io_decode_0_csr == 12'hb0a; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_48 = io_decode_0_csr == 12'hc0a; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_49 = io_decode_0_csr == 12'h32b; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_50 = io_decode_0_csr == 12'hb0b; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_51 = io_decode_0_csr == 12'hc0b; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_52 = io_decode_0_csr == 12'h32c; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_53 = io_decode_0_csr == 12'hb0c; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_54 = io_decode_0_csr == 12'hc0c; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_55 = io_decode_0_csr == 12'h32d; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_56 = io_decode_0_csr == 12'hb0d; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_57 = io_decode_0_csr == 12'hc0d; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_58 = io_decode_0_csr == 12'h32e; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_59 = io_decode_0_csr == 12'hb0e; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_60 = io_decode_0_csr == 12'hc0e; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_61 = io_decode_0_csr == 12'h32f; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_62 = io_decode_0_csr == 12'hb0f; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_63 = io_decode_0_csr == 12'hc0f; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_64 = io_decode_0_csr == 12'h330; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_65 = io_decode_0_csr == 12'hb10; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_66 = io_decode_0_csr == 12'hc10; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_67 = io_decode_0_csr == 12'h331; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_68 = io_decode_0_csr == 12'hb11; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_69 = io_decode_0_csr == 12'hc11; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_70 = io_decode_0_csr == 12'h332; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_71 = io_decode_0_csr == 12'hb12; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_72 = io_decode_0_csr == 12'hc12; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_73 = io_decode_0_csr == 12'h333; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_74 = io_decode_0_csr == 12'hb13; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_75 = io_decode_0_csr == 12'hc13; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_76 = io_decode_0_csr == 12'h334; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_77 = io_decode_0_csr == 12'hb14; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_78 = io_decode_0_csr == 12'hc14; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_79 = io_decode_0_csr == 12'h335; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_80 = io_decode_0_csr == 12'hb15; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_81 = io_decode_0_csr == 12'hc15; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_82 = io_decode_0_csr == 12'h336; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_83 = io_decode_0_csr == 12'hb16; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_84 = io_decode_0_csr == 12'hc16; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_85 = io_decode_0_csr == 12'h337; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_86 = io_decode_0_csr == 12'hb17; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_87 = io_decode_0_csr == 12'hc17; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_88 = io_decode_0_csr == 12'h338; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_89 = io_decode_0_csr == 12'hb18; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_90 = io_decode_0_csr == 12'hc18; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_91 = io_decode_0_csr == 12'h339; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_92 = io_decode_0_csr == 12'hb19; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_93 = io_decode_0_csr == 12'hc19; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_94 = io_decode_0_csr == 12'h33a; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_95 = io_decode_0_csr == 12'hb1a; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_96 = io_decode_0_csr == 12'hc1a; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_97 = io_decode_0_csr == 12'h33b; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_98 = io_decode_0_csr == 12'hb1b; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_99 = io_decode_0_csr == 12'hc1b; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_100 = io_decode_0_csr == 12'h33c; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_101 = io_decode_0_csr == 12'hb1c; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_102 = io_decode_0_csr == 12'hc1c; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_103 = io_decode_0_csr == 12'h33d; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_104 = io_decode_0_csr == 12'hb1d; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_105 = io_decode_0_csr == 12'hc1d; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_106 = io_decode_0_csr == 12'h33e; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_107 = io_decode_0_csr == 12'hb1e; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_108 = io_decode_0_csr == 12'hc1e; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_109 = io_decode_0_csr == 12'h33f; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_110 = io_decode_0_csr == 12'hb1f; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_111 = io_decode_0_csr == 12'hc1f; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_112 = io_decode_0_csr == 12'h306; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_113 = io_decode_0_csr == 12'hc00; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_114 = io_decode_0_csr == 12'hc02; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_115 = io_decode_0_csr == 12'h100; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_116 = io_decode_0_csr == 12'h144; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_117 = io_decode_0_csr == 12'h104; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_118 = io_decode_0_csr == 12'h140; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_119 = io_decode_0_csr == 12'h142; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_120 = io_decode_0_csr == 12'h143; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_121 = io_decode_0_csr == 12'h180; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_122 = io_decode_0_csr == 12'h141; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_123 = io_decode_0_csr == 12'h105; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_124 = io_decode_0_csr == 12'h106; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_125 = io_decode_0_csr == 12'h303; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_126 = io_decode_0_csr == 12'h302; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_127 = io_decode_0_csr == 12'h3a0; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_128 = io_decode_0_csr == 12'h3a2; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_129 = io_decode_0_csr == 12'h3b0; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_130 = io_decode_0_csr == 12'h3b1; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_131 = io_decode_0_csr == 12'h3b2; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_132 = io_decode_0_csr == 12'h3b3; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_133 = io_decode_0_csr == 12'h3b4; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_134 = io_decode_0_csr == 12'h3b5; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_135 = io_decode_0_csr == 12'h3b6; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_136 = io_decode_0_csr == 12'h3b7; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_137 = io_decode_0_csr == 12'h3b8; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_138 = io_decode_0_csr == 12'h3b9; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_139 = io_decode_0_csr == 12'h3ba; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_140 = io_decode_0_csr == 12'h3bb; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_141 = io_decode_0_csr == 12'h3bc; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_142 = io_decode_0_csr == 12'h3bd; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_143 = io_decode_0_csr == 12'h3be; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_144 = io_decode_0_csr == 12'h3bf; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_145 = io_decode_0_csr == 12'h7c1; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_146 = io_decode_0_csr == 12'hf12; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_147 = io_decode_0_csr == 12'hf11; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_148 = io_decode_0_csr == 12'hf13; // @[CSR.scala 655:99]
  assign _io_decode_0_read_illegal_T_149 = _io_decode_0_read_illegal_T_2 | _io_decode_0_read_illegal_T_3; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_150 = _io_decode_0_read_illegal_T_149 | _io_decode_0_read_illegal_T_4; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_151 = _io_decode_0_read_illegal_T_150 | _io_decode_0_read_illegal_T_5; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_152 = _io_decode_0_read_illegal_T_151 | _io_decode_0_read_illegal_T_6; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_153 = _io_decode_0_read_illegal_T_152 | _io_decode_0_read_illegal_T_7; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_154 = _io_decode_0_read_illegal_T_153 | _io_decode_0_read_illegal_T_8; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_155 = _io_decode_0_read_illegal_T_154 | _io_decode_0_read_illegal_T_9; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_156 = _io_decode_0_read_illegal_T_155 | _io_decode_0_read_illegal_T_10; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_157 = _io_decode_0_read_illegal_T_156 | _io_decode_0_read_illegal_T_11; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_158 = _io_decode_0_read_illegal_T_157 | _io_decode_0_read_illegal_T_12; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_159 = _io_decode_0_read_illegal_T_158 | _io_decode_0_read_illegal_T_13; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_160 = _io_decode_0_read_illegal_T_159 | _io_decode_0_read_illegal_T_14; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_161 = _io_decode_0_read_illegal_T_160 | _io_decode_0_read_illegal_T_15; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_162 = _io_decode_0_read_illegal_T_161 | _io_decode_0_read_illegal_T_16; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_163 = _io_decode_0_read_illegal_T_162 | _io_decode_0_read_illegal_T_17; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_164 = _io_decode_0_read_illegal_T_163 | _io_decode_0_read_illegal_T_18; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_165 = _io_decode_0_read_illegal_T_164 | _io_decode_0_read_illegal_T_19; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_166 = _io_decode_0_read_illegal_T_165 | _io_decode_0_read_illegal_T_20; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_167 = _io_decode_0_read_illegal_T_166 | _io_decode_0_read_illegal_T_21; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_168 = _io_decode_0_read_illegal_T_167 | _io_decode_0_read_illegal_T_22; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_169 = _io_decode_0_read_illegal_T_168 | _io_decode_0_read_illegal_T_23; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_170 = _io_decode_0_read_illegal_T_169 | _io_decode_0_read_illegal_T_24; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_171 = _io_decode_0_read_illegal_T_170 | _io_decode_0_read_illegal_T_25; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_172 = _io_decode_0_read_illegal_T_171 | _io_decode_0_read_illegal_T_26; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_173 = _io_decode_0_read_illegal_T_172 | _io_decode_0_read_illegal_T_27; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_174 = _io_decode_0_read_illegal_T_173 | _io_decode_0_read_illegal_T_28; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_175 = _io_decode_0_read_illegal_T_174 | _io_decode_0_read_illegal_T_29; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_176 = _io_decode_0_read_illegal_T_175 | _io_decode_0_read_illegal_T_30; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_177 = _io_decode_0_read_illegal_T_176 | _io_decode_0_read_illegal_T_31; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_178 = _io_decode_0_read_illegal_T_177 | _io_decode_0_read_illegal_T_32; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_179 = _io_decode_0_read_illegal_T_178 | _io_decode_0_read_illegal_T_33; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_180 = _io_decode_0_read_illegal_T_179 | _io_decode_0_read_illegal_T_34; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_181 = _io_decode_0_read_illegal_T_180 | _io_decode_0_read_illegal_T_35; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_182 = _io_decode_0_read_illegal_T_181 | _io_decode_0_read_illegal_T_36; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_183 = _io_decode_0_read_illegal_T_182 | _io_decode_0_read_illegal_T_37; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_184 = _io_decode_0_read_illegal_T_183 | _io_decode_0_read_illegal_T_38; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_185 = _io_decode_0_read_illegal_T_184 | _io_decode_0_read_illegal_T_39; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_186 = _io_decode_0_read_illegal_T_185 | _io_decode_0_read_illegal_T_40; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_187 = _io_decode_0_read_illegal_T_186 | _io_decode_0_read_illegal_T_41; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_188 = _io_decode_0_read_illegal_T_187 | _io_decode_0_read_illegal_T_42; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_189 = _io_decode_0_read_illegal_T_188 | _io_decode_0_read_illegal_T_43; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_190 = _io_decode_0_read_illegal_T_189 | _io_decode_0_read_illegal_T_44; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_191 = _io_decode_0_read_illegal_T_190 | _io_decode_0_read_illegal_T_45; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_192 = _io_decode_0_read_illegal_T_191 | _io_decode_0_read_illegal_T_46; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_193 = _io_decode_0_read_illegal_T_192 | _io_decode_0_read_illegal_T_47; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_194 = _io_decode_0_read_illegal_T_193 | _io_decode_0_read_illegal_T_48; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_195 = _io_decode_0_read_illegal_T_194 | _io_decode_0_read_illegal_T_49; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_196 = _io_decode_0_read_illegal_T_195 | _io_decode_0_read_illegal_T_50; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_197 = _io_decode_0_read_illegal_T_196 | _io_decode_0_read_illegal_T_51; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_198 = _io_decode_0_read_illegal_T_197 | _io_decode_0_read_illegal_T_52; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_199 = _io_decode_0_read_illegal_T_198 | _io_decode_0_read_illegal_T_53; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_200 = _io_decode_0_read_illegal_T_199 | _io_decode_0_read_illegal_T_54; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_201 = _io_decode_0_read_illegal_T_200 | _io_decode_0_read_illegal_T_55; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_202 = _io_decode_0_read_illegal_T_201 | _io_decode_0_read_illegal_T_56; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_203 = _io_decode_0_read_illegal_T_202 | _io_decode_0_read_illegal_T_57; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_204 = _io_decode_0_read_illegal_T_203 | _io_decode_0_read_illegal_T_58; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_205 = _io_decode_0_read_illegal_T_204 | _io_decode_0_read_illegal_T_59; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_206 = _io_decode_0_read_illegal_T_205 | _io_decode_0_read_illegal_T_60; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_207 = _io_decode_0_read_illegal_T_206 | _io_decode_0_read_illegal_T_61; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_208 = _io_decode_0_read_illegal_T_207 | _io_decode_0_read_illegal_T_62; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_209 = _io_decode_0_read_illegal_T_208 | _io_decode_0_read_illegal_T_63; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_210 = _io_decode_0_read_illegal_T_209 | _io_decode_0_read_illegal_T_64; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_211 = _io_decode_0_read_illegal_T_210 | _io_decode_0_read_illegal_T_65; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_212 = _io_decode_0_read_illegal_T_211 | _io_decode_0_read_illegal_T_66; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_213 = _io_decode_0_read_illegal_T_212 | _io_decode_0_read_illegal_T_67; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_214 = _io_decode_0_read_illegal_T_213 | _io_decode_0_read_illegal_T_68; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_215 = _io_decode_0_read_illegal_T_214 | _io_decode_0_read_illegal_T_69; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_216 = _io_decode_0_read_illegal_T_215 | _io_decode_0_read_illegal_T_70; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_217 = _io_decode_0_read_illegal_T_216 | _io_decode_0_read_illegal_T_71; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_218 = _io_decode_0_read_illegal_T_217 | _io_decode_0_read_illegal_T_72; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_219 = _io_decode_0_read_illegal_T_218 | _io_decode_0_read_illegal_T_73; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_220 = _io_decode_0_read_illegal_T_219 | _io_decode_0_read_illegal_T_74; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_221 = _io_decode_0_read_illegal_T_220 | _io_decode_0_read_illegal_T_75; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_222 = _io_decode_0_read_illegal_T_221 | _io_decode_0_read_illegal_T_76; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_223 = _io_decode_0_read_illegal_T_222 | _io_decode_0_read_illegal_T_77; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_224 = _io_decode_0_read_illegal_T_223 | _io_decode_0_read_illegal_T_78; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_225 = _io_decode_0_read_illegal_T_224 | _io_decode_0_read_illegal_T_79; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_226 = _io_decode_0_read_illegal_T_225 | _io_decode_0_read_illegal_T_80; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_227 = _io_decode_0_read_illegal_T_226 | _io_decode_0_read_illegal_T_81; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_228 = _io_decode_0_read_illegal_T_227 | _io_decode_0_read_illegal_T_82; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_229 = _io_decode_0_read_illegal_T_228 | _io_decode_0_read_illegal_T_83; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_230 = _io_decode_0_read_illegal_T_229 | _io_decode_0_read_illegal_T_84; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_231 = _io_decode_0_read_illegal_T_230 | _io_decode_0_read_illegal_T_85; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_232 = _io_decode_0_read_illegal_T_231 | _io_decode_0_read_illegal_T_86; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_233 = _io_decode_0_read_illegal_T_232 | _io_decode_0_read_illegal_T_87; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_234 = _io_decode_0_read_illegal_T_233 | _io_decode_0_read_illegal_T_88; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_235 = _io_decode_0_read_illegal_T_234 | _io_decode_0_read_illegal_T_89; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_236 = _io_decode_0_read_illegal_T_235 | _io_decode_0_read_illegal_T_90; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_237 = _io_decode_0_read_illegal_T_236 | _io_decode_0_read_illegal_T_91; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_238 = _io_decode_0_read_illegal_T_237 | _io_decode_0_read_illegal_T_92; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_239 = _io_decode_0_read_illegal_T_238 | _io_decode_0_read_illegal_T_93; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_240 = _io_decode_0_read_illegal_T_239 | _io_decode_0_read_illegal_T_94; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_241 = _io_decode_0_read_illegal_T_240 | _io_decode_0_read_illegal_T_95; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_242 = _io_decode_0_read_illegal_T_241 | _io_decode_0_read_illegal_T_96; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_243 = _io_decode_0_read_illegal_T_242 | _io_decode_0_read_illegal_T_97; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_244 = _io_decode_0_read_illegal_T_243 | _io_decode_0_read_illegal_T_98; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_245 = _io_decode_0_read_illegal_T_244 | _io_decode_0_read_illegal_T_99; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_246 = _io_decode_0_read_illegal_T_245 | _io_decode_0_read_illegal_T_100; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_247 = _io_decode_0_read_illegal_T_246 | _io_decode_0_read_illegal_T_101; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_248 = _io_decode_0_read_illegal_T_247 | _io_decode_0_read_illegal_T_102; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_249 = _io_decode_0_read_illegal_T_248 | _io_decode_0_read_illegal_T_103; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_250 = _io_decode_0_read_illegal_T_249 | _io_decode_0_read_illegal_T_104; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_251 = _io_decode_0_read_illegal_T_250 | _io_decode_0_read_illegal_T_105; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_252 = _io_decode_0_read_illegal_T_251 | _io_decode_0_read_illegal_T_106; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_253 = _io_decode_0_read_illegal_T_252 | _io_decode_0_read_illegal_T_107; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_254 = _io_decode_0_read_illegal_T_253 | _io_decode_0_read_illegal_T_108; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_255 = _io_decode_0_read_illegal_T_254 | _io_decode_0_read_illegal_T_109; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_256 = _io_decode_0_read_illegal_T_255 | _io_decode_0_read_illegal_T_110; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_257 = _io_decode_0_read_illegal_T_256 | _io_decode_0_read_illegal_T_111; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_258 = _io_decode_0_read_illegal_T_257 | _io_decode_0_read_illegal_T_112; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_259 = _io_decode_0_read_illegal_T_258 | _io_decode_0_read_illegal_T_113; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_260 = _io_decode_0_read_illegal_T_259 | _io_decode_0_read_illegal_T_114; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_261 = _io_decode_0_read_illegal_T_260 | _io_decode_0_read_illegal_T_115; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_262 = _io_decode_0_read_illegal_T_261 | _io_decode_0_read_illegal_T_116; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_263 = _io_decode_0_read_illegal_T_262 | _io_decode_0_read_illegal_T_117; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_264 = _io_decode_0_read_illegal_T_263 | _io_decode_0_read_illegal_T_118; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_265 = _io_decode_0_read_illegal_T_264 | _io_decode_0_read_illegal_T_119; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_266 = _io_decode_0_read_illegal_T_265 | _io_decode_0_read_illegal_T_120; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_267 = _io_decode_0_read_illegal_T_266 | _io_decode_0_read_illegal_T_121; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_268 = _io_decode_0_read_illegal_T_267 | _io_decode_0_read_illegal_T_122; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_269 = _io_decode_0_read_illegal_T_268 | _io_decode_0_read_illegal_T_123; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_270 = _io_decode_0_read_illegal_T_269 | _io_decode_0_read_illegal_T_124; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_271 = _io_decode_0_read_illegal_T_270 | _io_decode_0_read_illegal_T_125; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_272 = _io_decode_0_read_illegal_T_271 | _io_decode_0_read_illegal_T_126; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_273 = _io_decode_0_read_illegal_T_272 | _io_decode_0_read_illegal_T_127; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_274 = _io_decode_0_read_illegal_T_273 | _io_decode_0_read_illegal_T_128; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_275 = _io_decode_0_read_illegal_T_274 | _io_decode_0_read_illegal_T_129; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_276 = _io_decode_0_read_illegal_T_275 | _io_decode_0_read_illegal_T_130; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_277 = _io_decode_0_read_illegal_T_276 | _io_decode_0_read_illegal_T_131; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_278 = _io_decode_0_read_illegal_T_277 | _io_decode_0_read_illegal_T_132; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_279 = _io_decode_0_read_illegal_T_278 | _io_decode_0_read_illegal_T_133; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_280 = _io_decode_0_read_illegal_T_279 | _io_decode_0_read_illegal_T_134; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_281 = _io_decode_0_read_illegal_T_280 | _io_decode_0_read_illegal_T_135; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_282 = _io_decode_0_read_illegal_T_281 | _io_decode_0_read_illegal_T_136; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_283 = _io_decode_0_read_illegal_T_282 | _io_decode_0_read_illegal_T_137; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_284 = _io_decode_0_read_illegal_T_283 | _io_decode_0_read_illegal_T_138; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_285 = _io_decode_0_read_illegal_T_284 | _io_decode_0_read_illegal_T_139; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_286 = _io_decode_0_read_illegal_T_285 | _io_decode_0_read_illegal_T_140; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_287 = _io_decode_0_read_illegal_T_286 | _io_decode_0_read_illegal_T_141; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_288 = _io_decode_0_read_illegal_T_287 | _io_decode_0_read_illegal_T_142; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_289 = _io_decode_0_read_illegal_T_288 | _io_decode_0_read_illegal_T_143; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_290 = _io_decode_0_read_illegal_T_289 | _io_decode_0_read_illegal_T_144; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_291 = _io_decode_0_read_illegal_T_290 | _io_decode_0_read_illegal_T_145; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_292 = _io_decode_0_read_illegal_T_291 | _io_decode_0_read_illegal_T_146; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_293 = _io_decode_0_read_illegal_T_292 | _io_decode_0_read_illegal_T_147; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_294 = _io_decode_0_read_illegal_T_293 | _io_decode_0_read_illegal_T_148; // @[CSR.scala 655:115]
  assign _io_decode_0_read_illegal_T_296 = _io_decode_0_read_illegal_T_1 | ~_io_decode_0_read_illegal_T_294; // @[CSR.scala 671:62]
  assign _io_decode_0_read_illegal_T_299 = _io_decode_0_read_illegal_T_121 & ~allow_sfence_vma; // @[CSR.scala 673:32]
  assign _io_decode_0_read_illegal_T_300 = _io_decode_0_read_illegal_T_296 | _io_decode_0_read_illegal_T_299; // @[CSR.scala 672:32]
  assign _io_decode_0_read_illegal_T_301 = io_decode_0_csr >= 12'hc00; // @[package.scala 204:47]
  assign _io_decode_0_read_illegal_T_302 = io_decode_0_csr < 12'hc20; // @[package.scala 204:60]
  assign _io_decode_0_read_illegal_T_303 = _io_decode_0_read_illegal_T_301 & _io_decode_0_read_illegal_T_302; // @[package.scala 204:55]
  assign _io_decode_0_read_illegal_T_304 = io_decode_0_csr >= 12'hc80; // @[package.scala 204:47]
  assign _io_decode_0_read_illegal_T_305 = io_decode_0_csr < 12'hca0; // @[package.scala 204:60]
  assign _io_decode_0_read_illegal_T_306 = _io_decode_0_read_illegal_T_304 & _io_decode_0_read_illegal_T_305; // @[package.scala 204:55]
  assign _io_decode_0_read_illegal_T_307 = _io_decode_0_read_illegal_T_303 | _io_decode_0_read_illegal_T_306; // @[CSR.scala 674:66]
  assign _io_decode_0_read_illegal_T_309 = _io_decode_0_read_illegal_T_307 & ~allow_counter; // @[CSR.scala 674:130]
  assign _io_decode_0_read_illegal_T_310 = _io_decode_0_read_illegal_T_300 | _io_decode_0_read_illegal_T_309; // @[CSR.scala 673:53]
  assign _io_decode_0_read_illegal_T_311 = io_decode_0_csr & 12'hc10; // @[Decode.scala 14:65]
  assign _io_decode_0_read_illegal_T_312 = _io_decode_0_read_illegal_T_311 == 12'h410; // @[Decode.scala 14:121]
  assign _io_decode_0_read_illegal_T_316 = _io_decode_0_read_illegal_T_312 & ~reg_debug; // @[CSR.scala 675:42]
  assign _io_decode_0_read_illegal_T_317 = _io_decode_0_read_illegal_T_310 | _io_decode_0_read_illegal_T_316; // @[CSR.scala 674:148]
  assign _io_decode_0_read_illegal_T_320 = io_decode_0_fp_csr & io_decode_0_fp_illegal; // @[CSR.scala 677:21]
  assign _io_decode_0_write_flush_T = io_decode_0_csr >= 12'h340; // @[CSR.scala 679:40]
  assign _io_decode_0_write_flush_T_1 = io_decode_0_csr <= 12'h343; // @[CSR.scala 679:71]
  assign _io_decode_0_write_flush_T_2 = _io_decode_0_write_flush_T & _io_decode_0_write_flush_T_1; // @[CSR.scala 679:57]
  assign _io_decode_0_write_flush_T_3 = io_decode_0_csr >= 12'h140; // @[CSR.scala 679:99]
  assign _io_decode_0_write_flush_T_4 = io_decode_0_csr <= 12'h143; // @[CSR.scala 679:130]
  assign _io_decode_0_write_flush_T_5 = _io_decode_0_write_flush_T_3 & _io_decode_0_write_flush_T_4; // @[CSR.scala 679:116]
  assign _io_decode_0_write_flush_T_6 = _io_decode_0_write_flush_T_2 | _io_decode_0_write_flush_T_5; // @[CSR.scala 679:85]
  assign _io_decode_0_system_illegal_T_3 = is_wfi & ~allow_wfi; // @[CSR.scala 681:14]
  assign _io_decode_0_system_illegal_T_4 = _io_decode_0_read_illegal_T_1 | _io_decode_0_system_illegal_T_3; // @[CSR.scala 680:64]
  assign _io_decode_0_system_illegal_T_6 = is_ret & ~allow_sret; // @[CSR.scala 682:14]
  assign _io_decode_0_system_illegal_T_7 = _io_decode_0_system_illegal_T_4 | _io_decode_0_system_illegal_T_6; // @[CSR.scala 681:28]
  assign _io_decode_0_system_illegal_T_9 = is_ret & io_decode_0_csr[10]; // @[CSR.scala 683:14]
  assign _io_decode_0_system_illegal_T_11 = _io_decode_0_system_illegal_T_9 & io_decode_0_csr[7]; // @[CSR.scala 683:32]
  assign _io_decode_0_system_illegal_T_13 = _io_decode_0_system_illegal_T_11 & ~reg_debug; // @[CSR.scala 683:49]
  assign _io_decode_0_system_illegal_T_14 = _io_decode_0_system_illegal_T_7 | _io_decode_0_system_illegal_T_13; // @[CSR.scala 682:29]
  assign _io_decode_0_system_illegal_T_16 = is_sfence & ~allow_sfence_vma; // @[CSR.scala 684:17]
  assign _debugTVec_T = insn_break ? 12'h800 : 12'h808; // @[CSR.scala 697:37]
  assign debugTVec = reg_debug ? _debugTVec_T : 12'h800; // @[CSR.scala 697:22]
  assign notDebugTVec_base = delegate ? read_stvec : read_mtvec; // @[CSR.scala 705:19]
  assign notDebugTVec_interruptVec_lo = {cause[5:0], 2'h0}; // @[CSR.scala 706:59]
  assign notDebugTVec_interruptVec_hi = notDebugTVec_base[63:8]; // @[CSR.scala 707:33]
  assign notDebugTVec_interruptVec = {notDebugTVec_interruptVec_hi,notDebugTVec_interruptVec_lo}; // @[Cat.scala 30:58]
  assign _notDebugTVec_doVector_T_2 = notDebugTVec_base[0] & cause[63]; // @[CSR.scala 708:28]
  assign _notDebugTVec_doVector_T_4 = cause_lsbs[7:6] == 2'h0; // @[CSR.scala 708:94]
  assign notDebugTVec_doVector = _notDebugTVec_doVector_T_2 & _notDebugTVec_doVector_T_4; // @[CSR.scala 708:55]
  assign _notDebugTVec_T_1 = {notDebugTVec_base[63:2], 2'h0}; // @[CSR.scala 709:56]
  assign notDebugTVec = notDebugTVec_doVector ? notDebugTVec_interruptVec : _notDebugTVec_T_1; // @[CSR.scala 709:8]
  assign tvec = trapToDebug ? {{52'd0}, debugTVec} : notDebugTVec; // @[CSR.scala 723:17]
  assign _io_status_sd_T = &io_status_fs; // @[CSR.scala 729:32]
  assign _io_status_sd_T_1 = &io_status_xs; // @[CSR.scala 729:53]
  assign _io_status_sd_T_2 = _io_status_sd_T | _io_status_sd_T_1; // @[CSR.scala 729:37]
  assign _io_status_sd_T_3 = &io_status_vs; // @[CSR.scala 729:74]
  assign _io_status_dprv_x87_T_1 = reg_mstatus_mprv & ~reg_debug; // @[CSR.scala 734:53]
  assign _T_244 = insn_ret + insn_call; // @[Bitwise.scala 47:55]
  assign _T_246 = insn_break + io_exception; // @[Bitwise.scala 47:55]
  assign _T_248 = _T_244 + _T_246; // @[Bitwise.scala 47:55]
  assign _T_250 = _T_248 <= 3'h1; // @[CSR.scala 739:79]
  assign _T_252 = _T_250 | reset; // @[CSR.scala 739:9]
  assign _T_255 = insn_wfi & ~io_singleStep; // @[CSR.scala 741:18]
  assign _T_257 = _T_255 & ~reg_debug; // @[CSR.scala 741:36]
  assign _GEN_48 = _T_257 | reg_wfi; // @[CSR.scala 741:51]
  assign _T_258 = |pending_interrupts; // @[CSR.scala 742:28]
  assign _T_259 = _T_258 | io_interrupts_debug; // @[CSR.scala 742:32]
  assign _T_260 = _T_259 | exception; // @[CSR.scala 742:55]
  assign _T_262 = io_retire | exception; // @[CSR.scala 745:22]
  assign _GEN_50 = _T_262 | reg_singleStepped; // @[CSR.scala 745:36]
  assign _T_272 = ~reg_singleStepped | ~io_retire; // @[CSR.scala 748:29]
  assign _T_274 = _T_272 | reset; // @[CSR.scala 748:9]
  assign _epc_T_1 = ~io_pc | 40'h1; // @[CSR.scala 1207:31]
  assign epc = ~_epc_T_1; // @[CSR.scala 1207:26]
  assign _reg_dcsr_cause_T = causeIsDebugTrigger ? 2'h2 : 2'h1; // @[CSR.scala 759:86]
  assign _reg_dcsr_cause_T_1 = causeIsDebugInt ? 2'h3 : _reg_dcsr_cause_T; // @[CSR.scala 759:56]
  assign _GEN_52 = ~reg_debug | reg_debug; // @[CSR.scala 756:25]
  assign _GEN_53 = reg_debug ? reg_dpc : epc; // @[CSR.scala 756:25]
  assign _GEN_63 = _T_279 ? epc : reg_sepc; // @[CSR.scala 772:35]
  assign _GEN_67 = _T_279 ? reg_mstatus_sie : reg_mstatus_spie; // @[CSR.scala 772:35]
  assign _GEN_68 = _T_279 ? reg_mstatus_prv : {{1'd0}, reg_mstatus_spp}; // @[CSR.scala 772:35]
  assign _GEN_71 = _T_279 ? reg_mepc : epc; // @[CSR.scala 772:35]
  assign _GEN_74 = _T_279 ? reg_mstatus_mpie : reg_mstatus_mie; // @[CSR.scala 772:35]
  assign _GEN_75 = _T_279 ? reg_mstatus_mpp : reg_mstatus_prv; // @[CSR.scala 772:35]
  assign _GEN_76 = _T_279 & reg_mstatus_mie; // @[CSR.scala 772:35]
  assign _GEN_97 = trapToDebug ? _GEN_53 : reg_dpc; // @[CSR.scala 755:24]
  assign _GEN_106 = trapToDebug ? reg_sepc : _GEN_63; // @[CSR.scala 755:24]
  assign _GEN_110 = trapToDebug ? reg_mstatus_spie : _GEN_67; // @[CSR.scala 755:24]
  assign _GEN_111 = trapToDebug ? {{1'd0}, reg_mstatus_spp} : _GEN_68; // @[CSR.scala 755:24]
  assign _GEN_113 = trapToDebug ? reg_mepc : _GEN_71; // @[CSR.scala 755:24]
  assign _GEN_116 = trapToDebug ? reg_mstatus_mpie : _GEN_74; // @[CSR.scala 755:24]
  assign _GEN_117 = trapToDebug ? reg_mstatus_mpp : _GEN_75; // @[CSR.scala 755:24]
  assign _GEN_118 = trapToDebug ? reg_mstatus_mie : _GEN_76; // @[CSR.scala 755:24]
  assign _GEN_120 = exception ? _GEN_97 : reg_dpc; // @[CSR.scala 754:20]
  assign _GEN_129 = exception ? _GEN_106 : reg_sepc; // @[CSR.scala 754:20]
  assign _GEN_133 = exception ? _GEN_110 : reg_mstatus_spie; // @[CSR.scala 754:20]
  assign _GEN_134 = exception ? _GEN_111 : {{1'd0}, reg_mstatus_spp}; // @[CSR.scala 754:20]
  assign _GEN_136 = exception ? _GEN_113 : reg_mepc; // @[CSR.scala 754:20]
  assign _GEN_139 = exception ? _GEN_116 : reg_mstatus_mpie; // @[CSR.scala 754:20]
  assign _GEN_140 = exception ? _GEN_117 : reg_mstatus_mpp; // @[CSR.scala 754:20]
  assign _GEN_141 = exception ? _GEN_118 : reg_mstatus_mie; // @[CSR.scala 754:20]
  assign _GEN_151 = _T_406 ? lo_6 : lo_4; // @[CSR.scala 821:70]
  assign _GEN_158 = ~io_rw_addr[9] | _GEN_133; // @[CSR.scala 815:52]
  assign _GEN_159 = io_rw_addr[9] ? _GEN_134 : 2'h0; // @[CSR.scala 815:52]
  assign _GEN_161 = io_rw_addr[9] ? _GEN_151 : lo_8; // @[CSR.scala 815:52]
  assign _T_412 = ret_prv < 2'h3; // @[CSR.scala 839:32]
  assign _GEN_171 = insn_ret ? _GEN_159 : _GEN_134; // @[CSR.scala 813:19]
  assign _GEN_172 = insn_ret ? {{24'd0}, _GEN_161} : tvec; // @[CSR.scala 813:19]
  assign _GEN_181 = insn_cease | io_status_cease_r; // @[Reg.scala 28:19]
  assign _io_rw_rdata_T_1 = _T_46 ? _T_7 : 64'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_2 = _T_47 ? _T_10 : 64'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_4 = _T_49 ? reg_misa : 64'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_5 = _T_50 ? read_mstatus : 64'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_6 = _T_51 ? read_mtvec : 64'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_7 = _T_52 ? read_mip : 16'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_8 = _T_53 ? reg_mie : 64'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_9 = _T_54 ? reg_mscratch : 64'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_10 = _T_55 ? _T_18 : 64'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_11 = _T_56 ? _T_21 : 64'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_12 = _T_57 ? reg_mcause : 64'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_13 = _T_58 & io_hartid; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_14 = _T_59 ? _T_22 : 32'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_15 = _T_60 ? _T_29 : 64'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_16 = _T_61 ? reg_dscratch : 64'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_17 = _T_62 ? reg_fflags : 5'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_18 = _T_63 ? reg_frm : 3'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_19 = _T_64 ? read_fcsr : 8'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_20 = _T_65 ? reg_mcountinhibit : 3'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_21 = _T_66 ? value_1 : 64'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_22 = _T_67 ? value : 64'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_110 = _T_155 ? read_mcounteren : 32'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_111 = _T_156 ? value_1 : 64'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_112 = _T_157 ? value : 64'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_113 = _T_158 ? _T_30[63:0] : 64'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_114 = _T_159 ? read_sip : 64'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_115 = _T_160 ? read_sie : 64'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_116 = _T_161 ? reg_sscratch : 64'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_117 = _T_162 ? reg_scause : 64'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_118 = _T_163 ? _T_34 : 64'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_119 = _T_164 ? _T_35 : 64'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_120 = _T_165 ? _T_42 : 64'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_121 = _T_166 ? read_stvec : 64'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_122 = _T_167 ? read_scounteren : 32'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_123 = _T_168 ? read_mideleg : 64'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_124 = _T_169 ? read_medeleg : 64'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_125 = _T_170 ? _T_43 : 64'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_127 = _T_172 ? reg_pmp_0_addr : 30'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_128 = _T_173 ? reg_pmp_1_addr : 30'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_129 = _T_174 ? reg_pmp_2_addr : 30'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_130 = _T_175 ? reg_pmp_3_addr : 30'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_131 = _T_176 ? reg_pmp_4_addr : 30'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_132 = _T_177 ? reg_pmp_5_addr : 30'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_133 = _T_178 ? reg_pmp_6_addr : 30'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_134 = _T_179 ? reg_pmp_7_addr : 30'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_143 = _T_188 ? reg_custom_0 : 64'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_144 = _T_189 ? 64'h1 : 64'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_146 = _T_191 ? 64'h20181004 : 64'h0; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_148 = _io_rw_rdata_T_1 | _io_rw_rdata_T_2; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_150 = _io_rw_rdata_T_148 | _io_rw_rdata_T_4; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_151 = _io_rw_rdata_T_150 | _io_rw_rdata_T_5; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_152 = _io_rw_rdata_T_151 | _io_rw_rdata_T_6; // @[Mux.scala 27:72]
  assign _GEN_565 = {{48'd0}, _io_rw_rdata_T_7}; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_153 = _io_rw_rdata_T_152 | _GEN_565; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_154 = _io_rw_rdata_T_153 | _io_rw_rdata_T_8; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_155 = _io_rw_rdata_T_154 | _io_rw_rdata_T_9; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_156 = _io_rw_rdata_T_155 | _io_rw_rdata_T_10; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_157 = _io_rw_rdata_T_156 | _io_rw_rdata_T_11; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_158 = _io_rw_rdata_T_157 | _io_rw_rdata_T_12; // @[Mux.scala 27:72]
  assign _GEN_566 = {{63'd0}, _io_rw_rdata_T_13}; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_159 = _io_rw_rdata_T_158 | _GEN_566; // @[Mux.scala 27:72]
  assign _GEN_567 = {{32'd0}, _io_rw_rdata_T_14}; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_160 = _io_rw_rdata_T_159 | _GEN_567; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_161 = _io_rw_rdata_T_160 | _io_rw_rdata_T_15; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_162 = _io_rw_rdata_T_161 | _io_rw_rdata_T_16; // @[Mux.scala 27:72]
  assign _GEN_568 = {{59'd0}, _io_rw_rdata_T_17}; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_163 = _io_rw_rdata_T_162 | _GEN_568; // @[Mux.scala 27:72]
  assign _GEN_569 = {{61'd0}, _io_rw_rdata_T_18}; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_164 = _io_rw_rdata_T_163 | _GEN_569; // @[Mux.scala 27:72]
  assign _GEN_570 = {{56'd0}, _io_rw_rdata_T_19}; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_165 = _io_rw_rdata_T_164 | _GEN_570; // @[Mux.scala 27:72]
  assign _GEN_571 = {{61'd0}, _io_rw_rdata_T_20}; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_166 = _io_rw_rdata_T_165 | _GEN_571; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_167 = _io_rw_rdata_T_166 | _io_rw_rdata_T_21; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_168 = _io_rw_rdata_T_167 | _io_rw_rdata_T_22; // @[Mux.scala 27:72]
  assign _GEN_572 = {{32'd0}, _io_rw_rdata_T_110}; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_256 = _io_rw_rdata_T_168 | _GEN_572; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_257 = _io_rw_rdata_T_256 | _io_rw_rdata_T_111; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_258 = _io_rw_rdata_T_257 | _io_rw_rdata_T_112; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_259 = _io_rw_rdata_T_258 | _io_rw_rdata_T_113; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_260 = _io_rw_rdata_T_259 | _io_rw_rdata_T_114; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_261 = _io_rw_rdata_T_260 | _io_rw_rdata_T_115; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_262 = _io_rw_rdata_T_261 | _io_rw_rdata_T_116; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_263 = _io_rw_rdata_T_262 | _io_rw_rdata_T_117; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_264 = _io_rw_rdata_T_263 | _io_rw_rdata_T_118; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_265 = _io_rw_rdata_T_264 | _io_rw_rdata_T_119; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_266 = _io_rw_rdata_T_265 | _io_rw_rdata_T_120; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_267 = _io_rw_rdata_T_266 | _io_rw_rdata_T_121; // @[Mux.scala 27:72]
  assign _GEN_573 = {{32'd0}, _io_rw_rdata_T_122}; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_268 = _io_rw_rdata_T_267 | _GEN_573; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_269 = _io_rw_rdata_T_268 | _io_rw_rdata_T_123; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_270 = _io_rw_rdata_T_269 | _io_rw_rdata_T_124; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_271 = _io_rw_rdata_T_270 | _io_rw_rdata_T_125; // @[Mux.scala 27:72]
  assign _GEN_574 = {{34'd0}, _io_rw_rdata_T_127}; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_273 = _io_rw_rdata_T_271 | _GEN_574; // @[Mux.scala 27:72]
  assign _GEN_575 = {{34'd0}, _io_rw_rdata_T_128}; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_274 = _io_rw_rdata_T_273 | _GEN_575; // @[Mux.scala 27:72]
  assign _GEN_576 = {{34'd0}, _io_rw_rdata_T_129}; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_275 = _io_rw_rdata_T_274 | _GEN_576; // @[Mux.scala 27:72]
  assign _GEN_577 = {{34'd0}, _io_rw_rdata_T_130}; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_276 = _io_rw_rdata_T_275 | _GEN_577; // @[Mux.scala 27:72]
  assign _GEN_578 = {{34'd0}, _io_rw_rdata_T_131}; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_277 = _io_rw_rdata_T_276 | _GEN_578; // @[Mux.scala 27:72]
  assign _GEN_579 = {{34'd0}, _io_rw_rdata_T_132}; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_278 = _io_rw_rdata_T_277 | _GEN_579; // @[Mux.scala 27:72]
  assign _GEN_580 = {{34'd0}, _io_rw_rdata_T_133}; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_279 = _io_rw_rdata_T_278 | _GEN_580; // @[Mux.scala 27:72]
  assign _GEN_581 = {{34'd0}, _io_rw_rdata_T_134}; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_280 = _io_rw_rdata_T_279 | _GEN_581; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_289 = _io_rw_rdata_T_280 | _io_rw_rdata_T_143; // @[Mux.scala 27:72]
  assign _io_rw_rdata_T_290 = _io_rw_rdata_T_289 | _io_rw_rdata_T_144; // @[Mux.scala 27:72]
  assign _T_416 = io_rw_cmd == 3'h5; // @[package.scala 15:47]
  assign _T_417 = io_rw_cmd == 3'h6; // @[package.scala 15:47]
  assign _T_418 = io_rw_cmd == 3'h7; // @[package.scala 15:47]
  assign _lo_T = reg_fflags | io_fcsr_flags_bits; // @[CSR.scala 887:30]
  assign _GEN_182 = io_fcsr_flags_valid ? _lo_T : reg_fflags; // @[CSR.scala 886:30]
  assign _csr_wen_T_3 = _T_417 | _T_418; // @[package.scala 72:59]
  assign csr_wen = _csr_wen_T_3 | _T_416; // @[package.scala 72:59]
  assign _new_mstatus_WIRE = {{39'd0}, wdata};
  assign new_mstatus_sie = _new_mstatus_WIRE[1]; // @[CSR.scala 902:47]
  assign new_mstatus_mie = _new_mstatus_WIRE[3]; // @[CSR.scala 902:47]
  assign new_mstatus_spie = _new_mstatus_WIRE[5]; // @[CSR.scala 902:47]
  assign new_mstatus_mpie = _new_mstatus_WIRE[7]; // @[CSR.scala 902:47]
  assign new_mstatus_spp = _new_mstatus_WIRE[8]; // @[CSR.scala 902:47]
  assign new_mstatus_mpp = _new_mstatus_WIRE[12:11]; // @[CSR.scala 902:47]
  assign new_mstatus_fs = _new_mstatus_WIRE[14:13]; // @[CSR.scala 902:47]
  assign new_mstatus_mprv = _new_mstatus_WIRE[17]; // @[CSR.scala 902:47]
  assign new_mstatus_sum = _new_mstatus_WIRE[18]; // @[CSR.scala 902:47]
  assign new_mstatus_mxr = _new_mstatus_WIRE[19]; // @[CSR.scala 902:47]
  assign new_mstatus_tvm = _new_mstatus_WIRE[20]; // @[CSR.scala 902:47]
  assign new_mstatus_tw = _new_mstatus_WIRE[21]; // @[CSR.scala 902:47]
  assign new_mstatus_tsr = _new_mstatus_WIRE[22]; // @[CSR.scala 902:47]
  assign _reg_mstatus_mpp_T_2 = new_mstatus_mpp == 2'h2; // @[CSR.scala 1190:35]
  assign _reg_mstatus_fs_T = |new_mstatus_fs; // @[CSR.scala 1211:73]
  assign _GEN_188 = _T_50 ? {{1'd0}, new_mstatus_spp} : _GEN_171; // @[CSR.scala 901:39]
  assign f = wdata[5]; // @[CSR.scala 928:20]
  assign _T_1834 = ~io_pc[1] | wdata[2]; // @[CSR.scala 930:43]
  assign _reg_misa_T_2 = {~f, 3'h0}; // @[CSR.scala 932:38]
  assign _GEN_582 = {{60'd0}, _reg_misa_T_2}; // @[CSR.scala 932:32]
  assign _reg_misa_T_3 = ~wdata | _GEN_582; // @[CSR.scala 932:32]
  assign _reg_misa_T_5 = ~_reg_misa_T_3 & 64'h102d; // @[CSR.scala 932:55]
  assign _reg_misa_T_7 = reg_misa & 64'hffffffffffffefd2; // @[CSR.scala 932:73]
  assign _reg_misa_T_8 = _reg_misa_T_5 | _reg_misa_T_7; // @[CSR.scala 932:62]
  assign _new_mip_T = {4'h0,2'h0,reg_mip_seip,1'h0,2'h0,reg_mip_stip,1'h0,2'h0,reg_mip_ssip,1'h0}; // @[CSR.scala 940:59]
  assign _new_mip_T_2 = io_rw_cmd[1] ? _new_mip_T : 16'h0; // @[CSR.scala 1186:9]
  assign _GEN_583 = {{48'd0}, _new_mip_T_2}; // @[CSR.scala 1186:34]
  assign _new_mip_T_3 = _GEN_583 | io_rw_wdata; // @[CSR.scala 1186:34]
  assign _new_mip_T_8 = _new_mip_T_3 & ~_wdata_T_5; // @[CSR.scala 1186:43]
  assign new_mip_ssip = _new_mip_T_8[1]; // @[CSR.scala 940:88]
  assign new_mip_stip = _new_mip_T_8[5]; // @[CSR.scala 940:88]
  assign new_mip_seip = _new_mip_T_8[9]; // @[CSR.scala 940:88]
  assign _reg_mie_T = wdata & 64'haaa; // @[CSR.scala 947:59]
  assign _reg_mepc_T_1 = ~wdata | 64'h1; // @[CSR.scala 1207:31]
  assign _GEN_204 = _T_55 ? ~_reg_mepc_T_1 : {{24'd0}, _GEN_136}; // @[CSR.scala 948:40]
  assign _GEN_206 = _T_51 ? wdata : {{32'd0}, reg_mtvec}; // @[CSR.scala 951:40]
  assign _reg_mcause_T = wdata & 64'h800000000000000f; // @[CSR.scala 952:62]
  assign _reg_mcountinhibit_T_1 = wdata & 64'hfffffffffffffffd; // @[CSR.scala 968:76]
  assign _GEN_209 = _T_65 ? _reg_mcountinhibit_T_1 : {{61'd0}, reg_mcountinhibit}; // @[CSR.scala 968:47]
  assign _GEN_210 = _T_66 ? wdata : {{57'd0}, _GEN_2}; // @[CSR.scala 1204:31]
  assign _GEN_212 = _T_67 ? wdata : {{57'd0}, _GEN_0}; // @[CSR.scala 1204:31]
  assign _GEN_215 = _T_62 ? wdata : {{59'd0}, _GEN_182}; // @[CSR.scala 974:40]
  assign _GEN_217 = _T_63 ? wdata : {{61'd0}, reg_frm}; // @[CSR.scala 975:40]
  assign _GEN_219 = _T_64 ? wdata : _GEN_215; // @[CSR.scala 976:38]
  assign _GEN_220 = _T_64 ? {{5'd0}, wdata[63:5]} : _GEN_217; // @[CSR.scala 976:38]
  assign new_dcsr_prv = wdata[1:0]; // @[CSR.scala 984:43]
  assign new_dcsr_step = wdata[2]; // @[CSR.scala 984:43]
  assign new_dcsr_ebreaku = wdata[12]; // @[CSR.scala 984:43]
  assign new_dcsr_ebreaks = wdata[13]; // @[CSR.scala 984:43]
  assign new_dcsr_ebreakm = wdata[15]; // @[CSR.scala 984:43]
  assign _reg_dcsr_prv_T = new_dcsr_prv == 2'h2; // @[CSR.scala 1190:35]
  assign _GEN_226 = _T_60 ? ~_reg_mepc_T_1 : {{24'd0}, _GEN_120}; // @[CSR.scala 991:42]
  assign _GEN_230 = _T_158 ? {{1'd0}, new_mstatus_spp} : _GEN_188; // @[CSR.scala 998:41]
  assign _new_sip_T_1 = _GEN_45 & ~read_mideleg; // @[CSR.scala 1011:52]
  assign _new_sip_T_2 = wdata & read_mideleg; // @[CSR.scala 1011:78]
  assign _new_sip_T_3 = _new_sip_T_1 | _new_sip_T_2; // @[CSR.scala 1011:69]
  assign new_sip_ssip = _new_sip_T_3[1]; // @[CSR.scala 1011:41]
  assign new_satp_ppn = wdata[43:0]; // @[CSR.scala 1016:45]
  assign new_satp_mode = wdata[63:60]; // @[CSR.scala 1016:45]
  assign _T_1837 = new_satp_mode == 4'h0; // @[package.scala 15:47]
  assign _T_1838 = new_satp_mode == 4'h8; // @[package.scala 15:47]
  assign _T_1839 = _T_1837 | _T_1838; // @[package.scala 72:59]
  assign _reg_satp_mode_T = new_satp_mode & 4'h8; // @[CSR.scala 1019:44]
  assign _reg_mie_T_2 = reg_mie & ~read_mideleg; // @[CSR.scala 1025:64]
  assign _reg_mie_T_4 = _reg_mie_T_2 | _new_sip_T_2; // @[CSR.scala 1025:81]
  assign _GEN_242 = _T_165 ? ~_reg_mepc_T_1 : {{24'd0}, _GEN_129}; // @[CSR.scala 1027:42]
  assign _GEN_243 = _T_166 ? wdata : {{25'd0}, reg_stvec}; // @[CSR.scala 1028:42]
  assign _reg_scause_T = wdata & 64'h800000000000001f; // @[CSR.scala 1029:64]
  assign _GEN_248 = _T_167 ? wdata : {{32'd0}, reg_scounteren}; // @[CSR.scala 1033:44]
  assign _GEN_249 = _T_155 ? wdata : {{32'd0}, reg_mcounteren}; // @[CSR.scala 1036:44]
  assign _T_1842 = ~reg_bp_0_control_dmode | reg_debug; // @[CSR.scala 1042:55]
  assign _GEN_251 = _T_47 ? wdata : {{25'd0}, reg_bp_0_address}; // @[CSR.scala 1043:44]
  assign _newBPC_T_2 = io_rw_cmd[1] ? _T_7 : 64'h0; // @[CSR.scala 1186:9]
  assign _newBPC_T_3 = _newBPC_T_2 | io_rw_wdata; // @[CSR.scala 1186:34]
  assign _newBPC_T_8 = _newBPC_T_3 & ~_wdata_T_5; // @[CSR.scala 1186:43]
  assign newBPC_action = _newBPC_T_8[12]; // @[CSR.scala 1061:96]
  assign newBPC_dmode = _newBPC_T_8[59]; // @[CSR.scala 1061:96]
  assign dMode = newBPC_dmode & reg_debug; // @[CSR.scala 1062:38]
  assign _GEN_252 = dMode & newBPC_action; // @[CSR.scala 1064:51]
  assign _GEN_268 = _T_1842 ? _GEN_251 : {{25'd0}, reg_bp_0_address}; // @[CSR.scala 1042:70]
  assign _T_1853 = _T_170 & ~reg_pmp_0_cfg_l; // @[CSR.scala 1074:57]
  assign newCfg_r = wdata[0]; // @[CSR.scala 1075:46]
  assign newCfg_w = wdata[1]; // @[CSR.scala 1075:46]
  assign newCfg_x = wdata[2]; // @[CSR.scala 1075:46]
  assign newCfg_a = wdata[4:3]; // @[CSR.scala 1075:46]
  assign newCfg_l = wdata[7]; // @[CSR.scala 1075:46]
  assign _reg_pmp_0_cfg_w_T = newCfg_w & newCfg_r; // @[CSR.scala 1078:31]
  assign _T_1857 = ~reg_pmp_1_cfg_a[1] & pmp_mask_base_lo_1; // @[PMP.scala 49:20]
  assign _T_1858 = reg_pmp_1_cfg_l & _T_1857; // @[PMP.scala 51:62]
  assign _T_1859 = reg_pmp_0_cfg_l | _T_1858; // @[PMP.scala 51:44]
  assign _T_1861 = _T_172 & ~_T_1859; // @[CSR.scala 1083:45]
  assign _GEN_323 = _T_1861 ? wdata : {{34'd0}, reg_pmp_0_addr}; // @[CSR.scala 1083:71]
  assign _T_1863 = _T_170 & ~reg_pmp_1_cfg_l; // @[CSR.scala 1074:57]
  assign newCfg_1_r = wdata[8]; // @[CSR.scala 1075:46]
  assign newCfg_1_w = wdata[9]; // @[CSR.scala 1075:46]
  assign newCfg_1_x = wdata[10]; // @[CSR.scala 1075:46]
  assign newCfg_1_a = wdata[12:11]; // @[CSR.scala 1075:46]
  assign newCfg_1_l = wdata[15]; // @[CSR.scala 1075:46]
  assign _reg_pmp_1_cfg_w_T = newCfg_1_w & newCfg_1_r; // @[CSR.scala 1078:31]
  assign _T_1867 = ~reg_pmp_2_cfg_a[1] & pmp_mask_base_lo_2; // @[PMP.scala 49:20]
  assign _T_1868 = reg_pmp_2_cfg_l & _T_1867; // @[PMP.scala 51:62]
  assign _T_1869 = reg_pmp_1_cfg_l | _T_1868; // @[PMP.scala 51:44]
  assign _T_1871 = _T_173 & ~_T_1869; // @[CSR.scala 1083:45]
  assign _GEN_330 = _T_1871 ? wdata : {{34'd0}, reg_pmp_1_addr}; // @[CSR.scala 1083:71]
  assign _T_1873 = _T_170 & ~reg_pmp_2_cfg_l; // @[CSR.scala 1074:57]
  assign newCfg_2_r = wdata[16]; // @[CSR.scala 1075:46]
  assign newCfg_2_w = wdata[17]; // @[CSR.scala 1075:46]
  assign newCfg_2_x = wdata[18]; // @[CSR.scala 1075:46]
  assign newCfg_2_a = wdata[20:19]; // @[CSR.scala 1075:46]
  assign newCfg_2_l = wdata[23]; // @[CSR.scala 1075:46]
  assign _reg_pmp_2_cfg_w_T = newCfg_2_w & newCfg_2_r; // @[CSR.scala 1078:31]
  assign _T_1877 = ~reg_pmp_3_cfg_a[1] & pmp_mask_base_lo_3; // @[PMP.scala 49:20]
  assign _T_1878 = reg_pmp_3_cfg_l & _T_1877; // @[PMP.scala 51:62]
  assign _T_1879 = reg_pmp_2_cfg_l | _T_1878; // @[PMP.scala 51:44]
  assign _T_1881 = _T_174 & ~_T_1879; // @[CSR.scala 1083:45]
  assign _GEN_337 = _T_1881 ? wdata : {{34'd0}, reg_pmp_2_addr}; // @[CSR.scala 1083:71]
  assign _T_1883 = _T_170 & ~reg_pmp_3_cfg_l; // @[CSR.scala 1074:57]
  assign newCfg_3_r = wdata[24]; // @[CSR.scala 1075:46]
  assign newCfg_3_w = wdata[25]; // @[CSR.scala 1075:46]
  assign newCfg_3_x = wdata[26]; // @[CSR.scala 1075:46]
  assign newCfg_3_a = wdata[28:27]; // @[CSR.scala 1075:46]
  assign newCfg_3_l = wdata[31]; // @[CSR.scala 1075:46]
  assign _reg_pmp_3_cfg_w_T = newCfg_3_w & newCfg_3_r; // @[CSR.scala 1078:31]
  assign _T_1887 = ~reg_pmp_4_cfg_a[1] & pmp_mask_base_lo_4; // @[PMP.scala 49:20]
  assign _T_1888 = reg_pmp_4_cfg_l & _T_1887; // @[PMP.scala 51:62]
  assign _T_1889 = reg_pmp_3_cfg_l | _T_1888; // @[PMP.scala 51:44]
  assign _T_1891 = _T_175 & ~_T_1889; // @[CSR.scala 1083:45]
  assign _GEN_344 = _T_1891 ? wdata : {{34'd0}, reg_pmp_3_addr}; // @[CSR.scala 1083:71]
  assign _T_1893 = _T_170 & ~reg_pmp_4_cfg_l; // @[CSR.scala 1074:57]
  assign newCfg_4_r = wdata[32]; // @[CSR.scala 1075:46]
  assign newCfg_4_w = wdata[33]; // @[CSR.scala 1075:46]
  assign newCfg_4_x = wdata[34]; // @[CSR.scala 1075:46]
  assign newCfg_4_a = wdata[36:35]; // @[CSR.scala 1075:46]
  assign newCfg_4_l = wdata[39]; // @[CSR.scala 1075:46]
  assign _reg_pmp_4_cfg_w_T = newCfg_4_w & newCfg_4_r; // @[CSR.scala 1078:31]
  assign _T_1897 = ~reg_pmp_5_cfg_a[1] & pmp_mask_base_lo_5; // @[PMP.scala 49:20]
  assign _T_1898 = reg_pmp_5_cfg_l & _T_1897; // @[PMP.scala 51:62]
  assign _T_1899 = reg_pmp_4_cfg_l | _T_1898; // @[PMP.scala 51:44]
  assign _T_1901 = _T_176 & ~_T_1899; // @[CSR.scala 1083:45]
  assign _GEN_351 = _T_1901 ? wdata : {{34'd0}, reg_pmp_4_addr}; // @[CSR.scala 1083:71]
  assign _T_1903 = _T_170 & ~reg_pmp_5_cfg_l; // @[CSR.scala 1074:57]
  assign newCfg_5_r = wdata[40]; // @[CSR.scala 1075:46]
  assign newCfg_5_w = wdata[41]; // @[CSR.scala 1075:46]
  assign newCfg_5_x = wdata[42]; // @[CSR.scala 1075:46]
  assign newCfg_5_a = wdata[44:43]; // @[CSR.scala 1075:46]
  assign newCfg_5_l = wdata[47]; // @[CSR.scala 1075:46]
  assign _reg_pmp_5_cfg_w_T = newCfg_5_w & newCfg_5_r; // @[CSR.scala 1078:31]
  assign _T_1907 = ~reg_pmp_6_cfg_a[1] & pmp_mask_base_lo_6; // @[PMP.scala 49:20]
  assign _T_1908 = reg_pmp_6_cfg_l & _T_1907; // @[PMP.scala 51:62]
  assign _T_1909 = reg_pmp_5_cfg_l | _T_1908; // @[PMP.scala 51:44]
  assign _T_1911 = _T_177 & ~_T_1909; // @[CSR.scala 1083:45]
  assign _GEN_358 = _T_1911 ? wdata : {{34'd0}, reg_pmp_5_addr}; // @[CSR.scala 1083:71]
  assign _T_1913 = _T_170 & ~reg_pmp_6_cfg_l; // @[CSR.scala 1074:57]
  assign newCfg_6_r = wdata[48]; // @[CSR.scala 1075:46]
  assign newCfg_6_w = wdata[49]; // @[CSR.scala 1075:46]
  assign newCfg_6_x = wdata[50]; // @[CSR.scala 1075:46]
  assign newCfg_6_a = wdata[52:51]; // @[CSR.scala 1075:46]
  assign newCfg_6_l = wdata[55]; // @[CSR.scala 1075:46]
  assign _reg_pmp_6_cfg_w_T = newCfg_6_w & newCfg_6_r; // @[CSR.scala 1078:31]
  assign _T_1917 = ~reg_pmp_7_cfg_a[1] & pmp_mask_base_lo_7; // @[PMP.scala 49:20]
  assign _T_1918 = reg_pmp_7_cfg_l & _T_1917; // @[PMP.scala 51:62]
  assign _T_1919 = reg_pmp_6_cfg_l | _T_1918; // @[PMP.scala 51:44]
  assign _T_1921 = _T_178 & ~_T_1919; // @[CSR.scala 1083:45]
  assign _GEN_365 = _T_1921 ? wdata : {{34'd0}, reg_pmp_6_addr}; // @[CSR.scala 1083:71]
  assign _T_1923 = _T_170 & ~reg_pmp_7_cfg_l; // @[CSR.scala 1074:57]
  assign newCfg_7_r = wdata[56]; // @[CSR.scala 1075:46]
  assign newCfg_7_w = wdata[57]; // @[CSR.scala 1075:46]
  assign newCfg_7_x = wdata[58]; // @[CSR.scala 1075:46]
  assign newCfg_7_a = wdata[60:59]; // @[CSR.scala 1075:46]
  assign newCfg_7_l = wdata[63]; // @[CSR.scala 1075:46]
  assign _reg_pmp_7_cfg_w_T = newCfg_7_w & newCfg_7_r; // @[CSR.scala 1078:31]
  assign _T_1929 = reg_pmp_7_cfg_l | _T_1918; // @[PMP.scala 51:44]
  assign _T_1931 = _T_179 & ~_T_1929; // @[CSR.scala 1083:45]
  assign _GEN_372 = _T_1931 ? wdata : {{34'd0}, reg_pmp_7_addr}; // @[CSR.scala 1083:71]
  assign _reg_custom_0_T = wdata & 64'h208; // @[CSR.scala 1090:23]
  assign _reg_custom_0_T_2 = reg_custom_0 & 64'hfffffffffffffdf7; // @[CSR.scala 1090:38]
  assign _reg_custom_0_T_3 = _reg_custom_0_T | _reg_custom_0_T_2; // @[CSR.scala 1090:31]
  assign _GEN_385 = csr_wen ? _GEN_230 : _GEN_171; // @[CSR.scala 900:18]
  assign _GEN_400 = csr_wen ? _GEN_204 : {{24'd0}, _GEN_136}; // @[CSR.scala 900:18]
  assign _GEN_402 = csr_wen ? _GEN_206 : {{32'd0}, reg_mtvec}; // @[CSR.scala 900:18]
  assign _GEN_405 = csr_wen ? _GEN_209 : {{61'd0}, reg_mcountinhibit}; // @[CSR.scala 900:18]
  assign _GEN_406 = csr_wen ? _GEN_210 : {{57'd0}, _GEN_2}; // @[CSR.scala 900:18]
  assign _GEN_408 = csr_wen ? _GEN_212 : {{57'd0}, _GEN_0}; // @[CSR.scala 900:18]
  assign _GEN_411 = csr_wen ? _GEN_219 : {{59'd0}, _GEN_182}; // @[CSR.scala 900:18]
  assign _GEN_412 = csr_wen ? _GEN_220 : {{61'd0}, reg_frm}; // @[CSR.scala 900:18]
  assign _GEN_418 = csr_wen ? _GEN_226 : {{24'd0}, _GEN_120}; // @[CSR.scala 900:18]
  assign _GEN_423 = csr_wen ? _GEN_242 : {{24'd0}, _GEN_129}; // @[CSR.scala 900:18]
  assign _GEN_424 = csr_wen ? _GEN_243 : {{25'd0}, reg_stvec}; // @[CSR.scala 900:18]
  assign _GEN_429 = csr_wen ? _GEN_248 : {{32'd0}, reg_scounteren}; // @[CSR.scala 900:18]
  assign _GEN_430 = csr_wen ? _GEN_249 : {{32'd0}, reg_mcounteren}; // @[CSR.scala 900:18]
  assign _GEN_432 = csr_wen ? _GEN_268 : {{25'd0}, reg_bp_0_address}; // @[CSR.scala 900:18]
  assign _GEN_470 = csr_wen ? _GEN_323 : {{34'd0}, reg_pmp_0_addr}; // @[CSR.scala 900:18]
  assign _GEN_477 = csr_wen ? _GEN_330 : {{34'd0}, reg_pmp_1_addr}; // @[CSR.scala 900:18]
  assign _GEN_484 = csr_wen ? _GEN_337 : {{34'd0}, reg_pmp_2_addr}; // @[CSR.scala 900:18]
  assign _GEN_491 = csr_wen ? _GEN_344 : {{34'd0}, reg_pmp_3_addr}; // @[CSR.scala 900:18]
  assign _GEN_498 = csr_wen ? _GEN_351 : {{34'd0}, reg_pmp_4_addr}; // @[CSR.scala 900:18]
  assign _GEN_505 = csr_wen ? _GEN_358 : {{34'd0}, reg_pmp_5_addr}; // @[CSR.scala 900:18]
  assign _GEN_512 = csr_wen ? _GEN_365 : {{34'd0}, reg_pmp_6_addr}; // @[CSR.scala 900:18]
  assign _GEN_519 = csr_wen ? _GEN_372 : {{34'd0}, reg_pmp_7_addr}; // @[CSR.scala 900:18]
  assign _io_trace_0_valid_T = io_retire > 1'h0; // @[CSR.scala 1165:26]
  assign io_rw_rdata = _io_rw_rdata_T_290 | _io_rw_rdata_T_146; // @[CSR.scala 855:15]
  assign io_decode_0_fp_illegal = _io_decode_0_fp_illegal_T | ~reg_misa[5]; // @[CSR.scala 667:23]
  assign io_decode_0_fp_csr = _io_decode_0_fp_csr_T == 12'h0; // @[CSR.scala 669:19]
  assign io_decode_0_read_illegal = _io_decode_0_read_illegal_T_317 | _io_decode_0_read_illegal_T_320; // @[CSR.scala 671:25]
  assign io_decode_0_write_illegal = &io_decode_0_csr[11:10]; // @[CSR.scala 678:26]
  assign io_decode_0_write_flush = ~_io_decode_0_write_flush_T_6; // @[CSR.scala 679:24]
  assign io_decode_0_system_illegal = _io_decode_0_system_illegal_T_14 | _io_decode_0_system_illegal_T_16; // @[CSR.scala 680:27]
  assign io_csr_stall = reg_wfi | io_status_cease; // @[CSR.scala 845:16]
  assign io_eret = _exception_T | insn_ret; // @[CSR.scala 726:11]
  assign io_singleStep = reg_dcsr_step & ~reg_debug; // @[CSR.scala 727:17]
  assign io_status_debug = reg_debug; // @[CSR.scala 728:13 CSR.scala 730:19]
  assign io_status_cease = io_status_cease_r; // @[CSR.scala 728:13 CSR.scala 846:19]
  assign io_status_wfi = reg_wfi; // @[CSR.scala 728:13 CSR.scala 847:17]
  assign io_status_isa = reg_misa[31:0]; // @[CSR.scala 728:13 CSR.scala 731:17]
  assign io_status_dprv = io_status_dprv_REG; // @[CSR.scala 728:13 CSR.scala 734:18]
  assign io_status_prv = reg_mstatus_prv; // @[CSR.scala 728:13]
  assign io_status_sd = _io_status_sd_T_2 | _io_status_sd_T_3; // @[CSR.scala 728:13 CSR.scala 729:16]
  assign io_status_zero2 = 27'h0; // @[CSR.scala 728:13]
  assign io_status_sxl = 2'h2; // @[CSR.scala 728:13 CSR.scala 733:17]
  assign io_status_uxl = 2'h2; // @[CSR.scala 728:13 CSR.scala 732:17]
  assign io_status_sd_rv32 = 1'h0; // @[CSR.scala 728:13]
  assign io_status_zero1 = 8'h0; // @[CSR.scala 728:13]
  assign io_status_tsr = reg_mstatus_tsr; // @[CSR.scala 728:13]
  assign io_status_tw = reg_mstatus_tw; // @[CSR.scala 728:13]
  assign io_status_tvm = reg_mstatus_tvm; // @[CSR.scala 728:13]
  assign io_status_mxr = reg_mstatus_mxr; // @[CSR.scala 728:13]
  assign io_status_sum = reg_mstatus_sum; // @[CSR.scala 728:13]
  assign io_status_mprv = reg_mstatus_mprv; // @[CSR.scala 728:13]
  assign io_status_xs = 2'h0; // @[CSR.scala 728:13]
  assign io_status_fs = reg_mstatus_fs; // @[CSR.scala 728:13]
  assign io_status_mpp = reg_mstatus_mpp; // @[CSR.scala 728:13]
  assign io_status_vs = 2'h0; // @[CSR.scala 728:13]
  assign io_status_spp = reg_mstatus_spp; // @[CSR.scala 728:13]
  assign io_status_mpie = reg_mstatus_mpie; // @[CSR.scala 728:13]
  assign io_status_hpie = 1'h0; // @[CSR.scala 728:13]
  assign io_status_spie = reg_mstatus_spie; // @[CSR.scala 728:13]
  assign io_status_upie = 1'h0; // @[CSR.scala 728:13]
  assign io_status_mie = reg_mstatus_mie; // @[CSR.scala 728:13]
  assign io_status_hie = 1'h0; // @[CSR.scala 728:13]
  assign io_status_sie = reg_mstatus_sie; // @[CSR.scala 728:13]
  assign io_status_uie = 1'h0; // @[CSR.scala 728:13]
  assign io_ptbr_mode = reg_satp_mode; // @[CSR.scala 725:11]
  assign io_ptbr_ppn = reg_satp_ppn; // @[CSR.scala 725:11]
  assign io_evec = _GEN_172[39:0]; // @[CSR.scala 724:11 CSR.scala 820:15 CSR.scala 824:15 CSR.scala 829:15 CSR.scala 835:15]
  assign io_time = {value_hi_1,value_lo_1}; // @[CSR.scala 844:11]
  assign io_fcsr_rm = reg_frm; // @[CSR.scala 885:14]
  assign io_interrupt = _io_interrupt_T_2 & ~_io_interrupt_T_3; // @[CSR.scala 469:16]
  assign io_interrupt_cause = 64'h8000000000000000 + _GEN_556; // @[CSR.scala 470:22]
  assign io_bp_0_control_action = reg_bp_0_control_action; // @[CSR.scala 471:9]
  assign io_bp_0_control_tmatch = reg_bp_0_control_tmatch; // @[CSR.scala 471:9]
  assign io_bp_0_control_m = reg_bp_0_control_m; // @[CSR.scala 471:9]
  assign io_bp_0_control_s = reg_bp_0_control_s; // @[CSR.scala 471:9]
  assign io_bp_0_control_u = reg_bp_0_control_u; // @[CSR.scala 471:9]
  assign io_bp_0_control_x = reg_bp_0_control_x; // @[CSR.scala 471:9]
  assign io_bp_0_control_w = reg_bp_0_control_w; // @[CSR.scala 471:9]
  assign io_bp_0_control_r = reg_bp_0_control_r; // @[CSR.scala 471:9]
  assign io_bp_0_address = reg_bp_0_address; // @[CSR.scala 471:9]
  assign io_pmp_0_cfg_l = reg_pmp_0_cfg_l; // @[CSR.scala 474:10]
  assign io_pmp_0_cfg_a = reg_pmp_0_cfg_a; // @[CSR.scala 474:10]
  assign io_pmp_0_cfg_x = reg_pmp_0_cfg_x; // @[CSR.scala 474:10]
  assign io_pmp_0_cfg_w = reg_pmp_0_cfg_w; // @[CSR.scala 474:10]
  assign io_pmp_0_cfg_r = reg_pmp_0_cfg_r; // @[CSR.scala 474:10]
  assign io_pmp_0_addr = reg_pmp_0_addr; // @[CSR.scala 474:10]
  assign io_pmp_0_mask = _pmp_mask_T_3[31:0]; // @[CSR.scala 474:10]
  assign io_pmp_1_cfg_l = reg_pmp_1_cfg_l; // @[CSR.scala 474:10]
  assign io_pmp_1_cfg_a = reg_pmp_1_cfg_a; // @[CSR.scala 474:10]
  assign io_pmp_1_cfg_x = reg_pmp_1_cfg_x; // @[CSR.scala 474:10]
  assign io_pmp_1_cfg_w = reg_pmp_1_cfg_w; // @[CSR.scala 474:10]
  assign io_pmp_1_cfg_r = reg_pmp_1_cfg_r; // @[CSR.scala 474:10]
  assign io_pmp_1_addr = reg_pmp_1_addr; // @[CSR.scala 474:10]
  assign io_pmp_1_mask = _pmp_mask_T_7[31:0]; // @[CSR.scala 474:10]
  assign io_pmp_2_cfg_l = reg_pmp_2_cfg_l; // @[CSR.scala 474:10]
  assign io_pmp_2_cfg_a = reg_pmp_2_cfg_a; // @[CSR.scala 474:10]
  assign io_pmp_2_cfg_x = reg_pmp_2_cfg_x; // @[CSR.scala 474:10]
  assign io_pmp_2_cfg_w = reg_pmp_2_cfg_w; // @[CSR.scala 474:10]
  assign io_pmp_2_cfg_r = reg_pmp_2_cfg_r; // @[CSR.scala 474:10]
  assign io_pmp_2_addr = reg_pmp_2_addr; // @[CSR.scala 474:10]
  assign io_pmp_2_mask = _pmp_mask_T_11[31:0]; // @[CSR.scala 474:10]
  assign io_pmp_3_cfg_l = reg_pmp_3_cfg_l; // @[CSR.scala 474:10]
  assign io_pmp_3_cfg_a = reg_pmp_3_cfg_a; // @[CSR.scala 474:10]
  assign io_pmp_3_cfg_x = reg_pmp_3_cfg_x; // @[CSR.scala 474:10]
  assign io_pmp_3_cfg_w = reg_pmp_3_cfg_w; // @[CSR.scala 474:10]
  assign io_pmp_3_cfg_r = reg_pmp_3_cfg_r; // @[CSR.scala 474:10]
  assign io_pmp_3_addr = reg_pmp_3_addr; // @[CSR.scala 474:10]
  assign io_pmp_3_mask = _pmp_mask_T_15[31:0]; // @[CSR.scala 474:10]
  assign io_pmp_4_cfg_l = reg_pmp_4_cfg_l; // @[CSR.scala 474:10]
  assign io_pmp_4_cfg_a = reg_pmp_4_cfg_a; // @[CSR.scala 474:10]
  assign io_pmp_4_cfg_x = reg_pmp_4_cfg_x; // @[CSR.scala 474:10]
  assign io_pmp_4_cfg_w = reg_pmp_4_cfg_w; // @[CSR.scala 474:10]
  assign io_pmp_4_cfg_r = reg_pmp_4_cfg_r; // @[CSR.scala 474:10]
  assign io_pmp_4_addr = reg_pmp_4_addr; // @[CSR.scala 474:10]
  assign io_pmp_4_mask = _pmp_mask_T_19[31:0]; // @[CSR.scala 474:10]
  assign io_pmp_5_cfg_l = reg_pmp_5_cfg_l; // @[CSR.scala 474:10]
  assign io_pmp_5_cfg_a = reg_pmp_5_cfg_a; // @[CSR.scala 474:10]
  assign io_pmp_5_cfg_x = reg_pmp_5_cfg_x; // @[CSR.scala 474:10]
  assign io_pmp_5_cfg_w = reg_pmp_5_cfg_w; // @[CSR.scala 474:10]
  assign io_pmp_5_cfg_r = reg_pmp_5_cfg_r; // @[CSR.scala 474:10]
  assign io_pmp_5_addr = reg_pmp_5_addr; // @[CSR.scala 474:10]
  assign io_pmp_5_mask = _pmp_mask_T_23[31:0]; // @[CSR.scala 474:10]
  assign io_pmp_6_cfg_l = reg_pmp_6_cfg_l; // @[CSR.scala 474:10]
  assign io_pmp_6_cfg_a = reg_pmp_6_cfg_a; // @[CSR.scala 474:10]
  assign io_pmp_6_cfg_x = reg_pmp_6_cfg_x; // @[CSR.scala 474:10]
  assign io_pmp_6_cfg_w = reg_pmp_6_cfg_w; // @[CSR.scala 474:10]
  assign io_pmp_6_cfg_r = reg_pmp_6_cfg_r; // @[CSR.scala 474:10]
  assign io_pmp_6_addr = reg_pmp_6_addr; // @[CSR.scala 474:10]
  assign io_pmp_6_mask = _pmp_mask_T_27[31:0]; // @[CSR.scala 474:10]
  assign io_pmp_7_cfg_l = reg_pmp_7_cfg_l; // @[CSR.scala 474:10]
  assign io_pmp_7_cfg_a = reg_pmp_7_cfg_a; // @[CSR.scala 474:10]
  assign io_pmp_7_cfg_x = reg_pmp_7_cfg_x; // @[CSR.scala 474:10]
  assign io_pmp_7_cfg_w = reg_pmp_7_cfg_w; // @[CSR.scala 474:10]
  assign io_pmp_7_cfg_r = reg_pmp_7_cfg_r; // @[CSR.scala 474:10]
  assign io_pmp_7_addr = reg_pmp_7_addr; // @[CSR.scala 474:10]
  assign io_pmp_7_mask = _pmp_mask_T_31[31:0]; // @[CSR.scala 474:10]
  assign io_inhibit_cycle = reg_mcountinhibit[0]; // @[CSR.scala 437:20]
  assign io_trace_0_valid = _io_trace_0_valid_T | io_trace_0_exception; // @[CSR.scala 1165:13]
  assign io_trace_0_iaddr = io_pc; // @[CSR.scala 1167:13]
  assign io_trace_0_insn = io_inst_0; // @[CSR.scala 1166:12]
  assign io_trace_0_priv = {reg_debug,reg_mstatus_prv}; // @[CSR.scala 1168:12]
  assign io_trace_0_exception = _exception_T | io_exception; // @[CSR.scala 1164:17]
  assign io_trace_0_interrupt = cause[63]; // @[CSR.scala 1170:17]
  assign io_trace_0_cause = insn_call ? {{60'd0}, _cause_T_1} : _cause_T_2; // @[CSR.scala 1169:13]
  assign io_trace_0_tval = io_tval; // @[CSR.scala 1171:12]
  assign io_customCSRs_0_value = reg_custom_0; // @[CSR.scala 852:14]
  assign CSRFile_cov_read_addr = CSRFile_state;
  assign CSRFile_cov_read_data = CSRFile_cov[CSRFile_cov_read_addr]; // @[Coverage map for CSRFile]
  assign CSRFile_cov_write_data = 1'h1;
  assign CSRFile_cov_write_addr = CSRFile_state;
  assign CSRFile_cov_write_mask = 1'h1;
  assign CSRFile_cov_write_en = 1'h1;
  assign reg_pmp_5_cfg_l_shl = {reg_pmp_5_cfg_l, 19'h0};
  assign reg_pmp_5_cfg_l_pad = reg_pmp_5_cfg_l_shl;
  assign reg_debug_shl = {reg_debug, 1'h0};
  assign reg_debug_pad = {18'h0,reg_debug_shl};
  assign reg_mstatus_sie_shl = {reg_mstatus_sie, 16'h0};
  assign reg_mstatus_sie_pad = {3'h0,reg_mstatus_sie_shl};
  assign reg_dcsr_prv_shl = {reg_dcsr_prv, 13'h0};
  assign reg_dcsr_prv_pad = {5'h0,reg_dcsr_prv_shl};
  assign reg_mcountinhibit_shl = {reg_mcountinhibit, 15'h0};
  assign reg_mcountinhibit_pad = {2'h0,reg_mcountinhibit_shl};
  assign reg_unmie_shl = {reg_unmie, 2'h0};
  assign reg_unmie_pad = {17'h0,reg_unmie_shl};
  assign reg_pmp_7_cfg_a_shl = {reg_pmp_7_cfg_a, 13'h0};
  assign reg_pmp_7_cfg_a_pad = {5'h0,reg_pmp_7_cfg_a_shl};
  assign reg_mstatus_mpp_shl = reg_mstatus_mpp;
  assign reg_mstatus_mpp_pad = {18'h0,reg_mstatus_mpp_shl};
  assign reg_pmp_2_cfg_l_shl = {reg_pmp_2_cfg_l, 6'h0};
  assign reg_pmp_2_cfg_l_pad = {13'h0,reg_pmp_2_cfg_l_shl};
  assign reg_pmp_1_cfg_l_shl = {reg_pmp_1_cfg_l, 18'h0};
  assign reg_pmp_1_cfg_l_pad = {1'h0,reg_pmp_1_cfg_l_shl};
  assign reg_mip_seip_shl = {reg_mip_seip, 9'h0};
  assign reg_mip_seip_pad = {10'h0,reg_mip_seip_shl};
  assign reg_rnmie_shl = {reg_rnmie, 1'h0};
  assign reg_rnmie_pad = {18'h0,reg_rnmie_shl};
  assign reg_mip_ssip_shl = {reg_mip_ssip, 10'h0};
  assign reg_mip_ssip_pad = {9'h0,reg_mip_ssip_shl};
  assign reg_bp_0_control_dmode_shl = {reg_bp_0_control_dmode, 2'h0};
  assign reg_bp_0_control_dmode_pad = {17'h0,reg_bp_0_control_dmode_shl};
  assign reg_pmp_4_cfg_l_shl = {reg_pmp_4_cfg_l, 11'h0};
  assign reg_pmp_4_cfg_l_pad = {8'h0,reg_pmp_4_cfg_l_shl};
  assign reg_dcsr_ebreaks_shl = {reg_dcsr_ebreaks, 1'h0};
  assign reg_dcsr_ebreaks_pad = {18'h0,reg_dcsr_ebreaks_shl};
  assign reg_pmp_6_cfg_l_shl = {reg_pmp_6_cfg_l, 13'h0};
  assign reg_pmp_6_cfg_l_pad = {6'h0,reg_pmp_6_cfg_l_shl};
  assign reg_mstatus_prv_shl = {reg_mstatus_prv, 2'h0};
  assign reg_mstatus_prv_pad = {16'h0,reg_mstatus_prv_shl};
  assign reg_dcsr_ebreakm_shl = {reg_dcsr_ebreakm, 8'h0};
  assign reg_dcsr_ebreakm_pad = {11'h0,reg_dcsr_ebreakm_shl};
  assign reg_pmp_7_cfg_l_shl = reg_pmp_7_cfg_l;
  assign reg_pmp_7_cfg_l_pad = {19'h0,reg_pmp_7_cfg_l_shl};
  assign reg_pmp_0_cfg_l_shl = {reg_pmp_0_cfg_l, 18'h0};
  assign reg_pmp_0_cfg_l_pad = {1'h0,reg_pmp_0_cfg_l_shl};
  assign reg_pmp_3_cfg_l_shl = {reg_pmp_3_cfg_l, 1'h0};
  assign reg_pmp_3_cfg_l_pad = {18'h0,reg_pmp_3_cfg_l_shl};
  assign reg_mstatus_spp_shl = {reg_mstatus_spp, 13'h0};
  assign reg_mstatus_spp_pad = {6'h0,reg_mstatus_spp_shl};
  assign reg_mip_stip_shl = {reg_mip_stip, 12'h0};
  assign reg_mip_stip_pad = {7'h0,reg_mip_stip_shl};
  assign reg_dcsr_ebreaku_shl = {reg_dcsr_ebreaku, 13'h0};
  assign reg_dcsr_ebreaku_pad = {6'h0,reg_dcsr_ebreaku_shl};
  assign reg_mstatus_mprv_shl = reg_mstatus_mprv;
  assign reg_mstatus_mprv_pad = {19'h0,reg_mstatus_mprv_shl};
  assign reg_singleStepped_shl = {reg_singleStepped, 13'h0};
  assign reg_singleStepped_pad = {6'h0,reg_singleStepped_shl};
  assign reg_mstatus_mie_shl = {reg_mstatus_mie, 11'h0};
  assign reg_mstatus_mie_pad = {8'h0,reg_mstatus_mie_shl};
  assign CSRFile_xor16 = reg_debug_pad ^ reg_mstatus_sie_pad;
  assign CSRFile_xor7 = reg_pmp_5_cfg_l_pad ^ CSRFile_xor16;
  assign CSRFile_xor17 = reg_dcsr_prv_pad ^ reg_mcountinhibit_pad;
  assign CSRFile_xor18 = reg_unmie_pad ^ reg_pmp_7_cfg_a_pad;
  assign CSRFile_xor8 = CSRFile_xor17 ^ CSRFile_xor18;
  assign CSRFile_xor3 = CSRFile_xor7 ^ CSRFile_xor8;
  assign CSRFile_xor20 = reg_pmp_2_cfg_l_pad ^ reg_pmp_1_cfg_l_pad;
  assign CSRFile_xor9 = reg_mstatus_mpp_pad ^ CSRFile_xor20;
  assign CSRFile_xor21 = reg_mip_seip_pad ^ reg_rnmie_pad;
  assign CSRFile_xor22 = reg_mip_ssip_pad ^ reg_bp_0_control_dmode_pad;
  assign CSRFile_xor10 = CSRFile_xor21 ^ CSRFile_xor22;
  assign CSRFile_xor4 = CSRFile_xor9 ^ CSRFile_xor10;
  assign CSRFile_xor1 = CSRFile_xor3 ^ CSRFile_xor4;
  assign CSRFile_xor24 = reg_dcsr_ebreaks_pad ^ reg_pmp_6_cfg_l_pad;
  assign CSRFile_xor11 = reg_pmp_4_cfg_l_pad ^ CSRFile_xor24;
  assign CSRFile_xor25 = reg_mstatus_prv_pad ^ reg_dcsr_ebreakm_pad;
  assign CSRFile_xor26 = reg_pmp_7_cfg_l_pad ^ reg_pmp_0_cfg_l_pad;
  assign CSRFile_xor12 = CSRFile_xor25 ^ CSRFile_xor26;
  assign CSRFile_xor5 = CSRFile_xor11 ^ CSRFile_xor12;
  assign CSRFile_xor28 = reg_mstatus_spp_pad ^ reg_mip_stip_pad;
  assign CSRFile_xor13 = reg_pmp_3_cfg_l_pad ^ CSRFile_xor28;
  assign CSRFile_xor29 = reg_dcsr_ebreaku_pad ^ reg_mstatus_mprv_pad;
  assign CSRFile_xor30 = reg_singleStepped_pad ^ reg_mstatus_mie_pad;
  assign CSRFile_xor14 = CSRFile_xor29 ^ CSRFile_xor30;
  assign CSRFile_xor6 = CSRFile_xor13 ^ CSRFile_xor14;
  assign CSRFile_xor2 = CSRFile_xor5 ^ CSRFile_xor6;
  assign CSRFile_xor0 = CSRFile_xor1 ^ CSRFile_xor2;
  assign io_covSum = CSRFile_covSum;
  assign stopEn0 = ~_T_252;
  assign stopEn1 = ~_T_274;
  assign CSRFile_or0 = stopEn0 | stopEn1;
  assign metaAssert = CSRFile_metaAssert;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_mstatus_prv = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  reg_mstatus_tsr = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  reg_mstatus_tw = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  reg_mstatus_tvm = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  reg_mstatus_mxr = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  reg_mstatus_sum = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  reg_mstatus_mprv = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  reg_mstatus_fs = _RAND_7[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  reg_mstatus_mpp = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  reg_mstatus_spp = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  reg_mstatus_mpie = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  reg_mstatus_spie = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  reg_mstatus_mie = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  reg_mstatus_sie = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  reg_dcsr_prv = _RAND_14[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  reg_singleStepped = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  reg_dcsr_ebreakm = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  reg_dcsr_ebreaks = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  reg_dcsr_ebreaku = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  reg_debug = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  reg_rnmie = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  reg_unmie = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {2{`RANDOM}};
  reg_mideleg = _RAND_22[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {2{`RANDOM}};
  reg_medeleg = _RAND_23[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  reg_dcsr_cause = _RAND_24[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  reg_dcsr_step = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {2{`RANDOM}};
  reg_dpc = _RAND_26[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {2{`RANDOM}};
  reg_dscratch = _RAND_27[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  reg_bp_0_control_dmode = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  reg_bp_0_control_action = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  reg_bp_0_control_tmatch = _RAND_30[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  reg_bp_0_control_m = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  reg_bp_0_control_s = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  reg_bp_0_control_u = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  reg_bp_0_control_x = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  reg_bp_0_control_w = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  reg_bp_0_control_r = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {2{`RANDOM}};
  reg_bp_0_address = _RAND_37[38:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  reg_pmp_0_cfg_l = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  reg_pmp_0_cfg_a = _RAND_39[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  reg_pmp_0_cfg_x = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  reg_pmp_0_cfg_w = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  reg_pmp_0_cfg_r = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  reg_pmp_0_addr = _RAND_43[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  reg_pmp_1_cfg_l = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  reg_pmp_1_cfg_a = _RAND_45[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  reg_pmp_1_cfg_x = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  reg_pmp_1_cfg_w = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  reg_pmp_1_cfg_r = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  reg_pmp_1_addr = _RAND_49[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  reg_pmp_2_cfg_l = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  reg_pmp_2_cfg_a = _RAND_51[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  reg_pmp_2_cfg_x = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  reg_pmp_2_cfg_w = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  reg_pmp_2_cfg_r = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  reg_pmp_2_addr = _RAND_55[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  reg_pmp_3_cfg_l = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  reg_pmp_3_cfg_a = _RAND_57[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  reg_pmp_3_cfg_x = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  reg_pmp_3_cfg_w = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  reg_pmp_3_cfg_r = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  reg_pmp_3_addr = _RAND_61[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  reg_pmp_4_cfg_l = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  reg_pmp_4_cfg_a = _RAND_63[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  reg_pmp_4_cfg_x = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  reg_pmp_4_cfg_w = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  reg_pmp_4_cfg_r = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  reg_pmp_4_addr = _RAND_67[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  reg_pmp_5_cfg_l = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  reg_pmp_5_cfg_a = _RAND_69[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  reg_pmp_5_cfg_x = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  reg_pmp_5_cfg_w = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  reg_pmp_5_cfg_r = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  reg_pmp_5_addr = _RAND_73[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  reg_pmp_6_cfg_l = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  reg_pmp_6_cfg_a = _RAND_75[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  reg_pmp_6_cfg_x = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  reg_pmp_6_cfg_w = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  reg_pmp_6_cfg_r = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  reg_pmp_6_addr = _RAND_79[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  reg_pmp_7_cfg_l = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  reg_pmp_7_cfg_a = _RAND_81[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  reg_pmp_7_cfg_x = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  reg_pmp_7_cfg_w = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  reg_pmp_7_cfg_r = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  reg_pmp_7_addr = _RAND_85[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {2{`RANDOM}};
  reg_mie = _RAND_86[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  reg_mip_seip = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  reg_mip_stip = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  reg_mip_ssip = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {2{`RANDOM}};
  reg_mepc = _RAND_90[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {2{`RANDOM}};
  reg_mcause = _RAND_91[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {2{`RANDOM}};
  reg_mtval = _RAND_92[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {2{`RANDOM}};
  reg_mscratch = _RAND_93[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  reg_mtvec = _RAND_94[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  reg_mcounteren = _RAND_95[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  reg_scounteren = _RAND_96[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {2{`RANDOM}};
  reg_sepc = _RAND_97[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {2{`RANDOM}};
  reg_scause = _RAND_98[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {2{`RANDOM}};
  reg_stval = _RAND_99[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {2{`RANDOM}};
  reg_sscratch = _RAND_100[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {2{`RANDOM}};
  reg_stvec = _RAND_101[38:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  reg_satp_mode = _RAND_102[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {2{`RANDOM}};
  reg_satp_ppn = _RAND_103[43:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  reg_wfi = _RAND_104[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  reg_fflags = _RAND_105[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  reg_frm = _RAND_106[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  reg_mcountinhibit = _RAND_107[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  value_lo = _RAND_108[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {2{`RANDOM}};
  value_hi = _RAND_109[57:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  value_lo_1 = _RAND_110[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {2{`RANDOM}};
  value_hi_1 = _RAND_111[57:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {2{`RANDOM}};
  reg_misa = _RAND_112[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {2{`RANDOM}};
  reg_custom_0 = _RAND_113[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  io_status_dprv_REG = _RAND_114[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  io_status_cease_r = _RAND_115[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  CSRFile_state = _RAND_116[19:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1048576; initvar = initvar+1)
    CSRFile_cov[initvar] = _RAND_117[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  CSRFile_covSum = _RAND_118[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  CSRFile_metaAssert = _RAND_119[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      reg_mstatus_prv <= 2'h0;
    end else if (reset) begin
      reg_mstatus_prv <= 2'h3;
    end else if (_reg_mstatus_prv_T) begin
      reg_mstatus_prv <= 2'h0;
    end else if (insn_ret) begin
      if (~io_rw_addr[9]) begin
        reg_mstatus_prv <= {{1'd0}, reg_mstatus_spp};
      end else if (_T_406) begin
        reg_mstatus_prv <= reg_dcsr_prv;
      end else begin
        reg_mstatus_prv <= reg_mstatus_mpp;
      end
    end else if (exception) begin
      if (trapToDebug) begin
        if (~reg_debug) begin
          reg_mstatus_prv <= 2'h3;
        end
      end else if (_T_279) begin
        reg_mstatus_prv <= 2'h1;
      end else begin
        reg_mstatus_prv <= 2'h3;
      end
    end
    if (metaReset) begin
      reg_mstatus_tsr <= 1'h0;
    end else if (reset) begin
      reg_mstatus_tsr <= 1'h0;
    end else if (csr_wen) begin
      if (_T_50) begin
        reg_mstatus_tsr <= new_mstatus_tsr;
      end
    end
    if (metaReset) begin
      reg_mstatus_tw <= 1'h0;
    end else if (reset) begin
      reg_mstatus_tw <= 1'h0;
    end else if (csr_wen) begin
      if (_T_50) begin
        reg_mstatus_tw <= new_mstatus_tw;
      end
    end
    if (metaReset) begin
      reg_mstatus_tvm <= 1'h0;
    end else if (reset) begin
      reg_mstatus_tvm <= 1'h0;
    end else if (csr_wen) begin
      if (_T_50) begin
        reg_mstatus_tvm <= new_mstatus_tvm;
      end
    end
    if (metaReset) begin
      reg_mstatus_mxr <= 1'h0;
    end else if (reset) begin
      reg_mstatus_mxr <= 1'h0;
    end else if (csr_wen) begin
      if (_T_158) begin
        reg_mstatus_mxr <= new_mstatus_mxr;
      end else if (_T_50) begin
        reg_mstatus_mxr <= new_mstatus_mxr;
      end
    end
    if (metaReset) begin
      reg_mstatus_sum <= 1'h0;
    end else if (reset) begin
      reg_mstatus_sum <= 1'h0;
    end else if (csr_wen) begin
      if (_T_158) begin
        reg_mstatus_sum <= new_mstatus_sum;
      end else if (_T_50) begin
        reg_mstatus_sum <= new_mstatus_sum;
      end
    end
    if (metaReset) begin
      reg_mstatus_mprv <= 1'h0;
    end else if (reset) begin
      reg_mstatus_mprv <= 1'h0;
    end else if (csr_wen) begin
      if (_T_50) begin
        reg_mstatus_mprv <= new_mstatus_mprv;
      end else if (insn_ret) begin
        if (_T_412) begin
          reg_mstatus_mprv <= 1'h0;
        end
      end
    end else if (insn_ret) begin
      if (_T_412) begin
        reg_mstatus_mprv <= 1'h0;
      end
    end
    if (metaReset) begin
      reg_mstatus_fs <= 2'h0;
    end else if (reset) begin
      reg_mstatus_fs <= 2'h0;
    end else if (csr_wen) begin
      if (_T_158) begin
        if (_reg_mstatus_fs_T) begin
          reg_mstatus_fs <= 2'h3;
        end else begin
          reg_mstatus_fs <= 2'h0;
        end
      end else if (_T_50) begin
        if (_reg_mstatus_fs_T) begin
          reg_mstatus_fs <= 2'h3;
        end else begin
          reg_mstatus_fs <= 2'h0;
        end
      end
    end
    if (metaReset) begin
      reg_mstatus_mpp <= 2'h0;
    end else if (reset) begin
      reg_mstatus_mpp <= 2'h3;
    end else if (csr_wen) begin
      if (_T_50) begin
        if (_reg_mstatus_mpp_T_2) begin
          reg_mstatus_mpp <= 2'h0;
        end else begin
          reg_mstatus_mpp <= new_mstatus_mpp;
        end
      end else if (insn_ret) begin
        if (~io_rw_addr[9]) begin
          if (exception) begin
            if (!(trapToDebug)) begin
              if (!(_T_279)) begin
                reg_mstatus_mpp <= reg_mstatus_prv;
              end
            end
          end
        end else if (_T_406) begin
          if (exception) begin
            if (!(trapToDebug)) begin
              if (!(_T_279)) begin
                reg_mstatus_mpp <= reg_mstatus_prv;
              end
            end
          end
        end else begin
          reg_mstatus_mpp <= 2'h0;
        end
      end else if (exception) begin
        if (!(trapToDebug)) begin
          if (!(_T_279)) begin
            reg_mstatus_mpp <= reg_mstatus_prv;
          end
        end
      end
    end else if (insn_ret) begin
      if (~io_rw_addr[9]) begin
        if (exception) begin
          if (!(trapToDebug)) begin
            if (!(_T_279)) begin
              reg_mstatus_mpp <= reg_mstatus_prv;
            end
          end
        end
      end else if (_T_406) begin
        reg_mstatus_mpp <= _GEN_140;
      end else begin
        reg_mstatus_mpp <= 2'h0;
      end
    end else begin
      reg_mstatus_mpp <= _GEN_140;
    end
    if (metaReset) begin
      reg_mstatus_spp <= 1'h0;
    end else if (reset) begin
      reg_mstatus_spp <= 1'h0;
    end else begin
      reg_mstatus_spp <= _GEN_385[0];
    end
    if (metaReset) begin
      reg_mstatus_mpie <= 1'h0;
    end else if (reset) begin
      reg_mstatus_mpie <= 1'h0;
    end else if (csr_wen) begin
      if (_T_50) begin
        reg_mstatus_mpie <= new_mstatus_mpie;
      end else if (insn_ret) begin
        if (~io_rw_addr[9]) begin
          if (exception) begin
            if (!(trapToDebug)) begin
              if (!(_T_279)) begin
                reg_mstatus_mpie <= reg_mstatus_mie;
              end
            end
          end
        end else if (_T_406) begin
          if (exception) begin
            if (!(trapToDebug)) begin
              if (!(_T_279)) begin
                reg_mstatus_mpie <= reg_mstatus_mie;
              end
            end
          end
        end else begin
          reg_mstatus_mpie <= 1'h1;
        end
      end else if (exception) begin
        if (!(trapToDebug)) begin
          if (!(_T_279)) begin
            reg_mstatus_mpie <= reg_mstatus_mie;
          end
        end
      end
    end else if (insn_ret) begin
      if (~io_rw_addr[9]) begin
        if (exception) begin
          if (!(trapToDebug)) begin
            if (!(_T_279)) begin
              reg_mstatus_mpie <= reg_mstatus_mie;
            end
          end
        end
      end else if (_T_406) begin
        reg_mstatus_mpie <= _GEN_139;
      end else begin
        reg_mstatus_mpie <= 1'h1;
      end
    end else begin
      reg_mstatus_mpie <= _GEN_139;
    end
    if (metaReset) begin
      reg_mstatus_spie <= 1'h0;
    end else if (reset) begin
      reg_mstatus_spie <= 1'h0;
    end else if (csr_wen) begin
      if (_T_158) begin
        reg_mstatus_spie <= new_mstatus_spie;
      end else if (_T_50) begin
        reg_mstatus_spie <= new_mstatus_spie;
      end else if (insn_ret) begin
        reg_mstatus_spie <= _GEN_158;
      end else if (exception) begin
        if (!(trapToDebug)) begin
          if (_T_279) begin
            reg_mstatus_spie <= reg_mstatus_sie;
          end
        end
      end
    end else if (insn_ret) begin
      reg_mstatus_spie <= _GEN_158;
    end else if (exception) begin
      if (!(trapToDebug)) begin
        if (_T_279) begin
          reg_mstatus_spie <= reg_mstatus_sie;
        end
      end
    end
    if (metaReset) begin
      reg_mstatus_mie <= 1'h0;
    end else if (reset) begin
      reg_mstatus_mie <= 1'h0;
    end else if (csr_wen) begin
      if (_T_50) begin
        reg_mstatus_mie <= new_mstatus_mie;
      end else if (insn_ret) begin
        if (~io_rw_addr[9]) begin
          if (exception) begin
            if (!(trapToDebug)) begin
              reg_mstatus_mie <= _GEN_76;
            end
          end
        end else if (_T_406) begin
          if (exception) begin
            if (!(trapToDebug)) begin
              reg_mstatus_mie <= _GEN_76;
            end
          end
        end else begin
          reg_mstatus_mie <= reg_mstatus_mpie;
        end
      end else if (exception) begin
        if (!(trapToDebug)) begin
          reg_mstatus_mie <= _GEN_76;
        end
      end
    end else if (insn_ret) begin
      if (~io_rw_addr[9]) begin
        if (exception) begin
          if (!(trapToDebug)) begin
            reg_mstatus_mie <= _GEN_76;
          end
        end
      end else if (_T_406) begin
        reg_mstatus_mie <= _GEN_141;
      end else begin
        reg_mstatus_mie <= reg_mstatus_mpie;
      end
    end else begin
      reg_mstatus_mie <= _GEN_141;
    end
    if (metaReset) begin
      reg_mstatus_sie <= 1'h0;
    end else if (reset) begin
      reg_mstatus_sie <= 1'h0;
    end else if (csr_wen) begin
      if (_T_158) begin
        reg_mstatus_sie <= new_mstatus_sie;
      end else if (_T_50) begin
        reg_mstatus_sie <= new_mstatus_sie;
      end else if (insn_ret) begin
        if (~io_rw_addr[9]) begin
          reg_mstatus_sie <= reg_mstatus_spie;
        end else if (exception) begin
          if (!(trapToDebug)) begin
            if (_T_279) begin
              reg_mstatus_sie <= 1'h0;
            end
          end
        end
      end else if (exception) begin
        if (!(trapToDebug)) begin
          if (_T_279) begin
            reg_mstatus_sie <= 1'h0;
          end
        end
      end
    end else if (insn_ret) begin
      if (~io_rw_addr[9]) begin
        reg_mstatus_sie <= reg_mstatus_spie;
      end else if (exception) begin
        if (!(trapToDebug)) begin
          if (_T_279) begin
            reg_mstatus_sie <= 1'h0;
          end
        end
      end
    end else if (exception) begin
      if (!(trapToDebug)) begin
        if (_T_279) begin
          reg_mstatus_sie <= 1'h0;
        end
      end
    end
    if (metaReset) begin
      reg_dcsr_prv <= 2'h0;
    end else if (reset) begin
      reg_dcsr_prv <= 2'h3;
    end else if (csr_wen) begin
      if (_T_59) begin
        if (_reg_dcsr_prv_T) begin
          reg_dcsr_prv <= 2'h0;
        end else begin
          reg_dcsr_prv <= new_dcsr_prv;
        end
      end else if (exception) begin
        if (trapToDebug) begin
          if (~reg_debug) begin
            reg_dcsr_prv <= reg_mstatus_prv;
          end
        end
      end
    end else if (exception) begin
      if (trapToDebug) begin
        if (~reg_debug) begin
          reg_dcsr_prv <= reg_mstatus_prv;
        end
      end
    end
    if (metaReset) begin
      reg_singleStepped <= 1'h0;
    end else if (~io_singleStep) begin
      reg_singleStepped <= 1'h0;
    end else begin
      reg_singleStepped <= _GEN_50;
    end
    if (metaReset) begin
      reg_dcsr_ebreakm <= 1'h0;
    end else if (reset) begin
      reg_dcsr_ebreakm <= 1'h0;
    end else if (csr_wen) begin
      if (_T_59) begin
        reg_dcsr_ebreakm <= new_dcsr_ebreakm;
      end
    end
    if (metaReset) begin
      reg_dcsr_ebreaks <= 1'h0;
    end else if (reset) begin
      reg_dcsr_ebreaks <= 1'h0;
    end else if (csr_wen) begin
      if (_T_59) begin
        reg_dcsr_ebreaks <= new_dcsr_ebreaks;
      end
    end
    if (metaReset) begin
      reg_dcsr_ebreaku <= 1'h0;
    end else if (reset) begin
      reg_dcsr_ebreaku <= 1'h0;
    end else if (csr_wen) begin
      if (_T_59) begin
        reg_dcsr_ebreaku <= new_dcsr_ebreaku;
      end
    end
    if (metaReset) begin
      //if (rv_dv) begin
        reg_debug <= 1'h0; //SC
      //end
      //else begin
      //  reg_debug <= 1'h1;
      //end	
    end else if (reset) begin
      //if (rv_dv) begin
        reg_debug <= 1'h0; //SC
      //end
      //else begin
      //  reg_debug <= 1'h1;
      //end
    end else if (insn_ret) begin
      if (~io_rw_addr[9]) begin
        if (exception) begin
          if (trapToDebug) begin
            reg_debug <= _GEN_52;
          end
        end
      end else if (_T_406) begin
        reg_debug <= 1'h0;
      end else if (exception) begin
        if (trapToDebug) begin
          reg_debug <= _GEN_52;
        end
      end
    end else if (exception) begin
      if (trapToDebug) begin
        reg_debug <= _GEN_52;
      end
    end
    if (metaReset) begin
      reg_rnmie <= 1'h0;
    end else begin
      reg_rnmie <= reset | reg_rnmie;
    end
    if (metaReset) begin
      reg_unmie <= 1'h0;
    end else begin
      reg_unmie <= reset | reg_unmie;
    end
    if (metaReset) begin
      reg_mideleg <= 64'h0;
    end else if (csr_wen) begin
      if (_T_168) begin
        reg_mideleg <= wdata;
      end
    end
    if (metaReset) begin
      reg_medeleg <= 64'h0;
    end else if (csr_wen) begin
      if (_T_169) begin
        reg_medeleg <= wdata;
      end
    end
    if (metaReset) begin
      reg_dcsr_cause <= 3'h0;
    end else if (reset) begin
      reg_dcsr_cause <= 3'h0;
    end else if (exception) begin
      if (trapToDebug) begin
        if (~reg_debug) begin
          if (reg_singleStepped) begin
            reg_dcsr_cause <= 3'h4;
          end else begin
            reg_dcsr_cause <= {{1'd0}, _reg_dcsr_cause_T_1};
          end
        end
      end
    end
    if (metaReset) begin
      reg_dcsr_step <= 1'h0;
    end else if (reset) begin
      reg_dcsr_step <= 1'h0;
    end else if (csr_wen) begin
      if (_T_59) begin
        reg_dcsr_step <= new_dcsr_step;
      end
    end
    if (metaReset) begin
      reg_dpc <= 40'h0;
    end else begin
      reg_dpc <= _GEN_418[39:0];
    end
    if (metaReset) begin
      reg_dscratch <= 64'h0;
    end else if (csr_wen) begin
      if (_T_61) begin
        reg_dscratch <= wdata;
      end
    end
    if (metaReset) begin
      reg_bp_0_control_dmode <= 1'h0;
    end else if (reset) begin
      reg_bp_0_control_dmode <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1842) begin
        if (_T_46) begin
          reg_bp_0_control_dmode <= dMode;
        end
      end
    end
    if (metaReset) begin
      reg_bp_0_control_action <= 1'h0;
    end else if (reset) begin
      reg_bp_0_control_action <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1842) begin
        if (_T_46) begin
          reg_bp_0_control_action <= _GEN_252;
        end
      end
    end
    if (metaReset) begin
      reg_bp_0_control_tmatch <= 2'h0;
    end else if (csr_wen) begin
      if (_T_1842) begin
        if (_T_46) begin
          reg_bp_0_control_tmatch <= wdata[8:7];
        end
      end
    end
    if (metaReset) begin
      reg_bp_0_control_m <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1842) begin
        if (_T_46) begin
          reg_bp_0_control_m <= wdata[6];
        end
      end
    end
    if (metaReset) begin
      reg_bp_0_control_s <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1842) begin
        if (_T_46) begin
          reg_bp_0_control_s <= wdata[4];
        end
      end
    end
    if (metaReset) begin
      reg_bp_0_control_u <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1842) begin
        if (_T_46) begin
          reg_bp_0_control_u <= wdata[3];
        end
      end
    end
    if (metaReset) begin
      reg_bp_0_control_x <= 1'h0;
    end else if (reset) begin
      reg_bp_0_control_x <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1842) begin
        if (_T_46) begin
          reg_bp_0_control_x <= wdata[2];
        end
      end
    end
    if (metaReset) begin
      reg_bp_0_control_w <= 1'h0;
    end else if (reset) begin
      reg_bp_0_control_w <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1842) begin
        if (_T_46) begin
          reg_bp_0_control_w <= wdata[1];
        end
      end
    end
    if (metaReset) begin
      reg_bp_0_control_r <= 1'h0;
    end else if (reset) begin
      reg_bp_0_control_r <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1842) begin
        if (_T_46) begin
          reg_bp_0_control_r <= wdata[0];
        end
      end
    end
    if (metaReset) begin
      reg_bp_0_address <= 39'h0;
    end else begin
      reg_bp_0_address <= _GEN_432[38:0];
    end
    if (metaReset) begin
      reg_pmp_0_cfg_l <= 1'h0;
    end else if (reset) begin
      reg_pmp_0_cfg_l <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1853) begin
        reg_pmp_0_cfg_l <= newCfg_l;
      end
    end
    if (metaReset) begin
      reg_pmp_0_cfg_a <= 2'h0;
    end else if (reset) begin
      reg_pmp_0_cfg_a <= 2'h0;
    end else if (csr_wen) begin
      if (_T_1853) begin
        reg_pmp_0_cfg_a <= newCfg_a;
      end
    end
    if (metaReset) begin
      reg_pmp_0_cfg_x <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1853) begin
        reg_pmp_0_cfg_x <= newCfg_x;
      end
    end
    if (metaReset) begin
      reg_pmp_0_cfg_w <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1853) begin
        reg_pmp_0_cfg_w <= _reg_pmp_0_cfg_w_T;
      end
    end
    if (metaReset) begin
      reg_pmp_0_cfg_r <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1853) begin
        reg_pmp_0_cfg_r <= newCfg_r;
      end
    end
    if (metaReset) begin
      reg_pmp_0_addr <= 30'h0;
    end else begin
      reg_pmp_0_addr <= _GEN_470[29:0];
    end
    if (metaReset) begin
      reg_pmp_1_cfg_l <= 1'h0;
    end else if (reset) begin
      reg_pmp_1_cfg_l <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1863) begin
        reg_pmp_1_cfg_l <= newCfg_1_l;
      end
    end
    if (metaReset) begin
      reg_pmp_1_cfg_a <= 2'h0;
    end else if (reset) begin
      reg_pmp_1_cfg_a <= 2'h0;
    end else if (csr_wen) begin
      if (_T_1863) begin
        reg_pmp_1_cfg_a <= newCfg_1_a;
      end
    end
    if (metaReset) begin
      reg_pmp_1_cfg_x <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1863) begin
        reg_pmp_1_cfg_x <= newCfg_1_x;
      end
    end
    if (metaReset) begin
      reg_pmp_1_cfg_w <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1863) begin
        reg_pmp_1_cfg_w <= _reg_pmp_1_cfg_w_T;
      end
    end
    if (metaReset) begin
      reg_pmp_1_cfg_r <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1863) begin
        reg_pmp_1_cfg_r <= newCfg_1_r;
      end
    end
    if (metaReset) begin
      reg_pmp_1_addr <= 30'h0;
    end else begin
      reg_pmp_1_addr <= _GEN_477[29:0];
    end
    if (metaReset) begin
      reg_pmp_2_cfg_l <= 1'h0;
    end else if (reset) begin
      reg_pmp_2_cfg_l <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1873) begin
        reg_pmp_2_cfg_l <= newCfg_2_l;
      end
    end
    if (metaReset) begin
      reg_pmp_2_cfg_a <= 2'h0;
    end else if (reset) begin
      reg_pmp_2_cfg_a <= 2'h0;
    end else if (csr_wen) begin
      if (_T_1873) begin
        reg_pmp_2_cfg_a <= newCfg_2_a;
      end
    end
    if (metaReset) begin
      reg_pmp_2_cfg_x <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1873) begin
        reg_pmp_2_cfg_x <= newCfg_2_x;
      end
    end
    if (metaReset) begin
      reg_pmp_2_cfg_w <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1873) begin
        reg_pmp_2_cfg_w <= _reg_pmp_2_cfg_w_T;
      end
    end
    if (metaReset) begin
      reg_pmp_2_cfg_r <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1873) begin
        reg_pmp_2_cfg_r <= newCfg_2_r;
      end
    end
    if (metaReset) begin
      reg_pmp_2_addr <= 30'h0;
    end else begin
      reg_pmp_2_addr <= _GEN_484[29:0];
    end
    if (metaReset) begin
      reg_pmp_3_cfg_l <= 1'h0;
    end else if (reset) begin
      reg_pmp_3_cfg_l <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1883) begin
        reg_pmp_3_cfg_l <= newCfg_3_l;
      end
    end
    if (metaReset) begin
      reg_pmp_3_cfg_a <= 2'h0;
    end else if (reset) begin
      reg_pmp_3_cfg_a <= 2'h0;
    end else if (csr_wen) begin
      if (_T_1883) begin
        reg_pmp_3_cfg_a <= newCfg_3_a;
      end
    end
    if (metaReset) begin
      reg_pmp_3_cfg_x <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1883) begin
        reg_pmp_3_cfg_x <= newCfg_3_x;
      end
    end
    if (metaReset) begin
      reg_pmp_3_cfg_w <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1883) begin
        reg_pmp_3_cfg_w <= _reg_pmp_3_cfg_w_T;
      end
    end
    if (metaReset) begin
      reg_pmp_3_cfg_r <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1883) begin
        reg_pmp_3_cfg_r <= newCfg_3_r;
      end
    end
    if (metaReset) begin
      reg_pmp_3_addr <= 30'h0;
    end else begin
      reg_pmp_3_addr <= _GEN_491[29:0];
    end
    if (metaReset) begin
      reg_pmp_4_cfg_l <= 1'h0;
    end else if (reset) begin
      reg_pmp_4_cfg_l <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1893) begin
        reg_pmp_4_cfg_l <= newCfg_4_l;
      end
    end
    if (metaReset) begin
      reg_pmp_4_cfg_a <= 2'h0;
    end else if (reset) begin
      reg_pmp_4_cfg_a <= 2'h0;
    end else if (csr_wen) begin
      if (_T_1893) begin
        reg_pmp_4_cfg_a <= newCfg_4_a;
      end
    end
    if (metaReset) begin
      reg_pmp_4_cfg_x <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1893) begin
        reg_pmp_4_cfg_x <= newCfg_4_x;
      end
    end
    if (metaReset) begin
      reg_pmp_4_cfg_w <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1893) begin
        reg_pmp_4_cfg_w <= _reg_pmp_4_cfg_w_T;
      end
    end
    if (metaReset) begin
      reg_pmp_4_cfg_r <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1893) begin
        reg_pmp_4_cfg_r <= newCfg_4_r;
      end
    end
    if (metaReset) begin
      reg_pmp_4_addr <= 30'h0;
    end else begin
      reg_pmp_4_addr <= _GEN_498[29:0];
    end
    if (metaReset) begin
      reg_pmp_5_cfg_l <= 1'h0;
    end else if (reset) begin
      reg_pmp_5_cfg_l <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1903) begin
        reg_pmp_5_cfg_l <= newCfg_5_l;
      end
    end
    if (metaReset) begin
      reg_pmp_5_cfg_a <= 2'h0;
    end else if (reset) begin
      reg_pmp_5_cfg_a <= 2'h0;
    end else if (csr_wen) begin
      if (_T_1903) begin
        reg_pmp_5_cfg_a <= newCfg_5_a;
      end
    end
    if (metaReset) begin
      reg_pmp_5_cfg_x <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1903) begin
        reg_pmp_5_cfg_x <= newCfg_5_x;
      end
    end
    if (metaReset) begin
      reg_pmp_5_cfg_w <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1903) begin
        reg_pmp_5_cfg_w <= _reg_pmp_5_cfg_w_T;
      end
    end
    if (metaReset) begin
      reg_pmp_5_cfg_r <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1903) begin
        reg_pmp_5_cfg_r <= newCfg_5_r;
      end
    end
    if (metaReset) begin
      reg_pmp_5_addr <= 30'h0;
    end else begin
      reg_pmp_5_addr <= _GEN_505[29:0];
    end
    if (metaReset) begin
      reg_pmp_6_cfg_l <= 1'h0;
    end else if (reset) begin
      reg_pmp_6_cfg_l <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1913) begin
        reg_pmp_6_cfg_l <= newCfg_6_l;
      end
    end
    if (metaReset) begin
      reg_pmp_6_cfg_a <= 2'h0;
    end else if (reset) begin
      reg_pmp_6_cfg_a <= 2'h0;
    end else if (csr_wen) begin
      if (_T_1913) begin
        reg_pmp_6_cfg_a <= newCfg_6_a;
      end
    end
    if (metaReset) begin
      reg_pmp_6_cfg_x <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1913) begin
        reg_pmp_6_cfg_x <= newCfg_6_x;
      end
    end
    if (metaReset) begin
      reg_pmp_6_cfg_w <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1913) begin
        reg_pmp_6_cfg_w <= _reg_pmp_6_cfg_w_T;
      end
    end
    if (metaReset) begin
      reg_pmp_6_cfg_r <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1913) begin
        reg_pmp_6_cfg_r <= newCfg_6_r;
      end
    end
    if (metaReset) begin
      reg_pmp_6_addr <= 30'h0;
    end else begin
      reg_pmp_6_addr <= _GEN_512[29:0];
    end
    if (metaReset) begin
      reg_pmp_7_cfg_l <= 1'h0;
    end else if (reset) begin
      reg_pmp_7_cfg_l <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1923) begin
        reg_pmp_7_cfg_l <= newCfg_7_l;
      end
    end
    if (metaReset) begin
      reg_pmp_7_cfg_a <= 2'h0;
    end else if (reset) begin
      reg_pmp_7_cfg_a <= 2'h0;
    end else if (csr_wen) begin
      if (_T_1923) begin
        reg_pmp_7_cfg_a <= newCfg_7_a;
      end
    end
    if (metaReset) begin
      reg_pmp_7_cfg_x <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1923) begin
        reg_pmp_7_cfg_x <= newCfg_7_x;
      end
    end
    if (metaReset) begin
      reg_pmp_7_cfg_w <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1923) begin
        reg_pmp_7_cfg_w <= _reg_pmp_7_cfg_w_T;
      end
    end
    if (metaReset) begin
      reg_pmp_7_cfg_r <= 1'h0;
    end else if (csr_wen) begin
      if (_T_1923) begin
        reg_pmp_7_cfg_r <= newCfg_7_r;
      end
    end
    if (metaReset) begin
      reg_pmp_7_addr <= 30'h0;
    end else begin
      reg_pmp_7_addr <= _GEN_519[29:0];
    end
    if (metaReset) begin
      reg_mie <= 64'h0;
    end else if (csr_wen) begin
      if (_T_160) begin
        reg_mie <= _reg_mie_T_4;
      end else if (_T_53) begin
        reg_mie <= _reg_mie_T;
      end
    end
    if (metaReset) begin
      reg_mip_seip <= 1'h0;
    end else if (csr_wen) begin
      if (_T_52) begin
        reg_mip_seip <= new_mip_seip;
      end
    end
    if (metaReset) begin
      reg_mip_stip <= 1'h0;
    end else if (csr_wen) begin
      if (_T_52) begin
        reg_mip_stip <= new_mip_stip;
      end
    end
    if (metaReset) begin
      reg_mip_ssip <= 1'h0;
    end else if (csr_wen) begin
      if (_T_159) begin
        reg_mip_ssip <= new_sip_ssip;
      end else if (_T_52) begin
        reg_mip_ssip <= new_mip_ssip;
      end
    end
    if (metaReset) begin
      reg_mepc <= 40'h0;
    end else begin
      reg_mepc <= _GEN_400[39:0];
    end
    if (metaReset) begin
      reg_mcause <= 64'h0;
    end else if (reset) begin
      reg_mcause <= 64'h0;
    end else if (csr_wen) begin
      if (_T_57) begin
        reg_mcause <= _reg_mcause_T;
      end else if (exception) begin
        if (!(trapToDebug)) begin
          if (!(_T_279)) begin
            if (insn_call) begin
              reg_mcause <= {{60'd0}, _cause_T_1};
            end else if (insn_break) begin
              reg_mcause <= 64'h3;
            end else begin
              reg_mcause <= io_cause;
            end
          end
        end
      end
    end else if (exception) begin
      if (!(trapToDebug)) begin
        if (!(_T_279)) begin
          if (insn_call) begin
            reg_mcause <= {{60'd0}, _cause_T_1};
          end else if (insn_break) begin
            reg_mcause <= 64'h3;
          end else begin
            reg_mcause <= io_cause;
          end
        end
      end
    end
    if (metaReset) begin
      reg_mtval <= 40'h0;
    end else if (csr_wen) begin
      if (_T_56) begin
        reg_mtval <= wdata[39:0];
      end else if (exception) begin
        if (!(trapToDebug)) begin
          if (!(_T_279)) begin
            reg_mtval <= io_tval;
          end
        end
      end
    end else if (exception) begin
      if (!(trapToDebug)) begin
        if (!(_T_279)) begin
          reg_mtval <= io_tval;
        end
      end
    end
    if (metaReset) begin
      reg_mscratch <= 64'h0;
    end else if (csr_wen) begin
      if (_T_54) begin
        reg_mscratch <= wdata;
      end
    end
    if (metaReset) begin
      reg_mtvec <= 32'h0;
    end else if (reset) begin
      reg_mtvec <= 32'h0;
    end else begin
      reg_mtvec <= _GEN_402[31:0];
    end
    if (metaReset) begin
      reg_mcounteren <= 32'h0;
    end else begin
      reg_mcounteren <= _GEN_430[31:0];
    end
    if (metaReset) begin
      reg_scounteren <= 32'h0;
    end else begin
      reg_scounteren <= _GEN_429[31:0];
    end
    if (metaReset) begin
      reg_sepc <= 40'h0;
    end else begin
      reg_sepc <= _GEN_423[39:0];
    end
    if (metaReset) begin
      reg_scause <= 64'h0;
    end else if (csr_wen) begin
      if (_T_162) begin
        reg_scause <= _reg_scause_T;
      end else if (exception) begin
        if (!(trapToDebug)) begin
          if (_T_279) begin
            if (insn_call) begin
              reg_scause <= {{60'd0}, _cause_T_1};
            end else if (insn_break) begin
              reg_scause <= 64'h3;
            end else begin
              reg_scause <= io_cause;
            end
          end
        end
      end
    end else if (exception) begin
      if (!(trapToDebug)) begin
        if (_T_279) begin
          if (insn_call) begin
            reg_scause <= {{60'd0}, _cause_T_1};
          end else if (insn_break) begin
            reg_scause <= 64'h3;
          end else begin
            reg_scause <= io_cause;
          end
        end
      end
    end
    if (metaReset) begin
      reg_stval <= 40'h0;
    end else if (csr_wen) begin
      if (_T_163) begin
        reg_stval <= wdata[39:0];
      end else if (exception) begin
        if (!(trapToDebug)) begin
          if (_T_279) begin
            reg_stval <= io_tval;
          end
        end
      end
    end else if (exception) begin
      if (!(trapToDebug)) begin
        if (_T_279) begin
          reg_stval <= io_tval;
        end
      end
    end
    if (metaReset) begin
      reg_sscratch <= 64'h0;
    end else if (csr_wen) begin
      if (_T_161) begin
        reg_sscratch <= wdata;
      end
    end
    if (metaReset) begin
      reg_stvec <= 39'h0;
    end else begin
      reg_stvec <= _GEN_424[38:0];
    end
    if (metaReset) begin
      reg_satp_mode <= 4'h0;
    end else if (csr_wen) begin
      if (_T_164) begin
        if (_T_1839) begin
          reg_satp_mode <= _reg_satp_mode_T;
        end
      end
    end
    if (metaReset) begin
      reg_satp_ppn <= 44'h0;
    end else if (csr_wen) begin
      if (_T_164) begin
        if (_T_1839) begin
          reg_satp_ppn <= {{24'd0}, new_satp_ppn[19:0]};
        end
      end
    end
    if (metaReset) begin
      reg_fflags <= 5'h0;
    end else begin
      reg_fflags <= _GEN_411[4:0];
    end
    if (metaReset) begin
      reg_frm <= 3'h0;
    end else begin
      reg_frm <= _GEN_412[2:0];
    end
    if (metaReset) begin
      reg_mcountinhibit <= 3'h0;
    end else if (reset) begin
      reg_mcountinhibit <= 3'h0;
    end else begin
      reg_mcountinhibit <= _GEN_405[2:0];
    end
    if (metaReset) begin
      value_lo <= 6'h0;
    end else if (reset) begin
      value_lo <= 6'h0;
    end else begin
      value_lo <= _GEN_408[5:0];
    end
    if (metaReset) begin
      value_hi <= 58'h0;
    end else if (reset) begin
      value_hi <= 58'h0;
    end else if (csr_wen) begin
      if (_T_67) begin
        value_hi <= wdata[63:6];
      end else if (_large_T_2) begin
        value_hi <= _large_r_T_1;
      end
    end else if (_large_T_2) begin
      value_hi <= _large_r_T_1;
    end
    if (metaReset) begin
      value_lo_1 <= 6'h0;
    end else if (reset) begin
      value_lo_1 <= 6'h0;
    end else begin
      value_lo_1 <= _GEN_406[5:0];
    end
    if (metaReset) begin
      value_hi_1 <= 58'h0;
    end else if (reset) begin
      value_hi_1 <= 58'h0;
    end else if (csr_wen) begin
      if (_T_66) begin
        value_hi_1 <= wdata[63:6];
      end else if (_large_T_5) begin
        value_hi_1 <= _large_r_T_3;
      end
    end else if (_large_T_5) begin
      value_hi_1 <= _large_r_T_3;
    end
    if (metaReset) begin
      reg_misa <= 64'h0;
    end else if (reset) begin
      reg_misa <= 64'h800000000094112d;
    end else if (csr_wen) begin
      if (_T_49) begin
        if (_T_1834) begin
          reg_misa <= _reg_misa_T_8;
        end
      end
    end
    if (metaReset) begin
      reg_custom_0 <= 64'h0;
    end else if (reset) begin
      reg_custom_0 <= 64'h208;
    end else if (csr_wen) begin
      if (_T_188) begin
        reg_custom_0 <= _reg_custom_0_T_3;
      end
    end
    if (metaReset) begin
      io_status_dprv_REG <= 2'h0;
    end else if (_io_status_dprv_x87_T_1) begin
      io_status_dprv_REG <= reg_mstatus_mpp;
    end else begin
      io_status_dprv_REG <= reg_mstatus_prv;
    end
    if (metaReset) begin
      io_status_cease_r <= 1'h0;
    end else if (reset) begin
      io_status_cease_r <= 1'h0;
    end else begin
      io_status_cease_r <= _GEN_181;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_252) begin
          $fwrite(32'h80000002,"Assertion failed: these conditions must be mutually exclusive\n    at CSR.scala:739 assert(PopCount(insn_ret :: insn_call :: insn_break :: io.exception :: Nil) <= 1, \"these conditions must be mutually exclusive\")\n"); // @[CSR.scala 739:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_252) begin
          $fatal; // @[CSR.scala 739:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_274) begin
          $fwrite(32'h80000002,"Assertion failed\n    at CSR.scala:748 assert(!reg_singleStepped || io.retire === UInt(0))\n"); // @[CSR.scala 748:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_274) begin
          $fatal; // @[CSR.scala 748:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    CSRFile_state <= CSRFile_xor0;
    if (!(CSRFile_cov_read_data)) begin
      CSRFile_covSum <= CSRFile_covSum + 1'h1;
    end
    if (metaReset) begin
      CSRFile_metaAssert <= 1'h0;
    end else begin
      CSRFile_metaAssert <= CSRFile_metaAssert | CSRFile_or0;
    end
  end
  always @(posedge io_ungated_clock) begin
    if (metaReset) begin
      reg_wfi <= 1'h0;
    end else if (reset) begin
      reg_wfi <= 1'h0;
    end else if (_T_260) begin
      reg_wfi <= 1'h0;
    end else begin
      reg_wfi <= _GEN_48;
    end
  end
  always @(posedge clock) begin
    if(CSRFile_cov_write_en & CSRFile_cov_write_mask) begin
      CSRFile_cov[CSRFile_cov_write_addr] <= CSRFile_cov_write_data; // @[Coverage map for CSRFile]
    end
  end
endmodule
module BreakpointUnit(
  input         io_status_debug,
  input  [1:0]  io_status_prv,
  input         io_bp_0_control_action,
  input  [1:0]  io_bp_0_control_tmatch,
  input         io_bp_0_control_m,
  input         io_bp_0_control_s,
  input         io_bp_0_control_u,
  input         io_bp_0_control_x,
  input         io_bp_0_control_w,
  input         io_bp_0_control_r,
  input  [38:0] io_bp_0_address,
  input  [38:0] io_pc,
  input  [38:0] io_ea,
  output        io_xcpt_if,
  output        io_xcpt_ld,
  output        io_xcpt_st,
  output        io_debug_if,
  output        io_debug_ld,
  output        io_debug_st,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire [3:0] _en_T_1; // @[Cat.scala 30:58]
  wire [3:0] _en_T_2; // @[Breakpoint.scala 31:68]
  wire  en; // @[Breakpoint.scala 31:50]
  wire  _r_T; // @[Breakpoint.scala 107:16]
  wire  _r_T_2; // @[Breakpoint.scala 66:8]
  wire  _r_T_4; // @[Breakpoint.scala 66:20]
  wire  r_lo_hi; // @[Breakpoint.scala 60:73]
  wire  r_hi_lo; // @[Breakpoint.scala 60:73]
  wire  r_hi_hi; // @[Breakpoint.scala 60:73]
  wire [3:0] _r_T_9; // @[Cat.scala 30:58]
  wire [38:0] _GEN_11; // @[Breakpoint.scala 63:9]
  wire [38:0] _r_T_10; // @[Breakpoint.scala 63:9]
  wire [38:0] _r_T_16; // @[Breakpoint.scala 63:33]
  wire  _r_T_17; // @[Breakpoint.scala 63:19]
  wire  _r_T_18; // @[Breakpoint.scala 69:8]
  wire  r; // @[Breakpoint.scala 107:32]
  wire  _w_T; // @[Breakpoint.scala 108:16]
  wire  w; // @[Breakpoint.scala 108:32]
  wire  _x_T; // @[Breakpoint.scala 109:16]
  wire  _x_T_2; // @[Breakpoint.scala 66:8]
  wire  _x_T_4; // @[Breakpoint.scala 66:20]
  wire [38:0] _x_T_10; // @[Breakpoint.scala 63:9]
  wire  _x_T_17; // @[Breakpoint.scala 63:19]
  wire  _x_T_18; // @[Breakpoint.scala 69:8]
  wire  x; // @[Breakpoint.scala 109:32]
  wire [29:0] BreakpointUnit_covSum;
  assign _en_T_1 = {io_bp_0_control_m,1'h0,io_bp_0_control_s,io_bp_0_control_u}; // @[Cat.scala 30:58]
  assign _en_T_2 = _en_T_1 >> io_status_prv; // @[Breakpoint.scala 31:68]
  assign en = ~io_status_debug & _en_T_2[0]; // @[Breakpoint.scala 31:50]
  assign _r_T = en & io_bp_0_control_r; // @[Breakpoint.scala 107:16]
  assign _r_T_2 = io_ea >= io_bp_0_address; // @[Breakpoint.scala 66:8]
  assign _r_T_4 = _r_T_2 ^ io_bp_0_control_tmatch[0]; // @[Breakpoint.scala 66:20]
  assign r_lo_hi = io_bp_0_control_tmatch[0] & io_bp_0_address[0]; // @[Breakpoint.scala 60:73]
  assign r_hi_lo = r_lo_hi & io_bp_0_address[1]; // @[Breakpoint.scala 60:73]
  assign r_hi_hi = r_hi_lo & io_bp_0_address[2]; // @[Breakpoint.scala 60:73]
  assign _r_T_9 = {r_hi_hi,r_hi_lo,r_lo_hi,io_bp_0_control_tmatch[0]}; // @[Cat.scala 30:58]
  assign _GEN_11 = {{35'd0}, _r_T_9}; // @[Breakpoint.scala 63:9]
  assign _r_T_10 = ~io_ea | _GEN_11; // @[Breakpoint.scala 63:9]
  assign _r_T_16 = ~io_bp_0_address | _GEN_11; // @[Breakpoint.scala 63:33]
  assign _r_T_17 = _r_T_10 == _r_T_16; // @[Breakpoint.scala 63:19]
  assign _r_T_18 = io_bp_0_control_tmatch[1] ? _r_T_4 : _r_T_17; // @[Breakpoint.scala 69:8]
  assign r = _r_T & _r_T_18; // @[Breakpoint.scala 107:32]
  assign _w_T = en & io_bp_0_control_w; // @[Breakpoint.scala 108:16]
  assign w = _w_T & _r_T_18; // @[Breakpoint.scala 108:32]
  assign _x_T = en & io_bp_0_control_x; // @[Breakpoint.scala 109:16]
  assign _x_T_2 = io_pc >= io_bp_0_address; // @[Breakpoint.scala 66:8]
  assign _x_T_4 = _x_T_2 ^ io_bp_0_control_tmatch[0]; // @[Breakpoint.scala 66:20]
  assign _x_T_10 = ~io_pc | _GEN_11; // @[Breakpoint.scala 63:9]
  assign _x_T_17 = _x_T_10 == _r_T_16; // @[Breakpoint.scala 63:19]
  assign _x_T_18 = io_bp_0_control_tmatch[1] ? _x_T_4 : _x_T_17; // @[Breakpoint.scala 69:8]
  assign x = _x_T & _x_T_18; // @[Breakpoint.scala 109:32]
  assign io_xcpt_if = x & ~io_bp_0_control_action; // @[Breakpoint.scala 97:14 Breakpoint.scala 121:40]
  assign io_xcpt_ld = r & ~io_bp_0_control_action; // @[Breakpoint.scala 98:14 Breakpoint.scala 119:40]
  assign io_xcpt_st = w & ~io_bp_0_control_action; // @[Breakpoint.scala 99:14 Breakpoint.scala 120:40]
  assign io_debug_if = x & io_bp_0_control_action; // @[Breakpoint.scala 100:15 Breakpoint.scala 121:73]
  assign io_debug_ld = r & io_bp_0_control_action; // @[Breakpoint.scala 101:15 Breakpoint.scala 119:73]
  assign io_debug_st = w & io_bp_0_control_action; // @[Breakpoint.scala 102:15 Breakpoint.scala 120:73]
  assign BreakpointUnit_covSum = 30'h0;
  assign io_covSum = BreakpointUnit_covSum;
  assign metaAssert = 1'h0;
endmodule
module ALU(
  input         io_dw,
  input  [3:0]  io_fn,
  input  [63:0] io_in2,
  input  [63:0] io_in1,
  output [63:0] io_out,
  output [63:0] io_adder_out,
  output        io_cmp_out,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire [63:0] in2_inv; // @[ALU.scala 61:20]
  wire [63:0] in1_xor_in2; // @[ALU.scala 62:28]
  wire [63:0] _io_adder_out_T_1; // @[ALU.scala 63:26]
  wire [63:0] _GEN_1; // @[ALU.scala 63:36]
  wire  _slt_T_2; // @[ALU.scala 67:24]
  wire  _slt_T_7; // @[ALU.scala 68:8]
  wire  slt; // @[ALU.scala 67:8]
  wire  _io_cmp_out_T_3; // @[ALU.scala 69:68]
  wire  _io_cmp_out_T_4; // @[ALU.scala 69:41]
  wire  _T_2; // @[ALU.scala 76:46]
  wire [31:0] _T_4; // @[Bitwise.scala 72:12]
  wire [31:0] hi; // @[ALU.scala 77:24]
  wire  hi_1; // @[ALU.scala 78:33]
  wire [4:0] lo; // @[ALU.scala 78:60]
  wire [5:0] shamt; // @[Cat.scala 30:58]
  wire [31:0] lo_1; // @[ALU.scala 79:34]
  wire [63:0] shin_r; // @[Cat.scala 30:58]
  wire  _shin_T; // @[ALU.scala 81:24]
  wire  _shin_T_1; // @[ALU.scala 81:44]
  wire  _shin_T_2; // @[ALU.scala 81:35]
  wire [63:0] _shin_T_6; // @[Bitwise.scala 103:31]
  wire [63:0] _shin_T_8; // @[Bitwise.scala 103:65]
  wire [63:0] _shin_T_10; // @[Bitwise.scala 103:75]
  wire [63:0] _shin_T_11; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_2; // @[Bitwise.scala 103:31]
  wire [63:0] _shin_T_16; // @[Bitwise.scala 103:31]
  wire [63:0] _shin_T_18; // @[Bitwise.scala 103:65]
  wire [63:0] _shin_T_20; // @[Bitwise.scala 103:75]
  wire [63:0] _shin_T_21; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_3; // @[Bitwise.scala 103:31]
  wire [63:0] _shin_T_26; // @[Bitwise.scala 103:31]
  wire [63:0] _shin_T_28; // @[Bitwise.scala 103:65]
  wire [63:0] _shin_T_30; // @[Bitwise.scala 103:75]
  wire [63:0] _shin_T_31; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_4; // @[Bitwise.scala 103:31]
  wire [63:0] _shin_T_36; // @[Bitwise.scala 103:31]
  wire [63:0] _shin_T_38; // @[Bitwise.scala 103:65]
  wire [63:0] _shin_T_40; // @[Bitwise.scala 103:75]
  wire [63:0] _shin_T_41; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_5; // @[Bitwise.scala 103:31]
  wire [63:0] _shin_T_46; // @[Bitwise.scala 103:31]
  wire [63:0] _shin_T_48; // @[Bitwise.scala 103:65]
  wire [63:0] _shin_T_50; // @[Bitwise.scala 103:75]
  wire [63:0] _shin_T_51; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_6; // @[Bitwise.scala 103:31]
  wire [63:0] _shin_T_56; // @[Bitwise.scala 103:31]
  wire [63:0] _shin_T_58; // @[Bitwise.scala 103:65]
  wire [63:0] _shin_T_60; // @[Bitwise.scala 103:75]
  wire [63:0] _shin_T_61; // @[Bitwise.scala 103:39]
  wire [63:0] shin; // @[ALU.scala 81:17]
  wire  shout_r_hi; // @[ALU.scala 82:35]
  wire [64:0] _shout_r_T_3; // @[ALU.scala 82:57]
  wire [64:0] _shout_r_T_4; // @[ALU.scala 82:64]
  wire [63:0] shout_r; // @[ALU.scala 82:73]
  wire [63:0] _shout_l_T_3; // @[Bitwise.scala 103:31]
  wire [63:0] _shout_l_T_5; // @[Bitwise.scala 103:65]
  wire [63:0] _shout_l_T_7; // @[Bitwise.scala 103:75]
  wire [63:0] _shout_l_T_8; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_7; // @[Bitwise.scala 103:31]
  wire [63:0] _shout_l_T_13; // @[Bitwise.scala 103:31]
  wire [63:0] _shout_l_T_15; // @[Bitwise.scala 103:65]
  wire [63:0] _shout_l_T_17; // @[Bitwise.scala 103:75]
  wire [63:0] _shout_l_T_18; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_8; // @[Bitwise.scala 103:31]
  wire [63:0] _shout_l_T_23; // @[Bitwise.scala 103:31]
  wire [63:0] _shout_l_T_25; // @[Bitwise.scala 103:65]
  wire [63:0] _shout_l_T_27; // @[Bitwise.scala 103:75]
  wire [63:0] _shout_l_T_28; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_9; // @[Bitwise.scala 103:31]
  wire [63:0] _shout_l_T_33; // @[Bitwise.scala 103:31]
  wire [63:0] _shout_l_T_35; // @[Bitwise.scala 103:65]
  wire [63:0] _shout_l_T_37; // @[Bitwise.scala 103:75]
  wire [63:0] _shout_l_T_38; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_10; // @[Bitwise.scala 103:31]
  wire [63:0] _shout_l_T_43; // @[Bitwise.scala 103:31]
  wire [63:0] _shout_l_T_45; // @[Bitwise.scala 103:65]
  wire [63:0] _shout_l_T_47; // @[Bitwise.scala 103:75]
  wire [63:0] _shout_l_T_48; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_11; // @[Bitwise.scala 103:31]
  wire [63:0] _shout_l_T_53; // @[Bitwise.scala 103:31]
  wire [63:0] _shout_l_T_55; // @[Bitwise.scala 103:65]
  wire [63:0] _shout_l_T_57; // @[Bitwise.scala 103:75]
  wire [63:0] shout_l; // @[Bitwise.scala 103:39]
  wire [63:0] _shout_T_3; // @[ALU.scala 84:18]
  wire  _shout_T_4; // @[ALU.scala 85:25]
  wire [63:0] _shout_T_5; // @[ALU.scala 85:18]
  wire [63:0] shout; // @[ALU.scala 84:74]
  wire  _logic_T; // @[ALU.scala 88:25]
  wire  _logic_T_1; // @[ALU.scala 88:45]
  wire  _logic_T_2; // @[ALU.scala 88:36]
  wire [63:0] _logic_T_3; // @[ALU.scala 88:18]
  wire  _logic_T_5; // @[ALU.scala 89:44]
  wire  _logic_T_6; // @[ALU.scala 89:35]
  wire [63:0] _logic_T_7; // @[ALU.scala 89:63]
  wire [63:0] _logic_T_8; // @[ALU.scala 89:18]
  wire [63:0] logic_; // @[ALU.scala 88:78]
  wire  _shift_logic_T; // @[ALU.scala 41:30]
  wire  _shift_logic_T_1; // @[ALU.scala 90:35]
  wire [63:0] _GEN_12; // @[ALU.scala 90:43]
  wire [63:0] _shift_logic_T_2; // @[ALU.scala 90:43]
  wire [63:0] shift_logic; // @[ALU.scala 90:51]
  wire  _out_T; // @[ALU.scala 91:23]
  wire  _out_T_1; // @[ALU.scala 91:43]
  wire  _out_T_2; // @[ALU.scala 91:34]
  wire [63:0] out; // @[ALU.scala 91:16]
  wire [31:0] io_out_hi; // @[Bitwise.scala 72:12]
  wire [31:0] io_out_lo; // @[ALU.scala 96:66]
  wire [63:0] _io_out_T_2; // @[Cat.scala 30:58]
  wire [29:0] ALU_covSum;
  assign in2_inv = io_fn[3] ? ~io_in2 : io_in2; // @[ALU.scala 61:20]
  assign in1_xor_in2 = io_in1 ^ in2_inv; // @[ALU.scala 62:28]
  assign _io_adder_out_T_1 = io_in1 + in2_inv; // @[ALU.scala 63:26]
  assign _GEN_1 = {{63'd0}, io_fn[3]}; // @[ALU.scala 63:36]
  assign _slt_T_2 = io_in1[63] == io_in2[63]; // @[ALU.scala 67:24]
  assign _slt_T_7 = io_fn[1] ? io_in2[63] : io_in1[63]; // @[ALU.scala 68:8]
  assign slt = _slt_T_2 ? io_adder_out[63] : _slt_T_7; // @[ALU.scala 67:8]
  assign _io_cmp_out_T_3 = in1_xor_in2 == 64'h0; // @[ALU.scala 69:68]
  assign _io_cmp_out_T_4 = io_fn[3] ? slt : _io_cmp_out_T_3; // @[ALU.scala 69:41]
  assign _T_2 = io_fn[3] & io_in1[31]; // @[ALU.scala 76:46]
  assign _T_4 = _T_2 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  assign hi = io_dw ? io_in1[63:32] : _T_4; // @[ALU.scala 77:24]
  assign hi_1 = io_in2[5] & io_dw; // @[ALU.scala 78:33]
  assign lo = io_in2[4:0]; // @[ALU.scala 78:60]
  assign shamt = {hi_1,lo}; // @[Cat.scala 30:58]
  assign lo_1 = io_in1[31:0]; // @[ALU.scala 79:34]
  assign shin_r = {hi,lo_1}; // @[Cat.scala 30:58]
  assign _shin_T = io_fn == 4'h5; // @[ALU.scala 81:24]
  assign _shin_T_1 = io_fn == 4'hb; // @[ALU.scala 81:44]
  assign _shin_T_2 = _shin_T | _shin_T_1; // @[ALU.scala 81:35]
  assign _shin_T_6 = {{32'd0}, shin_r[63:32]}; // @[Bitwise.scala 103:31]
  assign _shin_T_8 = {shin_r[31:0], 32'h0}; // @[Bitwise.scala 103:65]
  assign _shin_T_10 = _shin_T_8 & 64'hffffffff00000000; // @[Bitwise.scala 103:75]
  assign _shin_T_11 = _shin_T_6 | _shin_T_10; // @[Bitwise.scala 103:39]
  assign _GEN_2 = {{16'd0}, _shin_T_11[63:16]}; // @[Bitwise.scala 103:31]
  assign _shin_T_16 = _GEN_2 & 64'hffff0000ffff; // @[Bitwise.scala 103:31]
  assign _shin_T_18 = {_shin_T_11[47:0], 16'h0}; // @[Bitwise.scala 103:65]
  assign _shin_T_20 = _shin_T_18 & 64'hffff0000ffff0000; // @[Bitwise.scala 103:75]
  assign _shin_T_21 = _shin_T_16 | _shin_T_20; // @[Bitwise.scala 103:39]
  assign _GEN_3 = {{8'd0}, _shin_T_21[63:8]}; // @[Bitwise.scala 103:31]
  assign _shin_T_26 = _GEN_3 & 64'hff00ff00ff00ff; // @[Bitwise.scala 103:31]
  assign _shin_T_28 = {_shin_T_21[55:0], 8'h0}; // @[Bitwise.scala 103:65]
  assign _shin_T_30 = _shin_T_28 & 64'hff00ff00ff00ff00; // @[Bitwise.scala 103:75]
  assign _shin_T_31 = _shin_T_26 | _shin_T_30; // @[Bitwise.scala 103:39]
  assign _GEN_4 = {{4'd0}, _shin_T_31[63:4]}; // @[Bitwise.scala 103:31]
  assign _shin_T_36 = _GEN_4 & 64'hf0f0f0f0f0f0f0f; // @[Bitwise.scala 103:31]
  assign _shin_T_38 = {_shin_T_31[59:0], 4'h0}; // @[Bitwise.scala 103:65]
  assign _shin_T_40 = _shin_T_38 & 64'hf0f0f0f0f0f0f0f0; // @[Bitwise.scala 103:75]
  assign _shin_T_41 = _shin_T_36 | _shin_T_40; // @[Bitwise.scala 103:39]
  assign _GEN_5 = {{2'd0}, _shin_T_41[63:2]}; // @[Bitwise.scala 103:31]
  assign _shin_T_46 = _GEN_5 & 64'h3333333333333333; // @[Bitwise.scala 103:31]
  assign _shin_T_48 = {_shin_T_41[61:0], 2'h0}; // @[Bitwise.scala 103:65]
  assign _shin_T_50 = _shin_T_48 & 64'hcccccccccccccccc; // @[Bitwise.scala 103:75]
  assign _shin_T_51 = _shin_T_46 | _shin_T_50; // @[Bitwise.scala 103:39]
  assign _GEN_6 = {{1'd0}, _shin_T_51[63:1]}; // @[Bitwise.scala 103:31]
  assign _shin_T_56 = _GEN_6 & 64'h5555555555555555; // @[Bitwise.scala 103:31]
  assign _shin_T_58 = {_shin_T_51[62:0], 1'h0}; // @[Bitwise.scala 103:65]
  assign _shin_T_60 = _shin_T_58 & 64'haaaaaaaaaaaaaaaa; // @[Bitwise.scala 103:75]
  assign _shin_T_61 = _shin_T_56 | _shin_T_60; // @[Bitwise.scala 103:39]
  assign shin = _shin_T_2 ? shin_r : _shin_T_61; // @[ALU.scala 81:17]
  assign shout_r_hi = io_fn[3] & shin[63]; // @[ALU.scala 82:35]
  assign _shout_r_T_3 = {shout_r_hi,shin}; // @[ALU.scala 82:57]
  assign _shout_r_T_4 = $signed(_shout_r_T_3) >>> shamt; // @[ALU.scala 82:64]
  assign shout_r = _shout_r_T_4[63:0]; // @[ALU.scala 82:73]
  assign _shout_l_T_3 = {{32'd0}, shout_r[63:32]}; // @[Bitwise.scala 103:31]
  assign _shout_l_T_5 = {shout_r[31:0], 32'h0}; // @[Bitwise.scala 103:65]
  assign _shout_l_T_7 = _shout_l_T_5 & 64'hffffffff00000000; // @[Bitwise.scala 103:75]
  assign _shout_l_T_8 = _shout_l_T_3 | _shout_l_T_7; // @[Bitwise.scala 103:39]
  assign _GEN_7 = {{16'd0}, _shout_l_T_8[63:16]}; // @[Bitwise.scala 103:31]
  assign _shout_l_T_13 = _GEN_7 & 64'hffff0000ffff; // @[Bitwise.scala 103:31]
  assign _shout_l_T_15 = {_shout_l_T_8[47:0], 16'h0}; // @[Bitwise.scala 103:65]
  assign _shout_l_T_17 = _shout_l_T_15 & 64'hffff0000ffff0000; // @[Bitwise.scala 103:75]
  assign _shout_l_T_18 = _shout_l_T_13 | _shout_l_T_17; // @[Bitwise.scala 103:39]
  assign _GEN_8 = {{8'd0}, _shout_l_T_18[63:8]}; // @[Bitwise.scala 103:31]
  assign _shout_l_T_23 = _GEN_8 & 64'hff00ff00ff00ff; // @[Bitwise.scala 103:31]
  assign _shout_l_T_25 = {_shout_l_T_18[55:0], 8'h0}; // @[Bitwise.scala 103:65]
  assign _shout_l_T_27 = _shout_l_T_25 & 64'hff00ff00ff00ff00; // @[Bitwise.scala 103:75]
  assign _shout_l_T_28 = _shout_l_T_23 | _shout_l_T_27; // @[Bitwise.scala 103:39]
  assign _GEN_9 = {{4'd0}, _shout_l_T_28[63:4]}; // @[Bitwise.scala 103:31]
  assign _shout_l_T_33 = _GEN_9 & 64'hf0f0f0f0f0f0f0f; // @[Bitwise.scala 103:31]
  assign _shout_l_T_35 = {_shout_l_T_28[59:0], 4'h0}; // @[Bitwise.scala 103:65]
  assign _shout_l_T_37 = _shout_l_T_35 & 64'hf0f0f0f0f0f0f0f0; // @[Bitwise.scala 103:75]
  assign _shout_l_T_38 = _shout_l_T_33 | _shout_l_T_37; // @[Bitwise.scala 103:39]
  assign _GEN_10 = {{2'd0}, _shout_l_T_38[63:2]}; // @[Bitwise.scala 103:31]
  assign _shout_l_T_43 = _GEN_10 & 64'h3333333333333333; // @[Bitwise.scala 103:31]
  assign _shout_l_T_45 = {_shout_l_T_38[61:0], 2'h0}; // @[Bitwise.scala 103:65]
  assign _shout_l_T_47 = _shout_l_T_45 & 64'hcccccccccccccccc; // @[Bitwise.scala 103:75]
  assign _shout_l_T_48 = _shout_l_T_43 | _shout_l_T_47; // @[Bitwise.scala 103:39]
  assign _GEN_11 = {{1'd0}, _shout_l_T_48[63:1]}; // @[Bitwise.scala 103:31]
  assign _shout_l_T_53 = _GEN_11 & 64'h5555555555555555; // @[Bitwise.scala 103:31]
  assign _shout_l_T_55 = {_shout_l_T_48[62:0], 1'h0}; // @[Bitwise.scala 103:65]
  assign _shout_l_T_57 = _shout_l_T_55 & 64'haaaaaaaaaaaaaaaa; // @[Bitwise.scala 103:75]
  assign shout_l = _shout_l_T_53 | _shout_l_T_57; // @[Bitwise.scala 103:39]
  assign _shout_T_3 = _shin_T_2 ? shout_r : 64'h0; // @[ALU.scala 84:18]
  assign _shout_T_4 = io_fn == 4'h1; // @[ALU.scala 85:25]
  assign _shout_T_5 = _shout_T_4 ? shout_l : 64'h0; // @[ALU.scala 85:18]
  assign shout = _shout_T_3 | _shout_T_5; // @[ALU.scala 84:74]
  assign _logic_T = io_fn == 4'h4; // @[ALU.scala 88:25]
  assign _logic_T_1 = io_fn == 4'h6; // @[ALU.scala 88:45]
  assign _logic_T_2 = _logic_T | _logic_T_1; // @[ALU.scala 88:36]
  assign _logic_T_3 = _logic_T_2 ? in1_xor_in2 : 64'h0; // @[ALU.scala 88:18]
  assign _logic_T_5 = io_fn == 4'h7; // @[ALU.scala 89:44]
  assign _logic_T_6 = _logic_T_1 | _logic_T_5; // @[ALU.scala 89:35]
  assign _logic_T_7 = io_in1 & io_in2; // @[ALU.scala 89:63]
  assign _logic_T_8 = _logic_T_6 ? _logic_T_7 : 64'h0; // @[ALU.scala 89:18]
  assign logic_ = _logic_T_3 | _logic_T_8; // @[ALU.scala 88:78]
  assign _shift_logic_T = io_fn >= 4'hc; // @[ALU.scala 41:30]
  assign _shift_logic_T_1 = _shift_logic_T & slt; // @[ALU.scala 90:35]
  assign _GEN_12 = {{63'd0}, _shift_logic_T_1}; // @[ALU.scala 90:43]
  assign _shift_logic_T_2 = _GEN_12 | logic_; // @[ALU.scala 90:43]
  assign shift_logic = _shift_logic_T_2 | shout; // @[ALU.scala 90:51]
  assign _out_T = io_fn == 4'h0; // @[ALU.scala 91:23]
  assign _out_T_1 = io_fn == 4'ha; // @[ALU.scala 91:43]
  assign _out_T_2 = _out_T | _out_T_1; // @[ALU.scala 91:34]
  assign out = _out_T_2 ? io_adder_out : shift_logic; // @[ALU.scala 91:16]
  assign io_out_hi = out[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  assign io_out_lo = out[31:0]; // @[ALU.scala 96:66]
  assign _io_out_T_2 = {io_out_hi,io_out_lo}; // @[Cat.scala 30:58]
  assign io_out = io_dw ? out : _io_out_T_2; // @[ALU.scala 93:10 ALU.scala 96:37]
  assign io_adder_out = _io_adder_out_T_1 + _GEN_1; // @[ALU.scala 63:16]
  assign io_cmp_out = io_fn[0] ^ _io_cmp_out_T_4; // @[ALU.scala 69:14]
  assign ALU_covSum = 30'h0;
  assign io_covSum = ALU_covSum;
  assign metaAssert = 1'h0;
endmodule
module MulDiv(
  input         clock,
  input         reset,
  output        io_req_ready,
  input         io_req_valid,
  input  [3:0]  io_req_bits_fn,
  input         io_req_bits_dw,
  input  [63:0] io_req_bits_in1,
  input  [63:0] io_req_bits_in2,
  input  [4:0]  io_req_bits_tag,
  input         io_kill,
  input         io_resp_ready,
  output        io_resp_valid,
  output [63:0] io_resp_bits_data,
  output [4:0]  io_resp_bits_tag,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  reg [2:0] state; // @[Multiplier.scala 52:22]
  reg [31:0] _RAND_0;
  reg  req_dw; // @[Multiplier.scala 54:16]
  reg [31:0] _RAND_1;
  reg [4:0] req_tag; // @[Multiplier.scala 54:16]
  reg [31:0] _RAND_2;
  reg [6:0] count; // @[Multiplier.scala 55:18]
  reg [31:0] _RAND_3;
  reg  neg_out; // @[Multiplier.scala 58:20]
  reg [31:0] _RAND_4;
  reg  isHi; // @[Multiplier.scala 59:17]
  reg [31:0] _RAND_5;
  reg  resHi; // @[Multiplier.scala 60:18]
  reg [31:0] _RAND_6;
  reg [64:0] divisor; // @[Multiplier.scala 61:20]
  reg [95:0] _RAND_7;
  reg [129:0] remainder; // @[Multiplier.scala 62:22]
  reg [159:0] _RAND_8;
  wire [3:0] _T; // @[Decode.scala 14:65]
  wire  cmdMul; // @[Decode.scala 14:121]
  wire [3:0] _T_3; // @[Decode.scala 14:65]
  wire  _T_4; // @[Decode.scala 14:121]
  wire [3:0] _T_5; // @[Decode.scala 14:65]
  wire  _T_6; // @[Decode.scala 14:121]
  wire  cmdHi; // @[Decode.scala 15:30]
  wire [3:0] _T_9; // @[Decode.scala 14:65]
  wire  _T_10; // @[Decode.scala 14:121]
  wire [3:0] _T_11; // @[Decode.scala 14:65]
  wire  _T_12; // @[Decode.scala 14:121]
  wire  lhsSigned; // @[Decode.scala 15:30]
  wire  _T_16; // @[Decode.scala 14:121]
  wire  rhsSigned; // @[Decode.scala 15:30]
  wire  _sign_T_2; // @[Multiplier.scala 82:29]
  wire  lhs_sign; // @[Multiplier.scala 82:23]
  wire [31:0] _hi_T_1; // @[Bitwise.scala 72:12]
  wire [31:0] hi; // @[Multiplier.scala 83:17]
  wire [31:0] lo; // @[Multiplier.scala 84:15]
  wire [63:0] lhs_in; // @[Cat.scala 30:58]
  wire  _sign_T_5; // @[Multiplier.scala 82:29]
  wire  rhs_sign; // @[Multiplier.scala 82:23]
  wire [31:0] _hi_T_4; // @[Bitwise.scala 72:12]
  wire [31:0] hi_1; // @[Multiplier.scala 83:17]
  wire [31:0] lo_1; // @[Multiplier.scala 84:15]
  wire [64:0] subtractor; // @[Multiplier.scala 89:37]
  wire [63:0] result; // @[Multiplier.scala 90:19]
  wire [63:0] negated_remainder; // @[Multiplier.scala 91:27]
  wire  _T_23; // @[Multiplier.scala 93:39]
  wire  _T_26; // @[Multiplier.scala 102:39]
  wire  _T_27; // @[Multiplier.scala 107:39]
  wire [64:0] mulReg_hi; // @[Multiplier.scala 108:31]
  wire [128:0] mulReg; // @[Cat.scala 30:58]
  wire  prod_hi; // @[Multiplier.scala 109:31]
  wire [63:0] mplier; // @[Multiplier.scala 110:24]
  wire [64:0] accum; // @[Multiplier.scala 111:37]
  wire [7:0] prod_lo; // @[Multiplier.scala 113:38]
  wire [8:0] _prod_T_1; // @[Multiplier.scala 113:60]
  wire [64:0] _GEN_37; // @[Multiplier.scala 113:67]
  wire [73:0] _prod_T_2; // @[Multiplier.scala 113:67]
  wire [73:0] _GEN_38; // @[Multiplier.scala 113:76]
  wire [55:0] nextMulReg_lo; // @[Multiplier.scala 114:38]
  wire [73:0] nextMulReg_hi; // @[Cat.scala 30:58]
  wire [129:0] nextMulReg; // @[Cat.scala 30:58]
  wire  _nextMplierSign_T; // @[Multiplier.scala 115:32]
  wire  remainder_hi_lo; // @[Multiplier.scala 115:57]
  wire [10:0] _eOutMask_T; // @[Multiplier.scala 117:54]
  wire [64:0] _eOutMask_T_2; // @[Multiplier.scala 117:44]
  wire [63:0] eOutMask; // @[Multiplier.scala 117:89]
  wire  _eOut_T; // @[Multiplier.scala 118:45]
  wire  _eOut_T_2; // @[Multiplier.scala 118:79]
  wire  _eOut_T_3; // @[Multiplier.scala 118:70]
  wire  _eOut_T_5; // @[Multiplier.scala 118:85]
  wire [63:0] _eOut_T_7; // @[Multiplier.scala 119:24]
  wire  _eOut_T_8; // @[Multiplier.scala 119:37]
  wire  eOut; // @[Multiplier.scala 119:13]
  wire [10:0] _eOutRes_T_2; // @[Multiplier.scala 120:36]
  wire [128:0] eOutRes; // @[Multiplier.scala 120:27]
  wire [64:0] nextMulReg1_hi; // @[Multiplier.scala 121:37]
  wire [129:0] _nextMulReg1_T; // @[Multiplier.scala 121:55]
  wire [63:0] nextMulReg1_lo; // @[Multiplier.scala 121:82]
  wire [128:0] nextMulReg1; // @[Cat.scala 30:58]
  wire [64:0] remainder_hi_hi; // @[Multiplier.scala 122:34]
  wire [63:0] remainder_lo; // @[Multiplier.scala 122:67]
  wire [129:0] _remainder_T; // @[Cat.scala 30:58]
  wire [6:0] _count_T_1; // @[Multiplier.scala 124:20]
  wire  _T_28; // @[Multiplier.scala 125:25]
  wire  _T_29; // @[Multiplier.scala 125:16]
  wire  _T_30; // @[Multiplier.scala 130:39]
  wire  unrolls_less; // @[Multiplier.scala 134:28]
  wire [63:0] unrolls_hi_hi; // @[Multiplier.scala 135:14]
  wire  unrolls_lo; // @[Multiplier.scala 135:67]
  wire [128:0] unrolls_0; // @[Cat.scala 30:58]
  wire  _T_31; // @[Multiplier.scala 139:17]
  wire  _divby0_T; // @[Multiplier.scala 147:24]
  wire  divby0; // @[Multiplier.scala 147:30]
  wire [31:0] divisorMSB_hi; // @[CircuitMath.scala 35:17]
  wire [31:0] divisorMSB_lo; // @[CircuitMath.scala 36:17]
  wire  divisorMSB_hi_1; // @[CircuitMath.scala 37:22]
  wire [15:0] divisorMSB_hi_2; // @[CircuitMath.scala 35:17]
  wire [15:0] divisorMSB_lo_1; // @[CircuitMath.scala 36:17]
  wire  divisorMSB_hi_3; // @[CircuitMath.scala 37:22]
  wire [7:0] divisorMSB_hi_4; // @[CircuitMath.scala 35:17]
  wire [7:0] divisorMSB_lo_2; // @[CircuitMath.scala 36:17]
  wire  divisorMSB_hi_5; // @[CircuitMath.scala 37:22]
  wire [3:0] divisorMSB_hi_6; // @[CircuitMath.scala 35:17]
  wire [3:0] divisorMSB_lo_3; // @[CircuitMath.scala 36:17]
  wire  divisorMSB_hi_7; // @[CircuitMath.scala 37:22]
  wire [1:0] _divisorMSB_T_4; // @[CircuitMath.scala 32:10]
  wire [1:0] _divisorMSB_T_5; // @[CircuitMath.scala 32:10]
  wire [1:0] _divisorMSB_T_9; // @[CircuitMath.scala 32:10]
  wire [1:0] _divisorMSB_T_10; // @[CircuitMath.scala 32:10]
  wire [1:0] divisorMSB_lo_4; // @[CircuitMath.scala 38:21]
  wire [2:0] _divisorMSB_T_11; // @[Cat.scala 30:58]
  wire [3:0] divisorMSB_hi_8; // @[CircuitMath.scala 35:17]
  wire [3:0] divisorMSB_lo_5; // @[CircuitMath.scala 36:17]
  wire  divisorMSB_hi_9; // @[CircuitMath.scala 37:22]
  wire [1:0] _divisorMSB_T_15; // @[CircuitMath.scala 32:10]
  wire [1:0] _divisorMSB_T_16; // @[CircuitMath.scala 32:10]
  wire [1:0] _divisorMSB_T_20; // @[CircuitMath.scala 32:10]
  wire [1:0] _divisorMSB_T_21; // @[CircuitMath.scala 32:10]
  wire [1:0] divisorMSB_lo_6; // @[CircuitMath.scala 38:21]
  wire [2:0] _divisorMSB_T_22; // @[Cat.scala 30:58]
  wire [2:0] divisorMSB_lo_7; // @[CircuitMath.scala 38:21]
  wire [3:0] _divisorMSB_T_23; // @[Cat.scala 30:58]
  wire [7:0] divisorMSB_hi_10; // @[CircuitMath.scala 35:17]
  wire [7:0] divisorMSB_lo_8; // @[CircuitMath.scala 36:17]
  wire  divisorMSB_hi_11; // @[CircuitMath.scala 37:22]
  wire [3:0] divisorMSB_hi_12; // @[CircuitMath.scala 35:17]
  wire [3:0] divisorMSB_lo_9; // @[CircuitMath.scala 36:17]
  wire  divisorMSB_hi_13; // @[CircuitMath.scala 37:22]
  wire [1:0] _divisorMSB_T_27; // @[CircuitMath.scala 32:10]
  wire [1:0] _divisorMSB_T_28; // @[CircuitMath.scala 32:10]
  wire [1:0] _divisorMSB_T_32; // @[CircuitMath.scala 32:10]
  wire [1:0] _divisorMSB_T_33; // @[CircuitMath.scala 32:10]
  wire [1:0] divisorMSB_lo_10; // @[CircuitMath.scala 38:21]
  wire [2:0] _divisorMSB_T_34; // @[Cat.scala 30:58]
  wire [3:0] divisorMSB_hi_14; // @[CircuitMath.scala 35:17]
  wire [3:0] divisorMSB_lo_11; // @[CircuitMath.scala 36:17]
  wire  divisorMSB_hi_15; // @[CircuitMath.scala 37:22]
  wire [1:0] _divisorMSB_T_38; // @[CircuitMath.scala 32:10]
  wire [1:0] _divisorMSB_T_39; // @[CircuitMath.scala 32:10]
  wire [1:0] _divisorMSB_T_43; // @[CircuitMath.scala 32:10]
  wire [1:0] _divisorMSB_T_44; // @[CircuitMath.scala 32:10]
  wire [1:0] divisorMSB_lo_12; // @[CircuitMath.scala 38:21]
  wire [2:0] _divisorMSB_T_45; // @[Cat.scala 30:58]
  wire [2:0] divisorMSB_lo_13; // @[CircuitMath.scala 38:21]
  wire [3:0] _divisorMSB_T_46; // @[Cat.scala 30:58]
  wire [3:0] divisorMSB_lo_14; // @[CircuitMath.scala 38:21]
  wire [4:0] _divisorMSB_T_47; // @[Cat.scala 30:58]
  wire [15:0] divisorMSB_hi_16; // @[CircuitMath.scala 35:17]
  wire [15:0] divisorMSB_lo_15; // @[CircuitMath.scala 36:17]
  wire  divisorMSB_hi_17; // @[CircuitMath.scala 37:22]
  wire [7:0] divisorMSB_hi_18; // @[CircuitMath.scala 35:17]
  wire [7:0] divisorMSB_lo_16; // @[CircuitMath.scala 36:17]
  wire  divisorMSB_hi_19; // @[CircuitMath.scala 37:22]
  wire [3:0] divisorMSB_hi_20; // @[CircuitMath.scala 35:17]
  wire [3:0] divisorMSB_lo_17; // @[CircuitMath.scala 36:17]
  wire  divisorMSB_hi_21; // @[CircuitMath.scala 37:22]
  wire [1:0] _divisorMSB_T_51; // @[CircuitMath.scala 32:10]
  wire [1:0] _divisorMSB_T_52; // @[CircuitMath.scala 32:10]
  wire [1:0] _divisorMSB_T_56; // @[CircuitMath.scala 32:10]
  wire [1:0] _divisorMSB_T_57; // @[CircuitMath.scala 32:10]
  wire [1:0] divisorMSB_lo_18; // @[CircuitMath.scala 38:21]
  wire [2:0] _divisorMSB_T_58; // @[Cat.scala 30:58]
  wire [3:0] divisorMSB_hi_22; // @[CircuitMath.scala 35:17]
  wire [3:0] divisorMSB_lo_19; // @[CircuitMath.scala 36:17]
  wire  divisorMSB_hi_23; // @[CircuitMath.scala 37:22]
  wire [1:0] _divisorMSB_T_62; // @[CircuitMath.scala 32:10]
  wire [1:0] _divisorMSB_T_63; // @[CircuitMath.scala 32:10]
  wire [1:0] _divisorMSB_T_67; // @[CircuitMath.scala 32:10]
  wire [1:0] _divisorMSB_T_68; // @[CircuitMath.scala 32:10]
  wire [1:0] divisorMSB_lo_20; // @[CircuitMath.scala 38:21]
  wire [2:0] _divisorMSB_T_69; // @[Cat.scala 30:58]
  wire [2:0] divisorMSB_lo_21; // @[CircuitMath.scala 38:21]
  wire [3:0] _divisorMSB_T_70; // @[Cat.scala 30:58]
  wire [7:0] divisorMSB_hi_24; // @[CircuitMath.scala 35:17]
  wire [7:0] divisorMSB_lo_22; // @[CircuitMath.scala 36:17]
  wire  divisorMSB_hi_25; // @[CircuitMath.scala 37:22]
  wire [3:0] divisorMSB_hi_26; // @[CircuitMath.scala 35:17]
  wire [3:0] divisorMSB_lo_23; // @[CircuitMath.scala 36:17]
  wire  divisorMSB_hi_27; // @[CircuitMath.scala 37:22]
  wire [1:0] _divisorMSB_T_74; // @[CircuitMath.scala 32:10]
  wire [1:0] _divisorMSB_T_75; // @[CircuitMath.scala 32:10]
  wire [1:0] _divisorMSB_T_79; // @[CircuitMath.scala 32:10]
  wire [1:0] _divisorMSB_T_80; // @[CircuitMath.scala 32:10]
  wire [1:0] divisorMSB_lo_24; // @[CircuitMath.scala 38:21]
  wire [2:0] _divisorMSB_T_81; // @[Cat.scala 30:58]
  wire [3:0] divisorMSB_hi_28; // @[CircuitMath.scala 35:17]
  wire [3:0] divisorMSB_lo_25; // @[CircuitMath.scala 36:17]
  wire  divisorMSB_hi_29; // @[CircuitMath.scala 37:22]
  wire [1:0] _divisorMSB_T_85; // @[CircuitMath.scala 32:10]
  wire [1:0] _divisorMSB_T_86; // @[CircuitMath.scala 32:10]
  wire [1:0] _divisorMSB_T_90; // @[CircuitMath.scala 32:10]
  wire [1:0] _divisorMSB_T_91; // @[CircuitMath.scala 32:10]
  wire [1:0] divisorMSB_lo_26; // @[CircuitMath.scala 38:21]
  wire [2:0] _divisorMSB_T_92; // @[Cat.scala 30:58]
  wire [2:0] divisorMSB_lo_27; // @[CircuitMath.scala 38:21]
  wire [3:0] _divisorMSB_T_93; // @[Cat.scala 30:58]
  wire [3:0] divisorMSB_lo_28; // @[CircuitMath.scala 38:21]
  wire [4:0] _divisorMSB_T_94; // @[Cat.scala 30:58]
  wire [4:0] divisorMSB_lo_29; // @[CircuitMath.scala 38:21]
  wire [5:0] divisorMSB; // @[Cat.scala 30:58]
  wire [31:0] dividendMSB_hi; // @[CircuitMath.scala 35:17]
  wire [31:0] dividendMSB_lo; // @[CircuitMath.scala 36:17]
  wire  dividendMSB_hi_1; // @[CircuitMath.scala 37:22]
  wire [15:0] dividendMSB_hi_2; // @[CircuitMath.scala 35:17]
  wire [15:0] dividendMSB_lo_1; // @[CircuitMath.scala 36:17]
  wire  dividendMSB_hi_3; // @[CircuitMath.scala 37:22]
  wire [7:0] dividendMSB_hi_4; // @[CircuitMath.scala 35:17]
  wire [7:0] dividendMSB_lo_2; // @[CircuitMath.scala 36:17]
  wire  dividendMSB_hi_5; // @[CircuitMath.scala 37:22]
  wire [3:0] dividendMSB_hi_6; // @[CircuitMath.scala 35:17]
  wire [3:0] dividendMSB_lo_3; // @[CircuitMath.scala 36:17]
  wire  dividendMSB_hi_7; // @[CircuitMath.scala 37:22]
  wire [1:0] _dividendMSB_T_4; // @[CircuitMath.scala 32:10]
  wire [1:0] _dividendMSB_T_5; // @[CircuitMath.scala 32:10]
  wire [1:0] _dividendMSB_T_9; // @[CircuitMath.scala 32:10]
  wire [1:0] _dividendMSB_T_10; // @[CircuitMath.scala 32:10]
  wire [1:0] dividendMSB_lo_4; // @[CircuitMath.scala 38:21]
  wire [2:0] _dividendMSB_T_11; // @[Cat.scala 30:58]
  wire [3:0] dividendMSB_hi_8; // @[CircuitMath.scala 35:17]
  wire [3:0] dividendMSB_lo_5; // @[CircuitMath.scala 36:17]
  wire  dividendMSB_hi_9; // @[CircuitMath.scala 37:22]
  wire [1:0] _dividendMSB_T_15; // @[CircuitMath.scala 32:10]
  wire [1:0] _dividendMSB_T_16; // @[CircuitMath.scala 32:10]
  wire [1:0] _dividendMSB_T_20; // @[CircuitMath.scala 32:10]
  wire [1:0] _dividendMSB_T_21; // @[CircuitMath.scala 32:10]
  wire [1:0] dividendMSB_lo_6; // @[CircuitMath.scala 38:21]
  wire [2:0] _dividendMSB_T_22; // @[Cat.scala 30:58]
  wire [2:0] dividendMSB_lo_7; // @[CircuitMath.scala 38:21]
  wire [3:0] _dividendMSB_T_23; // @[Cat.scala 30:58]
  wire [7:0] dividendMSB_hi_10; // @[CircuitMath.scala 35:17]
  wire [7:0] dividendMSB_lo_8; // @[CircuitMath.scala 36:17]
  wire  dividendMSB_hi_11; // @[CircuitMath.scala 37:22]
  wire [3:0] dividendMSB_hi_12; // @[CircuitMath.scala 35:17]
  wire [3:0] dividendMSB_lo_9; // @[CircuitMath.scala 36:17]
  wire  dividendMSB_hi_13; // @[CircuitMath.scala 37:22]
  wire [1:0] _dividendMSB_T_27; // @[CircuitMath.scala 32:10]
  wire [1:0] _dividendMSB_T_28; // @[CircuitMath.scala 32:10]
  wire [1:0] _dividendMSB_T_32; // @[CircuitMath.scala 32:10]
  wire [1:0] _dividendMSB_T_33; // @[CircuitMath.scala 32:10]
  wire [1:0] dividendMSB_lo_10; // @[CircuitMath.scala 38:21]
  wire [2:0] _dividendMSB_T_34; // @[Cat.scala 30:58]
  wire [3:0] dividendMSB_hi_14; // @[CircuitMath.scala 35:17]
  wire [3:0] dividendMSB_lo_11; // @[CircuitMath.scala 36:17]
  wire  dividendMSB_hi_15; // @[CircuitMath.scala 37:22]
  wire [1:0] _dividendMSB_T_38; // @[CircuitMath.scala 32:10]
  wire [1:0] _dividendMSB_T_39; // @[CircuitMath.scala 32:10]
  wire [1:0] _dividendMSB_T_43; // @[CircuitMath.scala 32:10]
  wire [1:0] _dividendMSB_T_44; // @[CircuitMath.scala 32:10]
  wire [1:0] dividendMSB_lo_12; // @[CircuitMath.scala 38:21]
  wire [2:0] _dividendMSB_T_45; // @[Cat.scala 30:58]
  wire [2:0] dividendMSB_lo_13; // @[CircuitMath.scala 38:21]
  wire [3:0] _dividendMSB_T_46; // @[Cat.scala 30:58]
  wire [3:0] dividendMSB_lo_14; // @[CircuitMath.scala 38:21]
  wire [4:0] _dividendMSB_T_47; // @[Cat.scala 30:58]
  wire [15:0] dividendMSB_hi_16; // @[CircuitMath.scala 35:17]
  wire [15:0] dividendMSB_lo_15; // @[CircuitMath.scala 36:17]
  wire  dividendMSB_hi_17; // @[CircuitMath.scala 37:22]
  wire [7:0] dividendMSB_hi_18; // @[CircuitMath.scala 35:17]
  wire [7:0] dividendMSB_lo_16; // @[CircuitMath.scala 36:17]
  wire  dividendMSB_hi_19; // @[CircuitMath.scala 37:22]
  wire [3:0] dividendMSB_hi_20; // @[CircuitMath.scala 35:17]
  wire [3:0] dividendMSB_lo_17; // @[CircuitMath.scala 36:17]
  wire  dividendMSB_hi_21; // @[CircuitMath.scala 37:22]
  wire [1:0] _dividendMSB_T_51; // @[CircuitMath.scala 32:10]
  wire [1:0] _dividendMSB_T_52; // @[CircuitMath.scala 32:10]
  wire [1:0] _dividendMSB_T_56; // @[CircuitMath.scala 32:10]
  wire [1:0] _dividendMSB_T_57; // @[CircuitMath.scala 32:10]
  wire [1:0] dividendMSB_lo_18; // @[CircuitMath.scala 38:21]
  wire [2:0] _dividendMSB_T_58; // @[Cat.scala 30:58]
  wire [3:0] dividendMSB_hi_22; // @[CircuitMath.scala 35:17]
  wire [3:0] dividendMSB_lo_19; // @[CircuitMath.scala 36:17]
  wire  dividendMSB_hi_23; // @[CircuitMath.scala 37:22]
  wire [1:0] _dividendMSB_T_62; // @[CircuitMath.scala 32:10]
  wire [1:0] _dividendMSB_T_63; // @[CircuitMath.scala 32:10]
  wire [1:0] _dividendMSB_T_67; // @[CircuitMath.scala 32:10]
  wire [1:0] _dividendMSB_T_68; // @[CircuitMath.scala 32:10]
  wire [1:0] dividendMSB_lo_20; // @[CircuitMath.scala 38:21]
  wire [2:0] _dividendMSB_T_69; // @[Cat.scala 30:58]
  wire [2:0] dividendMSB_lo_21; // @[CircuitMath.scala 38:21]
  wire [3:0] _dividendMSB_T_70; // @[Cat.scala 30:58]
  wire [7:0] dividendMSB_hi_24; // @[CircuitMath.scala 35:17]
  wire [7:0] dividendMSB_lo_22; // @[CircuitMath.scala 36:17]
  wire  dividendMSB_hi_25; // @[CircuitMath.scala 37:22]
  wire [3:0] dividendMSB_hi_26; // @[CircuitMath.scala 35:17]
  wire [3:0] dividendMSB_lo_23; // @[CircuitMath.scala 36:17]
  wire  dividendMSB_hi_27; // @[CircuitMath.scala 37:22]
  wire [1:0] _dividendMSB_T_74; // @[CircuitMath.scala 32:10]
  wire [1:0] _dividendMSB_T_75; // @[CircuitMath.scala 32:10]
  wire [1:0] _dividendMSB_T_79; // @[CircuitMath.scala 32:10]
  wire [1:0] _dividendMSB_T_80; // @[CircuitMath.scala 32:10]
  wire [1:0] dividendMSB_lo_24; // @[CircuitMath.scala 38:21]
  wire [2:0] _dividendMSB_T_81; // @[Cat.scala 30:58]
  wire [3:0] dividendMSB_hi_28; // @[CircuitMath.scala 35:17]
  wire [3:0] dividendMSB_lo_25; // @[CircuitMath.scala 36:17]
  wire  dividendMSB_hi_29; // @[CircuitMath.scala 37:22]
  wire [1:0] _dividendMSB_T_85; // @[CircuitMath.scala 32:10]
  wire [1:0] _dividendMSB_T_86; // @[CircuitMath.scala 32:10]
  wire [1:0] _dividendMSB_T_90; // @[CircuitMath.scala 32:10]
  wire [1:0] _dividendMSB_T_91; // @[CircuitMath.scala 32:10]
  wire [1:0] dividendMSB_lo_26; // @[CircuitMath.scala 38:21]
  wire [2:0] _dividendMSB_T_92; // @[Cat.scala 30:58]
  wire [2:0] dividendMSB_lo_27; // @[CircuitMath.scala 38:21]
  wire [3:0] _dividendMSB_T_93; // @[Cat.scala 30:58]
  wire [3:0] dividendMSB_lo_28; // @[CircuitMath.scala 38:21]
  wire [4:0] _dividendMSB_T_94; // @[Cat.scala 30:58]
  wire [4:0] dividendMSB_lo_29; // @[CircuitMath.scala 38:21]
  wire [5:0] dividendMSB; // @[Cat.scala 30:58]
  wire [5:0] _eOutPos_T_1; // @[Multiplier.scala 153:35]
  wire [5:0] eOutPos; // @[Multiplier.scala 153:21]
  wire  _eOut_T_11; // @[Multiplier.scala 154:30]
  wire  _eOut_T_12; // @[Multiplier.scala 154:52]
  wire  eOut_1; // @[Multiplier.scala 154:41]
  wire [126:0] _GEN_39; // @[Multiplier.scala 156:39]
  wire [126:0] _remainder_T_2; // @[Multiplier.scala 156:39]
  wire [128:0] _GEN_16; // @[Multiplier.scala 155:19]
  wire  _T_33; // @[Multiplier.scala 160:18]
  wire  _T_34; // @[Decoupled.scala 40:37]
  wire  _T_35; // @[Multiplier.scala 162:24]
  wire  _T_36; // @[Decoupled.scala 40:37]
  wire  _state_T_1; // @[Multiplier.scala 166:46]
  wire  _count_T_7; // @[Multiplier.scala 169:46]
  wire [2:0] _count_T_8; // @[Multiplier.scala 169:38]
  wire  _neg_out_T; // @[Multiplier.scala 170:46]
  wire [64:0] _divisor_T; // @[Cat.scala 30:58]
  wire [2:0] _outMul_T_1; // @[Multiplier.scala 176:23]
  wire  outMul; // @[Multiplier.scala 176:52]
  wire  _loOut_T_3; // @[Multiplier.scala 177:48]
  wire [31:0] loOut; // @[Multiplier.scala 177:18]
  wire [31:0] _hiOut_T_4; // @[Bitwise.scala 72:12]
  wire [31:0] hiOut; // @[Multiplier.scala 178:18]
  wire  _io_resp_valid_T; // @[Multiplier.scala 182:27]
  wire  _io_resp_valid_T_1; // @[Multiplier.scala 182:51]
  reg [19:0] MulDiv_state; // @[Register tracking MulDiv state]
  reg [31:0] _RAND_9;
  reg  MulDiv_cov [0:1048575]; // @[Coverage map for MulDiv]
  reg [31:0] _RAND_10;
  wire  MulDiv_cov_read_data; // @[Coverage map for MulDiv]
  wire [19:0] MulDiv_cov_read_addr; // @[Coverage map for MulDiv]
  wire  MulDiv_cov_write_data; // @[Coverage map for MulDiv]
  wire [19:0] MulDiv_cov_write_addr; // @[Coverage map for MulDiv]
  wire  MulDiv_cov_write_mask; // @[Coverage map for MulDiv]
  wire  MulDiv_cov_write_en; // @[Coverage map for MulDiv]
  reg [29:0] MulDiv_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_11;
  wire  mux_cond_0;
  wire  mux_cond_1;
  wire  mux_cond_2;
  wire  mux_cond_3;
  wire  mux_cond_4;
  wire  mux_cond_5;
  wire  mux_cond_6;
  wire  mux_cond_7;
  wire  mux_cond_8;
  wire  mux_cond_9;
  wire  mux_cond_10;
  wire  mux_cond_11;
  wire  mux_cond_12;
  wire  mux_cond_13;
  wire  mux_cond_14;
  wire  mux_cond_15;
  wire  mux_cond_16;
  wire  mux_cond_17;
  wire  mux_cond_18;
  wire  mux_cond_19;
  wire  mux_cond_20;
  wire  mux_cond_21;
  wire  mux_cond_22;
  wire  mux_cond_23;
  wire  mux_cond_24;
  wire  mux_cond_25;
  wire  mux_cond_26;
  wire  mux_cond_27;
  wire  mux_cond_28;
  wire  mux_cond_29;
  wire  mux_cond_30;
  wire  mux_cond_31;
  wire  mux_cond_32;
  wire  mux_cond_33;
  wire  mux_cond_34;
  wire  mux_cond_35;
  wire  mux_cond_36;
  wire  mux_cond_37;
  wire  mux_cond_38;
  wire  mux_cond_39;
  wire  mux_cond_40;
  wire  mux_cond_41;
  wire  mux_cond_42;
  wire  mux_cond_43;
  wire  mux_cond_44;
  wire  mux_cond_45;
  wire  mux_cond_46;
  wire  mux_cond_47;
  wire  mux_cond_48;
  wire  mux_cond_49;
  wire  mux_cond_50;
  wire  mux_cond_51;
  wire  mux_cond_52;
  wire  mux_cond_53;
  wire  mux_cond_54;
  wire  mux_cond_55;
  wire  mux_cond_56;
  wire  mux_cond_57;
  wire  mux_cond_58;
  wire  mux_cond_59;
  wire  mux_cond_60;
  wire  mux_cond_61;
  wire  mux_cond_62;
  wire  mux_cond_63;
  wire  mux_cond_64;
  wire  mux_cond_65;
  wire  mux_cond_66;
  wire  mux_cond_67;
  wire  mux_cond_68;
  wire  mux_cond_69;
  wire  mux_cond_70;
  wire  mux_cond_71;
  wire  mux_cond_72;
  wire  mux_cond_73;
  wire  mux_cond_74;
  wire  mux_cond_75;
  wire  mux_cond_76;
  wire  mux_cond_77;
  wire  mux_cond_78;
  wire  mux_cond_79;
  wire  mux_cond_80;
  wire  mux_cond_81;
  wire  mux_cond_82;
  wire  mux_cond_83;
  wire  mux_cond_84;
  wire  mux_cond_85;
  wire  mux_cond_86;
  wire  mux_cond_87;
  wire  mux_cond_88;
  wire  mux_cond_89;
  wire  mux_cond_90;
  wire  mux_cond_91;
  wire  mux_cond_92;
  wire  mux_cond_93;
  wire  mux_cond_94;
  wire  mux_cond_95;
  wire  mux_cond_96;
  wire  mux_cond_97;
  wire [4:0] isHi_shl;
  wire [19:0] isHi_pad;
  wire [12:0] neg_out_shl;
  wire [19:0] neg_out_pad;
  wire [4:0] req_dw_shl;
  wire [19:0] req_dw_pad;
  wire [10:0] state_shl;
  wire [19:0] state_pad;
  wire [1:0] resHi_shl;
  wire [19:0] resHi_pad;
  wire [12:0] mux_cond_0_shl;
  wire [19:0] mux_cond_0_pad;
  wire [1:0] mux_cond_1_shl;
  wire [19:0] mux_cond_1_pad;
  wire  mux_cond_2_shl;
  wire [19:0] mux_cond_2_pad;
  wire [12:0] mux_cond_3_shl;
  wire [19:0] mux_cond_3_pad;
  wire [15:0] mux_cond_4_shl;
  wire [19:0] mux_cond_4_pad;
  wire [11:0] mux_cond_5_shl;
  wire [19:0] mux_cond_5_pad;
  wire [7:0] mux_cond_6_shl;
  wire [19:0] mux_cond_6_pad;
  wire [17:0] mux_cond_7_shl;
  wire [19:0] mux_cond_7_pad;
  wire [11:0] mux_cond_8_shl;
  wire [19:0] mux_cond_8_pad;
  wire [15:0] mux_cond_9_shl;
  wire [19:0] mux_cond_9_pad;
  wire [13:0] mux_cond_10_shl;
  wire [19:0] mux_cond_10_pad;
  wire  mux_cond_11_shl;
  wire [19:0] mux_cond_11_pad;
  wire [7:0] mux_cond_12_shl;
  wire [19:0] mux_cond_12_pad;
  wire [13:0] mux_cond_13_shl;
  wire [19:0] mux_cond_13_pad;
  wire  mux_cond_14_shl;
  wire [19:0] mux_cond_14_pad;
  wire [9:0] mux_cond_15_shl;
  wire [19:0] mux_cond_15_pad;
  wire [8:0] mux_cond_16_shl;
  wire [19:0] mux_cond_16_pad;
  wire [8:0] mux_cond_17_shl;
  wire [19:0] mux_cond_17_pad;
  wire [8:0] mux_cond_18_shl;
  wire [19:0] mux_cond_18_pad;
  wire [2:0] mux_cond_19_shl;
  wire [19:0] mux_cond_19_pad;
  wire [16:0] mux_cond_20_shl;
  wire [19:0] mux_cond_20_pad;
  wire [6:0] mux_cond_21_shl;
  wire [19:0] mux_cond_21_pad;
  wire [11:0] mux_cond_22_shl;
  wire [19:0] mux_cond_22_pad;
  wire  mux_cond_23_shl;
  wire [19:0] mux_cond_23_pad;
  wire [6:0] mux_cond_24_shl;
  wire [19:0] mux_cond_24_pad;
  wire [12:0] mux_cond_25_shl;
  wire [19:0] mux_cond_25_pad;
  wire [4:0] mux_cond_26_shl;
  wire [19:0] mux_cond_26_pad;
  wire [11:0] mux_cond_27_shl;
  wire [19:0] mux_cond_27_pad;
  wire [6:0] mux_cond_28_shl;
  wire [19:0] mux_cond_28_pad;
  wire [12:0] mux_cond_29_shl;
  wire [19:0] mux_cond_29_pad;
  wire [1:0] mux_cond_30_shl;
  wire [19:0] mux_cond_30_pad;
  wire [11:0] mux_cond_31_shl;
  wire [19:0] mux_cond_31_pad;
  wire [6:0] mux_cond_32_shl;
  wire [19:0] mux_cond_32_pad;
  wire [5:0] mux_cond_33_shl;
  wire [19:0] mux_cond_33_pad;
  wire [18:0] mux_cond_34_shl;
  wire [19:0] mux_cond_34_pad;
  wire [12:0] mux_cond_35_shl;
  wire [19:0] mux_cond_35_pad;
  wire  mux_cond_36_shl;
  wire [19:0] mux_cond_36_pad;
  wire [8:0] mux_cond_37_shl;
  wire [19:0] mux_cond_37_pad;
  wire [5:0] mux_cond_38_shl;
  wire [19:0] mux_cond_38_pad;
  wire [16:0] mux_cond_39_shl;
  wire [19:0] mux_cond_39_pad;
  wire [3:0] mux_cond_40_shl;
  wire [19:0] mux_cond_40_pad;
  wire [9:0] mux_cond_41_shl;
  wire [19:0] mux_cond_41_pad;
  wire [15:0] mux_cond_42_shl;
  wire [19:0] mux_cond_42_pad;
  wire [13:0] mux_cond_43_shl;
  wire [19:0] mux_cond_43_pad;
  wire [12:0] mux_cond_44_shl;
  wire [19:0] mux_cond_44_pad;
  wire  mux_cond_45_shl;
  wire [19:0] mux_cond_45_pad;
  wire [3:0] mux_cond_46_shl;
  wire [19:0] mux_cond_46_pad;
  wire [14:0] mux_cond_47_shl;
  wire [19:0] mux_cond_47_pad;
  wire [16:0] mux_cond_48_shl;
  wire [19:0] mux_cond_48_pad;
  wire [18:0] mux_cond_49_shl;
  wire [19:0] mux_cond_49_pad;
  wire  mux_cond_50_shl;
  wire [19:0] mux_cond_50_pad;
  wire [7:0] mux_cond_51_shl;
  wire [19:0] mux_cond_51_pad;
  wire  mux_cond_52_shl;
  wire [19:0] mux_cond_52_pad;
  wire [19:0] mux_cond_53_shl;
  wire [19:0] mux_cond_53_pad;
  wire [10:0] mux_cond_54_shl;
  wire [19:0] mux_cond_54_pad;
  wire [13:0] mux_cond_55_shl;
  wire [19:0] mux_cond_55_pad;
  wire [9:0] mux_cond_56_shl;
  wire [19:0] mux_cond_56_pad;
  wire [6:0] mux_cond_57_shl;
  wire [19:0] mux_cond_57_pad;
  wire [17:0] mux_cond_58_shl;
  wire [19:0] mux_cond_58_pad;
  wire [19:0] mux_cond_59_shl;
  wire [19:0] mux_cond_59_pad;
  wire [3:0] mux_cond_60_shl;
  wire [19:0] mux_cond_60_pad;
  wire [14:0] mux_cond_61_shl;
  wire [19:0] mux_cond_61_pad;
  wire [4:0] mux_cond_62_shl;
  wire [19:0] mux_cond_62_pad;
  wire  mux_cond_63_shl;
  wire [19:0] mux_cond_63_pad;
  wire [10:0] mux_cond_64_shl;
  wire [19:0] mux_cond_64_pad;
  wire [17:0] mux_cond_65_shl;
  wire [19:0] mux_cond_65_pad;
  wire [9:0] mux_cond_66_shl;
  wire [19:0] mux_cond_66_pad;
  wire [6:0] mux_cond_67_shl;
  wire [19:0] mux_cond_67_pad;
  wire [19:0] mux_cond_68_shl;
  wire [19:0] mux_cond_68_pad;
  wire [10:0] mux_cond_69_shl;
  wire [19:0] mux_cond_69_pad;
  wire [10:0] mux_cond_70_shl;
  wire [19:0] mux_cond_70_pad;
  wire [13:0] mux_cond_71_shl;
  wire [19:0] mux_cond_71_pad;
  wire [18:0] mux_cond_72_shl;
  wire [19:0] mux_cond_72_pad;
  wire [12:0] mux_cond_73_shl;
  wire [19:0] mux_cond_73_pad;
  wire [13:0] mux_cond_74_shl;
  wire [19:0] mux_cond_74_pad;
  wire [13:0] mux_cond_75_shl;
  wire [19:0] mux_cond_75_pad;
  wire [13:0] mux_cond_76_shl;
  wire [19:0] mux_cond_76_pad;
  wire [13:0] mux_cond_77_shl;
  wire [19:0] mux_cond_77_pad;
  wire [17:0] mux_cond_78_shl;
  wire [19:0] mux_cond_78_pad;
  wire [12:0] mux_cond_79_shl;
  wire [19:0] mux_cond_79_pad;
  wire [17:0] mux_cond_80_shl;
  wire [19:0] mux_cond_80_pad;
  wire [13:0] mux_cond_81_shl;
  wire [19:0] mux_cond_81_pad;
  wire [12:0] mux_cond_82_shl;
  wire [19:0] mux_cond_82_pad;
  wire [4:0] mux_cond_83_shl;
  wire [19:0] mux_cond_83_pad;
  wire [16:0] mux_cond_84_shl;
  wire [19:0] mux_cond_84_pad;
  wire [9:0] mux_cond_85_shl;
  wire [19:0] mux_cond_85_pad;
  wire [10:0] mux_cond_86_shl;
  wire [19:0] mux_cond_86_pad;
  wire [2:0] mux_cond_87_shl;
  wire [19:0] mux_cond_87_pad;
  wire [6:0] mux_cond_88_shl;
  wire [19:0] mux_cond_88_pad;
  wire [11:0] mux_cond_89_shl;
  wire [19:0] mux_cond_89_pad;
  wire [7:0] mux_cond_90_shl;
  wire [19:0] mux_cond_90_pad;
  wire [16:0] mux_cond_91_shl;
  wire [19:0] mux_cond_91_pad;
  wire [17:0] mux_cond_92_shl;
  wire [19:0] mux_cond_92_pad;
  wire [5:0] mux_cond_93_shl;
  wire [19:0] mux_cond_93_pad;
  wire [18:0] mux_cond_94_shl;
  wire [19:0] mux_cond_94_pad;
  wire [1:0] mux_cond_95_shl;
  wire [19:0] mux_cond_95_pad;
  wire [17:0] mux_cond_96_shl;
  wire [19:0] mux_cond_96_pad;
  wire [1:0] mux_cond_97_shl;
  wire [19:0] mux_cond_97_pad;
  wire [19:0] MulDiv_xor64;
  wire [19:0] MulDiv_xor31;
  wire [19:0] MulDiv_xor66;
  wire [19:0] MulDiv_xor32;
  wire [19:0] MulDiv_xor15;
  wire [19:0] MulDiv_xor68;
  wire [19:0] MulDiv_xor33;
  wire [19:0] MulDiv_xor70;
  wire [19:0] MulDiv_xor34;
  wire [19:0] MulDiv_xor16;
  wire [19:0] MulDiv_xor7;
  wire [19:0] MulDiv_xor72;
  wire [19:0] MulDiv_xor35;
  wire [19:0] MulDiv_xor74;
  wire [19:0] MulDiv_xor36;
  wire [19:0] MulDiv_xor17;
  wire [19:0] MulDiv_xor76;
  wire [19:0] MulDiv_xor37;
  wire [19:0] MulDiv_xor77;
  wire [19:0] MulDiv_xor78;
  wire [19:0] MulDiv_xor38;
  wire [19:0] MulDiv_xor18;
  wire [19:0] MulDiv_xor8;
  wire [19:0] MulDiv_xor3;
  wire [19:0] MulDiv_xor80;
  wire [19:0] MulDiv_xor39;
  wire [19:0] MulDiv_xor82;
  wire [19:0] MulDiv_xor40;
  wire [19:0] MulDiv_xor19;
  wire [19:0] MulDiv_xor84;
  wire [19:0] MulDiv_xor41;
  wire [19:0] MulDiv_xor85;
  wire [19:0] MulDiv_xor86;
  wire [19:0] MulDiv_xor42;
  wire [19:0] MulDiv_xor20;
  wire [19:0] MulDiv_xor9;
  wire [19:0] MulDiv_xor88;
  wire [19:0] MulDiv_xor43;
  wire [19:0] MulDiv_xor90;
  wire [19:0] MulDiv_xor44;
  wire [19:0] MulDiv_xor21;
  wire [19:0] MulDiv_xor92;
  wire [19:0] MulDiv_xor45;
  wire [19:0] MulDiv_xor93;
  wire [19:0] MulDiv_xor94;
  wire [19:0] MulDiv_xor46;
  wire [19:0] MulDiv_xor22;
  wire [19:0] MulDiv_xor10;
  wire [19:0] MulDiv_xor4;
  wire [19:0] MulDiv_xor1;
  wire [19:0] MulDiv_xor96;
  wire [19:0] MulDiv_xor47;
  wire [19:0] MulDiv_xor98;
  wire [19:0] MulDiv_xor48;
  wire [19:0] MulDiv_xor23;
  wire [19:0] MulDiv_xor100;
  wire [19:0] MulDiv_xor49;
  wire [19:0] MulDiv_xor101;
  wire [19:0] MulDiv_xor102;
  wire [19:0] MulDiv_xor50;
  wire [19:0] MulDiv_xor24;
  wire [19:0] MulDiv_xor11;
  wire [19:0] MulDiv_xor104;
  wire [19:0] MulDiv_xor51;
  wire [19:0] MulDiv_xor106;
  wire [19:0] MulDiv_xor52;
  wire [19:0] MulDiv_xor25;
  wire [19:0] MulDiv_xor108;
  wire [19:0] MulDiv_xor53;
  wire [19:0] MulDiv_xor109;
  wire [19:0] MulDiv_xor110;
  wire [19:0] MulDiv_xor54;
  wire [19:0] MulDiv_xor26;
  wire [19:0] MulDiv_xor12;
  wire [19:0] MulDiv_xor5;
  wire [19:0] MulDiv_xor112;
  wire [19:0] MulDiv_xor55;
  wire [19:0] MulDiv_xor114;
  wire [19:0] MulDiv_xor56;
  wire [19:0] MulDiv_xor27;
  wire [19:0] MulDiv_xor116;
  wire [19:0] MulDiv_xor57;
  wire [19:0] MulDiv_xor117;
  wire [19:0] MulDiv_xor118;
  wire [19:0] MulDiv_xor58;
  wire [19:0] MulDiv_xor28;
  wire [19:0] MulDiv_xor13;
  wire [19:0] MulDiv_xor120;
  wire [19:0] MulDiv_xor59;
  wire [19:0] MulDiv_xor122;
  wire [19:0] MulDiv_xor60;
  wire [19:0] MulDiv_xor29;
  wire [19:0] MulDiv_xor124;
  wire [19:0] MulDiv_xor61;
  wire [19:0] MulDiv_xor125;
  wire [19:0] MulDiv_xor126;
  wire [19:0] MulDiv_xor62;
  wire [19:0] MulDiv_xor30;
  wire [19:0] MulDiv_xor14;
  wire [19:0] MulDiv_xor6;
  wire [19:0] MulDiv_xor2;
  wire [19:0] MulDiv_xor0;
  assign _T = io_req_bits_fn & 4'h4; // @[Decode.scala 14:65]
  assign cmdMul = _T == 4'h0; // @[Decode.scala 14:121]
  assign _T_3 = io_req_bits_fn & 4'h5; // @[Decode.scala 14:65]
  assign _T_4 = _T_3 == 4'h1; // @[Decode.scala 14:121]
  assign _T_5 = io_req_bits_fn & 4'h2; // @[Decode.scala 14:65]
  assign _T_6 = _T_5 == 4'h2; // @[Decode.scala 14:121]
  assign cmdHi = _T_4 | _T_6; // @[Decode.scala 15:30]
  assign _T_9 = io_req_bits_fn & 4'h6; // @[Decode.scala 14:65]
  assign _T_10 = _T_9 == 4'h0; // @[Decode.scala 14:121]
  assign _T_11 = io_req_bits_fn & 4'h1; // @[Decode.scala 14:65]
  assign _T_12 = _T_11 == 4'h0; // @[Decode.scala 14:121]
  assign lhsSigned = _T_10 | _T_12; // @[Decode.scala 15:30]
  assign _T_16 = _T_3 == 4'h4; // @[Decode.scala 14:121]
  assign rhsSigned = _T_10 | _T_16; // @[Decode.scala 15:30]
  assign _sign_T_2 = io_req_bits_dw ? io_req_bits_in1[63] : io_req_bits_in1[31]; // @[Multiplier.scala 82:29]
  assign lhs_sign = lhsSigned & _sign_T_2; // @[Multiplier.scala 82:23]
  assign _hi_T_1 = lhs_sign ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  assign hi = io_req_bits_dw ? io_req_bits_in1[63:32] : _hi_T_1; // @[Multiplier.scala 83:17]
  assign lo = io_req_bits_in1[31:0]; // @[Multiplier.scala 84:15]
  assign lhs_in = {hi,lo}; // @[Cat.scala 30:58]
  assign _sign_T_5 = io_req_bits_dw ? io_req_bits_in2[63] : io_req_bits_in2[31]; // @[Multiplier.scala 82:29]
  assign rhs_sign = rhsSigned & _sign_T_5; // @[Multiplier.scala 82:23]
  assign _hi_T_4 = rhs_sign ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  assign hi_1 = io_req_bits_dw ? io_req_bits_in2[63:32] : _hi_T_4; // @[Multiplier.scala 83:17]
  assign lo_1 = io_req_bits_in2[31:0]; // @[Multiplier.scala 84:15]
  assign subtractor = remainder[128:64] - divisor; // @[Multiplier.scala 89:37]
  assign result = resHi ? remainder[128:65] : remainder[63:0]; // @[Multiplier.scala 90:19]
  assign negated_remainder = 64'h0 - result; // @[Multiplier.scala 91:27]
  assign _T_23 = state == 3'h1; // @[Multiplier.scala 93:39]
  assign _T_26 = state == 3'h5; // @[Multiplier.scala 102:39]
  assign _T_27 = state == 3'h2; // @[Multiplier.scala 107:39]
  assign mulReg_hi = remainder[129:65]; // @[Multiplier.scala 108:31]
  assign mulReg = {mulReg_hi,remainder[63:0]}; // @[Cat.scala 30:58]
  assign prod_hi = remainder[64]; // @[Multiplier.scala 109:31]
  assign mplier = mulReg[63:0]; // @[Multiplier.scala 110:24]
  assign accum = mulReg[128:64]; // @[Multiplier.scala 111:37]
  assign prod_lo = mplier[7:0]; // @[Multiplier.scala 113:38]
  assign _prod_T_1 = {prod_hi,prod_lo}; // @[Multiplier.scala 113:60]
  assign _GEN_37 = {{56{_prod_T_1[8]}},_prod_T_1}; // @[Multiplier.scala 113:67]
  assign _prod_T_2 = $signed(_GEN_37) * $signed(divisor); // @[Multiplier.scala 113:67]
  assign _GEN_38 = {{9{accum[64]}},accum}; // @[Multiplier.scala 113:76]
  assign nextMulReg_lo = mplier[63:8]; // @[Multiplier.scala 114:38]
  assign nextMulReg_hi = $signed(_prod_T_2) + $signed(_GEN_38); // @[Cat.scala 30:58]
  assign nextMulReg = {nextMulReg_hi,nextMulReg_lo}; // @[Cat.scala 30:58]
  assign _nextMplierSign_T = count == 7'h6; // @[Multiplier.scala 115:32]
  assign remainder_hi_lo = _nextMplierSign_T & neg_out; // @[Multiplier.scala 115:57]
  assign _eOutMask_T = count * 7'h8; // @[Multiplier.scala 117:54]
  assign _eOutMask_T_2 = -65'sh10000000000000000 >>> _eOutMask_T[5:0]; // @[Multiplier.scala 117:44]
  assign eOutMask = _eOutMask_T_2[63:0]; // @[Multiplier.scala 117:89]
  assign _eOut_T = count != 7'h7; // @[Multiplier.scala 118:45]
  assign _eOut_T_2 = count != 7'h0; // @[Multiplier.scala 118:79]
  assign _eOut_T_3 = _eOut_T & _eOut_T_2; // @[Multiplier.scala 118:70]
  assign _eOut_T_5 = _eOut_T_3 & ~isHi; // @[Multiplier.scala 118:85]
  assign _eOut_T_7 = mplier & ~eOutMask; // @[Multiplier.scala 119:24]
  assign _eOut_T_8 = _eOut_T_7 == 64'h0; // @[Multiplier.scala 119:37]
  assign eOut = _eOut_T_5 & _eOut_T_8; // @[Multiplier.scala 119:13]
  assign _eOutRes_T_2 = 11'h40 - _eOutMask_T; // @[Multiplier.scala 120:36]
  assign eOutRes = mulReg >> _eOutRes_T_2[5:0]; // @[Multiplier.scala 120:27]
  assign nextMulReg1_hi = nextMulReg[128:64]; // @[Multiplier.scala 121:37]
  assign _nextMulReg1_T = eOut ? {{1'd0}, eOutRes} : nextMulReg; // @[Multiplier.scala 121:55]
  assign nextMulReg1_lo = _nextMulReg1_T[63:0]; // @[Multiplier.scala 121:82]
  assign nextMulReg1 = {nextMulReg1_hi,nextMulReg1_lo}; // @[Cat.scala 30:58]
  assign remainder_hi_hi = nextMulReg1[128:64]; // @[Multiplier.scala 122:34]
  assign remainder_lo = nextMulReg1[63:0]; // @[Multiplier.scala 122:67]
  assign _remainder_T = {remainder_hi_hi,remainder_hi_lo,remainder_lo}; // @[Cat.scala 30:58]
  assign _count_T_1 = count + 7'h1; // @[Multiplier.scala 124:20]
  assign _T_28 = count == 7'h7; // @[Multiplier.scala 125:25]
  assign _T_29 = eOut | _T_28; // @[Multiplier.scala 125:16]
  assign _T_30 = state == 3'h3; // @[Multiplier.scala 130:39]
  assign unrolls_less = subtractor[64]; // @[Multiplier.scala 134:28]
  assign unrolls_hi_hi = unrolls_less ? remainder[127:64] : subtractor[63:0]; // @[Multiplier.scala 135:14]
  assign unrolls_lo = ~unrolls_less; // @[Multiplier.scala 135:67]
  assign unrolls_0 = {unrolls_hi_hi,remainder[63:0],unrolls_lo}; // @[Cat.scala 30:58]
  assign _T_31 = count == 7'h40; // @[Multiplier.scala 139:17]
  assign _divby0_T = count == 7'h0; // @[Multiplier.scala 147:24]
  assign divby0 = _divby0_T & unrolls_lo; // @[Multiplier.scala 147:30]
  assign divisorMSB_hi = divisor[63:32]; // @[CircuitMath.scala 35:17]
  assign divisorMSB_lo = divisor[31:0]; // @[CircuitMath.scala 36:17]
  assign divisorMSB_hi_1 = |divisorMSB_hi; // @[CircuitMath.scala 37:22]
  assign divisorMSB_hi_2 = divisorMSB_hi[31:16]; // @[CircuitMath.scala 35:17]
  assign divisorMSB_lo_1 = divisorMSB_hi[15:0]; // @[CircuitMath.scala 36:17]
  assign divisorMSB_hi_3 = |divisorMSB_hi_2; // @[CircuitMath.scala 37:22]
  assign divisorMSB_hi_4 = divisorMSB_hi_2[15:8]; // @[CircuitMath.scala 35:17]
  assign divisorMSB_lo_2 = divisorMSB_hi_2[7:0]; // @[CircuitMath.scala 36:17]
  assign divisorMSB_hi_5 = |divisorMSB_hi_4; // @[CircuitMath.scala 37:22]
  assign divisorMSB_hi_6 = divisorMSB_hi_4[7:4]; // @[CircuitMath.scala 35:17]
  assign divisorMSB_lo_3 = divisorMSB_hi_4[3:0]; // @[CircuitMath.scala 36:17]
  assign divisorMSB_hi_7 = |divisorMSB_hi_6; // @[CircuitMath.scala 37:22]
  assign _divisorMSB_T_4 = divisorMSB_hi_6[2] ? 2'h2 : {{1'd0}, divisorMSB_hi_6[1]}; // @[CircuitMath.scala 32:10]
  assign _divisorMSB_T_5 = divisorMSB_hi_6[3] ? 2'h3 : _divisorMSB_T_4; // @[CircuitMath.scala 32:10]
  assign _divisorMSB_T_9 = divisorMSB_lo_3[2] ? 2'h2 : {{1'd0}, divisorMSB_lo_3[1]}; // @[CircuitMath.scala 32:10]
  assign _divisorMSB_T_10 = divisorMSB_lo_3[3] ? 2'h3 : _divisorMSB_T_9; // @[CircuitMath.scala 32:10]
  assign divisorMSB_lo_4 = divisorMSB_hi_7 ? _divisorMSB_T_5 : _divisorMSB_T_10; // @[CircuitMath.scala 38:21]
  assign _divisorMSB_T_11 = {divisorMSB_hi_7,divisorMSB_lo_4}; // @[Cat.scala 30:58]
  assign divisorMSB_hi_8 = divisorMSB_lo_2[7:4]; // @[CircuitMath.scala 35:17]
  assign divisorMSB_lo_5 = divisorMSB_lo_2[3:0]; // @[CircuitMath.scala 36:17]
  assign divisorMSB_hi_9 = |divisorMSB_hi_8; // @[CircuitMath.scala 37:22]
  assign _divisorMSB_T_15 = divisorMSB_hi_8[2] ? 2'h2 : {{1'd0}, divisorMSB_hi_8[1]}; // @[CircuitMath.scala 32:10]
  assign _divisorMSB_T_16 = divisorMSB_hi_8[3] ? 2'h3 : _divisorMSB_T_15; // @[CircuitMath.scala 32:10]
  assign _divisorMSB_T_20 = divisorMSB_lo_5[2] ? 2'h2 : {{1'd0}, divisorMSB_lo_5[1]}; // @[CircuitMath.scala 32:10]
  assign _divisorMSB_T_21 = divisorMSB_lo_5[3] ? 2'h3 : _divisorMSB_T_20; // @[CircuitMath.scala 32:10]
  assign divisorMSB_lo_6 = divisorMSB_hi_9 ? _divisorMSB_T_16 : _divisorMSB_T_21; // @[CircuitMath.scala 38:21]
  assign _divisorMSB_T_22 = {divisorMSB_hi_9,divisorMSB_lo_6}; // @[Cat.scala 30:58]
  assign divisorMSB_lo_7 = divisorMSB_hi_5 ? _divisorMSB_T_11 : _divisorMSB_T_22; // @[CircuitMath.scala 38:21]
  assign _divisorMSB_T_23 = {divisorMSB_hi_5,divisorMSB_lo_7}; // @[Cat.scala 30:58]
  assign divisorMSB_hi_10 = divisorMSB_lo_1[15:8]; // @[CircuitMath.scala 35:17]
  assign divisorMSB_lo_8 = divisorMSB_lo_1[7:0]; // @[CircuitMath.scala 36:17]
  assign divisorMSB_hi_11 = |divisorMSB_hi_10; // @[CircuitMath.scala 37:22]
  assign divisorMSB_hi_12 = divisorMSB_hi_10[7:4]; // @[CircuitMath.scala 35:17]
  assign divisorMSB_lo_9 = divisorMSB_hi_10[3:0]; // @[CircuitMath.scala 36:17]
  assign divisorMSB_hi_13 = |divisorMSB_hi_12; // @[CircuitMath.scala 37:22]
  assign _divisorMSB_T_27 = divisorMSB_hi_12[2] ? 2'h2 : {{1'd0}, divisorMSB_hi_12[1]}; // @[CircuitMath.scala 32:10]
  assign _divisorMSB_T_28 = divisorMSB_hi_12[3] ? 2'h3 : _divisorMSB_T_27; // @[CircuitMath.scala 32:10]
  assign _divisorMSB_T_32 = divisorMSB_lo_9[2] ? 2'h2 : {{1'd0}, divisorMSB_lo_9[1]}; // @[CircuitMath.scala 32:10]
  assign _divisorMSB_T_33 = divisorMSB_lo_9[3] ? 2'h3 : _divisorMSB_T_32; // @[CircuitMath.scala 32:10]
  assign divisorMSB_lo_10 = divisorMSB_hi_13 ? _divisorMSB_T_28 : _divisorMSB_T_33; // @[CircuitMath.scala 38:21]
  assign _divisorMSB_T_34 = {divisorMSB_hi_13,divisorMSB_lo_10}; // @[Cat.scala 30:58]
  assign divisorMSB_hi_14 = divisorMSB_lo_8[7:4]; // @[CircuitMath.scala 35:17]
  assign divisorMSB_lo_11 = divisorMSB_lo_8[3:0]; // @[CircuitMath.scala 36:17]
  assign divisorMSB_hi_15 = |divisorMSB_hi_14; // @[CircuitMath.scala 37:22]
  assign _divisorMSB_T_38 = divisorMSB_hi_14[2] ? 2'h2 : {{1'd0}, divisorMSB_hi_14[1]}; // @[CircuitMath.scala 32:10]
  assign _divisorMSB_T_39 = divisorMSB_hi_14[3] ? 2'h3 : _divisorMSB_T_38; // @[CircuitMath.scala 32:10]
  assign _divisorMSB_T_43 = divisorMSB_lo_11[2] ? 2'h2 : {{1'd0}, divisorMSB_lo_11[1]}; // @[CircuitMath.scala 32:10]
  assign _divisorMSB_T_44 = divisorMSB_lo_11[3] ? 2'h3 : _divisorMSB_T_43; // @[CircuitMath.scala 32:10]
  assign divisorMSB_lo_12 = divisorMSB_hi_15 ? _divisorMSB_T_39 : _divisorMSB_T_44; // @[CircuitMath.scala 38:21]
  assign _divisorMSB_T_45 = {divisorMSB_hi_15,divisorMSB_lo_12}; // @[Cat.scala 30:58]
  assign divisorMSB_lo_13 = divisorMSB_hi_11 ? _divisorMSB_T_34 : _divisorMSB_T_45; // @[CircuitMath.scala 38:21]
  assign _divisorMSB_T_46 = {divisorMSB_hi_11,divisorMSB_lo_13}; // @[Cat.scala 30:58]
  assign divisorMSB_lo_14 = divisorMSB_hi_3 ? _divisorMSB_T_23 : _divisorMSB_T_46; // @[CircuitMath.scala 38:21]
  assign _divisorMSB_T_47 = {divisorMSB_hi_3,divisorMSB_lo_14}; // @[Cat.scala 30:58]
  assign divisorMSB_hi_16 = divisorMSB_lo[31:16]; // @[CircuitMath.scala 35:17]
  assign divisorMSB_lo_15 = divisorMSB_lo[15:0]; // @[CircuitMath.scala 36:17]
  assign divisorMSB_hi_17 = |divisorMSB_hi_16; // @[CircuitMath.scala 37:22]
  assign divisorMSB_hi_18 = divisorMSB_hi_16[15:8]; // @[CircuitMath.scala 35:17]
  assign divisorMSB_lo_16 = divisorMSB_hi_16[7:0]; // @[CircuitMath.scala 36:17]
  assign divisorMSB_hi_19 = |divisorMSB_hi_18; // @[CircuitMath.scala 37:22]
  assign divisorMSB_hi_20 = divisorMSB_hi_18[7:4]; // @[CircuitMath.scala 35:17]
  assign divisorMSB_lo_17 = divisorMSB_hi_18[3:0]; // @[CircuitMath.scala 36:17]
  assign divisorMSB_hi_21 = |divisorMSB_hi_20; // @[CircuitMath.scala 37:22]
  assign _divisorMSB_T_51 = divisorMSB_hi_20[2] ? 2'h2 : {{1'd0}, divisorMSB_hi_20[1]}; // @[CircuitMath.scala 32:10]
  assign _divisorMSB_T_52 = divisorMSB_hi_20[3] ? 2'h3 : _divisorMSB_T_51; // @[CircuitMath.scala 32:10]
  assign _divisorMSB_T_56 = divisorMSB_lo_17[2] ? 2'h2 : {{1'd0}, divisorMSB_lo_17[1]}; // @[CircuitMath.scala 32:10]
  assign _divisorMSB_T_57 = divisorMSB_lo_17[3] ? 2'h3 : _divisorMSB_T_56; // @[CircuitMath.scala 32:10]
  assign divisorMSB_lo_18 = divisorMSB_hi_21 ? _divisorMSB_T_52 : _divisorMSB_T_57; // @[CircuitMath.scala 38:21]
  assign _divisorMSB_T_58 = {divisorMSB_hi_21,divisorMSB_lo_18}; // @[Cat.scala 30:58]
  assign divisorMSB_hi_22 = divisorMSB_lo_16[7:4]; // @[CircuitMath.scala 35:17]
  assign divisorMSB_lo_19 = divisorMSB_lo_16[3:0]; // @[CircuitMath.scala 36:17]
  assign divisorMSB_hi_23 = |divisorMSB_hi_22; // @[CircuitMath.scala 37:22]
  assign _divisorMSB_T_62 = divisorMSB_hi_22[2] ? 2'h2 : {{1'd0}, divisorMSB_hi_22[1]}; // @[CircuitMath.scala 32:10]
  assign _divisorMSB_T_63 = divisorMSB_hi_22[3] ? 2'h3 : _divisorMSB_T_62; // @[CircuitMath.scala 32:10]
  assign _divisorMSB_T_67 = divisorMSB_lo_19[2] ? 2'h2 : {{1'd0}, divisorMSB_lo_19[1]}; // @[CircuitMath.scala 32:10]
  assign _divisorMSB_T_68 = divisorMSB_lo_19[3] ? 2'h3 : _divisorMSB_T_67; // @[CircuitMath.scala 32:10]
  assign divisorMSB_lo_20 = divisorMSB_hi_23 ? _divisorMSB_T_63 : _divisorMSB_T_68; // @[CircuitMath.scala 38:21]
  assign _divisorMSB_T_69 = {divisorMSB_hi_23,divisorMSB_lo_20}; // @[Cat.scala 30:58]
  assign divisorMSB_lo_21 = divisorMSB_hi_19 ? _divisorMSB_T_58 : _divisorMSB_T_69; // @[CircuitMath.scala 38:21]
  assign _divisorMSB_T_70 = {divisorMSB_hi_19,divisorMSB_lo_21}; // @[Cat.scala 30:58]
  assign divisorMSB_hi_24 = divisorMSB_lo_15[15:8]; // @[CircuitMath.scala 35:17]
  assign divisorMSB_lo_22 = divisorMSB_lo_15[7:0]; // @[CircuitMath.scala 36:17]
  assign divisorMSB_hi_25 = |divisorMSB_hi_24; // @[CircuitMath.scala 37:22]
  assign divisorMSB_hi_26 = divisorMSB_hi_24[7:4]; // @[CircuitMath.scala 35:17]
  assign divisorMSB_lo_23 = divisorMSB_hi_24[3:0]; // @[CircuitMath.scala 36:17]
  assign divisorMSB_hi_27 = |divisorMSB_hi_26; // @[CircuitMath.scala 37:22]
  assign _divisorMSB_T_74 = divisorMSB_hi_26[2] ? 2'h2 : {{1'd0}, divisorMSB_hi_26[1]}; // @[CircuitMath.scala 32:10]
  assign _divisorMSB_T_75 = divisorMSB_hi_26[3] ? 2'h3 : _divisorMSB_T_74; // @[CircuitMath.scala 32:10]
  assign _divisorMSB_T_79 = divisorMSB_lo_23[2] ? 2'h2 : {{1'd0}, divisorMSB_lo_23[1]}; // @[CircuitMath.scala 32:10]
  assign _divisorMSB_T_80 = divisorMSB_lo_23[3] ? 2'h3 : _divisorMSB_T_79; // @[CircuitMath.scala 32:10]
  assign divisorMSB_lo_24 = divisorMSB_hi_27 ? _divisorMSB_T_75 : _divisorMSB_T_80; // @[CircuitMath.scala 38:21]
  assign _divisorMSB_T_81 = {divisorMSB_hi_27,divisorMSB_lo_24}; // @[Cat.scala 30:58]
  assign divisorMSB_hi_28 = divisorMSB_lo_22[7:4]; // @[CircuitMath.scala 35:17]
  assign divisorMSB_lo_25 = divisorMSB_lo_22[3:0]; // @[CircuitMath.scala 36:17]
  assign divisorMSB_hi_29 = |divisorMSB_hi_28; // @[CircuitMath.scala 37:22]
  assign _divisorMSB_T_85 = divisorMSB_hi_28[2] ? 2'h2 : {{1'd0}, divisorMSB_hi_28[1]}; // @[CircuitMath.scala 32:10]
  assign _divisorMSB_T_86 = divisorMSB_hi_28[3] ? 2'h3 : _divisorMSB_T_85; // @[CircuitMath.scala 32:10]
  assign _divisorMSB_T_90 = divisorMSB_lo_25[2] ? 2'h2 : {{1'd0}, divisorMSB_lo_25[1]}; // @[CircuitMath.scala 32:10]
  assign _divisorMSB_T_91 = divisorMSB_lo_25[3] ? 2'h3 : _divisorMSB_T_90; // @[CircuitMath.scala 32:10]
  assign divisorMSB_lo_26 = divisorMSB_hi_29 ? _divisorMSB_T_86 : _divisorMSB_T_91; // @[CircuitMath.scala 38:21]
  assign _divisorMSB_T_92 = {divisorMSB_hi_29,divisorMSB_lo_26}; // @[Cat.scala 30:58]
  assign divisorMSB_lo_27 = divisorMSB_hi_25 ? _divisorMSB_T_81 : _divisorMSB_T_92; // @[CircuitMath.scala 38:21]
  assign _divisorMSB_T_93 = {divisorMSB_hi_25,divisorMSB_lo_27}; // @[Cat.scala 30:58]
  assign divisorMSB_lo_28 = divisorMSB_hi_17 ? _divisorMSB_T_70 : _divisorMSB_T_93; // @[CircuitMath.scala 38:21]
  assign _divisorMSB_T_94 = {divisorMSB_hi_17,divisorMSB_lo_28}; // @[Cat.scala 30:58]
  assign divisorMSB_lo_29 = divisorMSB_hi_1 ? _divisorMSB_T_47 : _divisorMSB_T_94; // @[CircuitMath.scala 38:21]
  assign divisorMSB = {divisorMSB_hi_1,divisorMSB_lo_29}; // @[Cat.scala 30:58]
  assign dividendMSB_hi = remainder[63:32]; // @[CircuitMath.scala 35:17]
  assign dividendMSB_lo = remainder[31:0]; // @[CircuitMath.scala 36:17]
  assign dividendMSB_hi_1 = |dividendMSB_hi; // @[CircuitMath.scala 37:22]
  assign dividendMSB_hi_2 = dividendMSB_hi[31:16]; // @[CircuitMath.scala 35:17]
  assign dividendMSB_lo_1 = dividendMSB_hi[15:0]; // @[CircuitMath.scala 36:17]
  assign dividendMSB_hi_3 = |dividendMSB_hi_2; // @[CircuitMath.scala 37:22]
  assign dividendMSB_hi_4 = dividendMSB_hi_2[15:8]; // @[CircuitMath.scala 35:17]
  assign dividendMSB_lo_2 = dividendMSB_hi_2[7:0]; // @[CircuitMath.scala 36:17]
  assign dividendMSB_hi_5 = |dividendMSB_hi_4; // @[CircuitMath.scala 37:22]
  assign dividendMSB_hi_6 = dividendMSB_hi_4[7:4]; // @[CircuitMath.scala 35:17]
  assign dividendMSB_lo_3 = dividendMSB_hi_4[3:0]; // @[CircuitMath.scala 36:17]
  assign dividendMSB_hi_7 = |dividendMSB_hi_6; // @[CircuitMath.scala 37:22]
  assign _dividendMSB_T_4 = dividendMSB_hi_6[2] ? 2'h2 : {{1'd0}, dividendMSB_hi_6[1]}; // @[CircuitMath.scala 32:10]
  assign _dividendMSB_T_5 = dividendMSB_hi_6[3] ? 2'h3 : _dividendMSB_T_4; // @[CircuitMath.scala 32:10]
  assign _dividendMSB_T_9 = dividendMSB_lo_3[2] ? 2'h2 : {{1'd0}, dividendMSB_lo_3[1]}; // @[CircuitMath.scala 32:10]
  assign _dividendMSB_T_10 = dividendMSB_lo_3[3] ? 2'h3 : _dividendMSB_T_9; // @[CircuitMath.scala 32:10]
  assign dividendMSB_lo_4 = dividendMSB_hi_7 ? _dividendMSB_T_5 : _dividendMSB_T_10; // @[CircuitMath.scala 38:21]
  assign _dividendMSB_T_11 = {dividendMSB_hi_7,dividendMSB_lo_4}; // @[Cat.scala 30:58]
  assign dividendMSB_hi_8 = dividendMSB_lo_2[7:4]; // @[CircuitMath.scala 35:17]
  assign dividendMSB_lo_5 = dividendMSB_lo_2[3:0]; // @[CircuitMath.scala 36:17]
  assign dividendMSB_hi_9 = |dividendMSB_hi_8; // @[CircuitMath.scala 37:22]
  assign _dividendMSB_T_15 = dividendMSB_hi_8[2] ? 2'h2 : {{1'd0}, dividendMSB_hi_8[1]}; // @[CircuitMath.scala 32:10]
  assign _dividendMSB_T_16 = dividendMSB_hi_8[3] ? 2'h3 : _dividendMSB_T_15; // @[CircuitMath.scala 32:10]
  assign _dividendMSB_T_20 = dividendMSB_lo_5[2] ? 2'h2 : {{1'd0}, dividendMSB_lo_5[1]}; // @[CircuitMath.scala 32:10]
  assign _dividendMSB_T_21 = dividendMSB_lo_5[3] ? 2'h3 : _dividendMSB_T_20; // @[CircuitMath.scala 32:10]
  assign dividendMSB_lo_6 = dividendMSB_hi_9 ? _dividendMSB_T_16 : _dividendMSB_T_21; // @[CircuitMath.scala 38:21]
  assign _dividendMSB_T_22 = {dividendMSB_hi_9,dividendMSB_lo_6}; // @[Cat.scala 30:58]
  assign dividendMSB_lo_7 = dividendMSB_hi_5 ? _dividendMSB_T_11 : _dividendMSB_T_22; // @[CircuitMath.scala 38:21]
  assign _dividendMSB_T_23 = {dividendMSB_hi_5,dividendMSB_lo_7}; // @[Cat.scala 30:58]
  assign dividendMSB_hi_10 = dividendMSB_lo_1[15:8]; // @[CircuitMath.scala 35:17]
  assign dividendMSB_lo_8 = dividendMSB_lo_1[7:0]; // @[CircuitMath.scala 36:17]
  assign dividendMSB_hi_11 = |dividendMSB_hi_10; // @[CircuitMath.scala 37:22]
  assign dividendMSB_hi_12 = dividendMSB_hi_10[7:4]; // @[CircuitMath.scala 35:17]
  assign dividendMSB_lo_9 = dividendMSB_hi_10[3:0]; // @[CircuitMath.scala 36:17]
  assign dividendMSB_hi_13 = |dividendMSB_hi_12; // @[CircuitMath.scala 37:22]
  assign _dividendMSB_T_27 = dividendMSB_hi_12[2] ? 2'h2 : {{1'd0}, dividendMSB_hi_12[1]}; // @[CircuitMath.scala 32:10]
  assign _dividendMSB_T_28 = dividendMSB_hi_12[3] ? 2'h3 : _dividendMSB_T_27; // @[CircuitMath.scala 32:10]
  assign _dividendMSB_T_32 = dividendMSB_lo_9[2] ? 2'h2 : {{1'd0}, dividendMSB_lo_9[1]}; // @[CircuitMath.scala 32:10]
  assign _dividendMSB_T_33 = dividendMSB_lo_9[3] ? 2'h3 : _dividendMSB_T_32; // @[CircuitMath.scala 32:10]
  assign dividendMSB_lo_10 = dividendMSB_hi_13 ? _dividendMSB_T_28 : _dividendMSB_T_33; // @[CircuitMath.scala 38:21]
  assign _dividendMSB_T_34 = {dividendMSB_hi_13,dividendMSB_lo_10}; // @[Cat.scala 30:58]
  assign dividendMSB_hi_14 = dividendMSB_lo_8[7:4]; // @[CircuitMath.scala 35:17]
  assign dividendMSB_lo_11 = dividendMSB_lo_8[3:0]; // @[CircuitMath.scala 36:17]
  assign dividendMSB_hi_15 = |dividendMSB_hi_14; // @[CircuitMath.scala 37:22]
  assign _dividendMSB_T_38 = dividendMSB_hi_14[2] ? 2'h2 : {{1'd0}, dividendMSB_hi_14[1]}; // @[CircuitMath.scala 32:10]
  assign _dividendMSB_T_39 = dividendMSB_hi_14[3] ? 2'h3 : _dividendMSB_T_38; // @[CircuitMath.scala 32:10]
  assign _dividendMSB_T_43 = dividendMSB_lo_11[2] ? 2'h2 : {{1'd0}, dividendMSB_lo_11[1]}; // @[CircuitMath.scala 32:10]
  assign _dividendMSB_T_44 = dividendMSB_lo_11[3] ? 2'h3 : _dividendMSB_T_43; // @[CircuitMath.scala 32:10]
  assign dividendMSB_lo_12 = dividendMSB_hi_15 ? _dividendMSB_T_39 : _dividendMSB_T_44; // @[CircuitMath.scala 38:21]
  assign _dividendMSB_T_45 = {dividendMSB_hi_15,dividendMSB_lo_12}; // @[Cat.scala 30:58]
  assign dividendMSB_lo_13 = dividendMSB_hi_11 ? _dividendMSB_T_34 : _dividendMSB_T_45; // @[CircuitMath.scala 38:21]
  assign _dividendMSB_T_46 = {dividendMSB_hi_11,dividendMSB_lo_13}; // @[Cat.scala 30:58]
  assign dividendMSB_lo_14 = dividendMSB_hi_3 ? _dividendMSB_T_23 : _dividendMSB_T_46; // @[CircuitMath.scala 38:21]
  assign _dividendMSB_T_47 = {dividendMSB_hi_3,dividendMSB_lo_14}; // @[Cat.scala 30:58]
  assign dividendMSB_hi_16 = dividendMSB_lo[31:16]; // @[CircuitMath.scala 35:17]
  assign dividendMSB_lo_15 = dividendMSB_lo[15:0]; // @[CircuitMath.scala 36:17]
  assign dividendMSB_hi_17 = |dividendMSB_hi_16; // @[CircuitMath.scala 37:22]
  assign dividendMSB_hi_18 = dividendMSB_hi_16[15:8]; // @[CircuitMath.scala 35:17]
  assign dividendMSB_lo_16 = dividendMSB_hi_16[7:0]; // @[CircuitMath.scala 36:17]
  assign dividendMSB_hi_19 = |dividendMSB_hi_18; // @[CircuitMath.scala 37:22]
  assign dividendMSB_hi_20 = dividendMSB_hi_18[7:4]; // @[CircuitMath.scala 35:17]
  assign dividendMSB_lo_17 = dividendMSB_hi_18[3:0]; // @[CircuitMath.scala 36:17]
  assign dividendMSB_hi_21 = |dividendMSB_hi_20; // @[CircuitMath.scala 37:22]
  assign _dividendMSB_T_51 = dividendMSB_hi_20[2] ? 2'h2 : {{1'd0}, dividendMSB_hi_20[1]}; // @[CircuitMath.scala 32:10]
  assign _dividendMSB_T_52 = dividendMSB_hi_20[3] ? 2'h3 : _dividendMSB_T_51; // @[CircuitMath.scala 32:10]
  assign _dividendMSB_T_56 = dividendMSB_lo_17[2] ? 2'h2 : {{1'd0}, dividendMSB_lo_17[1]}; // @[CircuitMath.scala 32:10]
  assign _dividendMSB_T_57 = dividendMSB_lo_17[3] ? 2'h3 : _dividendMSB_T_56; // @[CircuitMath.scala 32:10]
  assign dividendMSB_lo_18 = dividendMSB_hi_21 ? _dividendMSB_T_52 : _dividendMSB_T_57; // @[CircuitMath.scala 38:21]
  assign _dividendMSB_T_58 = {dividendMSB_hi_21,dividendMSB_lo_18}; // @[Cat.scala 30:58]
  assign dividendMSB_hi_22 = dividendMSB_lo_16[7:4]; // @[CircuitMath.scala 35:17]
  assign dividendMSB_lo_19 = dividendMSB_lo_16[3:0]; // @[CircuitMath.scala 36:17]
  assign dividendMSB_hi_23 = |dividendMSB_hi_22; // @[CircuitMath.scala 37:22]
  assign _dividendMSB_T_62 = dividendMSB_hi_22[2] ? 2'h2 : {{1'd0}, dividendMSB_hi_22[1]}; // @[CircuitMath.scala 32:10]
  assign _dividendMSB_T_63 = dividendMSB_hi_22[3] ? 2'h3 : _dividendMSB_T_62; // @[CircuitMath.scala 32:10]
  assign _dividendMSB_T_67 = dividendMSB_lo_19[2] ? 2'h2 : {{1'd0}, dividendMSB_lo_19[1]}; // @[CircuitMath.scala 32:10]
  assign _dividendMSB_T_68 = dividendMSB_lo_19[3] ? 2'h3 : _dividendMSB_T_67; // @[CircuitMath.scala 32:10]
  assign dividendMSB_lo_20 = dividendMSB_hi_23 ? _dividendMSB_T_63 : _dividendMSB_T_68; // @[CircuitMath.scala 38:21]
  assign _dividendMSB_T_69 = {dividendMSB_hi_23,dividendMSB_lo_20}; // @[Cat.scala 30:58]
  assign dividendMSB_lo_21 = dividendMSB_hi_19 ? _dividendMSB_T_58 : _dividendMSB_T_69; // @[CircuitMath.scala 38:21]
  assign _dividendMSB_T_70 = {dividendMSB_hi_19,dividendMSB_lo_21}; // @[Cat.scala 30:58]
  assign dividendMSB_hi_24 = dividendMSB_lo_15[15:8]; // @[CircuitMath.scala 35:17]
  assign dividendMSB_lo_22 = dividendMSB_lo_15[7:0]; // @[CircuitMath.scala 36:17]
  assign dividendMSB_hi_25 = |dividendMSB_hi_24; // @[CircuitMath.scala 37:22]
  assign dividendMSB_hi_26 = dividendMSB_hi_24[7:4]; // @[CircuitMath.scala 35:17]
  assign dividendMSB_lo_23 = dividendMSB_hi_24[3:0]; // @[CircuitMath.scala 36:17]
  assign dividendMSB_hi_27 = |dividendMSB_hi_26; // @[CircuitMath.scala 37:22]
  assign _dividendMSB_T_74 = dividendMSB_hi_26[2] ? 2'h2 : {{1'd0}, dividendMSB_hi_26[1]}; // @[CircuitMath.scala 32:10]
  assign _dividendMSB_T_75 = dividendMSB_hi_26[3] ? 2'h3 : _dividendMSB_T_74; // @[CircuitMath.scala 32:10]
  assign _dividendMSB_T_79 = dividendMSB_lo_23[2] ? 2'h2 : {{1'd0}, dividendMSB_lo_23[1]}; // @[CircuitMath.scala 32:10]
  assign _dividendMSB_T_80 = dividendMSB_lo_23[3] ? 2'h3 : _dividendMSB_T_79; // @[CircuitMath.scala 32:10]
  assign dividendMSB_lo_24 = dividendMSB_hi_27 ? _dividendMSB_T_75 : _dividendMSB_T_80; // @[CircuitMath.scala 38:21]
  assign _dividendMSB_T_81 = {dividendMSB_hi_27,dividendMSB_lo_24}; // @[Cat.scala 30:58]
  assign dividendMSB_hi_28 = dividendMSB_lo_22[7:4]; // @[CircuitMath.scala 35:17]
  assign dividendMSB_lo_25 = dividendMSB_lo_22[3:0]; // @[CircuitMath.scala 36:17]
  assign dividendMSB_hi_29 = |dividendMSB_hi_28; // @[CircuitMath.scala 37:22]
  assign _dividendMSB_T_85 = dividendMSB_hi_28[2] ? 2'h2 : {{1'd0}, dividendMSB_hi_28[1]}; // @[CircuitMath.scala 32:10]
  assign _dividendMSB_T_86 = dividendMSB_hi_28[3] ? 2'h3 : _dividendMSB_T_85; // @[CircuitMath.scala 32:10]
  assign _dividendMSB_T_90 = dividendMSB_lo_25[2] ? 2'h2 : {{1'd0}, dividendMSB_lo_25[1]}; // @[CircuitMath.scala 32:10]
  assign _dividendMSB_T_91 = dividendMSB_lo_25[3] ? 2'h3 : _dividendMSB_T_90; // @[CircuitMath.scala 32:10]
  assign dividendMSB_lo_26 = dividendMSB_hi_29 ? _dividendMSB_T_86 : _dividendMSB_T_91; // @[CircuitMath.scala 38:21]
  assign _dividendMSB_T_92 = {dividendMSB_hi_29,dividendMSB_lo_26}; // @[Cat.scala 30:58]
  assign dividendMSB_lo_27 = dividendMSB_hi_25 ? _dividendMSB_T_81 : _dividendMSB_T_92; // @[CircuitMath.scala 38:21]
  assign _dividendMSB_T_93 = {dividendMSB_hi_25,dividendMSB_lo_27}; // @[Cat.scala 30:58]
  assign dividendMSB_lo_28 = dividendMSB_hi_17 ? _dividendMSB_T_70 : _dividendMSB_T_93; // @[CircuitMath.scala 38:21]
  assign _dividendMSB_T_94 = {dividendMSB_hi_17,dividendMSB_lo_28}; // @[Cat.scala 30:58]
  assign dividendMSB_lo_29 = dividendMSB_hi_1 ? _dividendMSB_T_47 : _dividendMSB_T_94; // @[CircuitMath.scala 38:21]
  assign dividendMSB = {dividendMSB_hi_1,dividendMSB_lo_29}; // @[Cat.scala 30:58]
  assign _eOutPos_T_1 = dividendMSB - divisorMSB; // @[Multiplier.scala 153:35]
  assign eOutPos = ~_eOutPos_T_1; // @[Multiplier.scala 153:21]
  assign _eOut_T_11 = _divby0_T & ~divby0; // @[Multiplier.scala 154:30]
  assign _eOut_T_12 = eOutPos >= 6'h1; // @[Multiplier.scala 154:52]
  assign eOut_1 = _eOut_T_11 & _eOut_T_12; // @[Multiplier.scala 154:41]
  assign _GEN_39 = {{63'd0}, remainder[63:0]}; // @[Multiplier.scala 156:39]
  assign _remainder_T_2 = _GEN_39 << eOutPos; // @[Multiplier.scala 156:39]
  assign _GEN_16 = eOut_1 ? {{2'd0}, _remainder_T_2} : unrolls_0; // @[Multiplier.scala 155:19]
  assign _T_33 = divby0 & ~isHi; // @[Multiplier.scala 160:18]
  assign _T_34 = io_resp_ready & io_resp_valid; // @[Decoupled.scala 40:37]
  assign _T_35 = _T_34 | io_kill; // @[Multiplier.scala 162:24]
  assign _T_36 = io_req_ready & io_req_valid; // @[Decoupled.scala 40:37]
  assign _state_T_1 = lhs_sign | rhs_sign; // @[Multiplier.scala 166:46]
  assign _count_T_7 = cmdMul & ~io_req_bits_dw; // @[Multiplier.scala 169:46]
  assign _count_T_8 = _count_T_7 ? 3'h4 : 3'h0; // @[Multiplier.scala 169:38]
  assign _neg_out_T = lhs_sign != rhs_sign; // @[Multiplier.scala 170:46]
  assign _divisor_T = {rhs_sign,hi_1,lo_1}; // @[Cat.scala 30:58]
  assign _outMul_T_1 = state & 3'h1; // @[Multiplier.scala 176:23]
  assign outMul = _outMul_T_1 == 3'h0; // @[Multiplier.scala 176:52]
  assign _loOut_T_3 = ~req_dw & outMul; // @[Multiplier.scala 177:48]
  assign loOut = _loOut_T_3 ? result[63:32] : result[31:0]; // @[Multiplier.scala 177:18]
  assign _hiOut_T_4 = loOut[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  assign hiOut = req_dw ? result[63:32] : _hiOut_T_4; // @[Multiplier.scala 178:18]
  assign _io_resp_valid_T = state == 3'h6; // @[Multiplier.scala 182:27]
  assign _io_resp_valid_T_1 = state == 3'h7; // @[Multiplier.scala 182:51]
  assign io_req_ready = state == 3'h0; // @[Multiplier.scala 183:16]
  assign io_resp_valid = _io_resp_valid_T | _io_resp_valid_T_1; // @[Multiplier.scala 182:17]
  assign io_resp_bits_data = {hiOut,loOut}; // @[Multiplier.scala 181:21]
  assign io_resp_bits_tag = req_tag; // @[Multiplier.scala 179:20]
  assign MulDiv_cov_read_addr = MulDiv_state;
  assign MulDiv_cov_read_data = MulDiv_cov[MulDiv_cov_read_addr]; // @[Coverage map for MulDiv]
  assign MulDiv_cov_write_data = 1'h1;
  assign MulDiv_cov_write_addr = MulDiv_state;
  assign MulDiv_cov_write_mask = 1'h1;
  assign MulDiv_cov_write_en = 1'h1;
  assign mux_cond_0 = dividendMSB_hi_13;
  assign mux_cond_1 = dividendMSB_lo_19[3];
  assign mux_cond_2 = divisorMSB_hi_21;
  assign mux_cond_3 = dividendMSB_hi_28[3];
  assign mux_cond_4 = divisorMSB_hi_3;
  assign mux_cond_5 = divisorMSB_lo_5[2];
  assign mux_cond_6 = dividendMSB_lo_19[2];
  assign mux_cond_7 = divisorMSB_hi_14[2];
  assign mux_cond_8 = divisorMSB_hi_26[3];
  assign mux_cond_9 = dividendMSB_hi_7;
  assign mux_cond_10 = divisorMSB_hi_28[3];
  assign mux_cond_11 = dividendMSB_hi_20[2];
  assign mux_cond_12 = dividendMSB_hi_8[3];
  assign mux_cond_13 = dividendMSB_hi_27;
  assign mux_cond_14 = divisorMSB_lo_19[2];
  assign mux_cond_15 = divisorMSB_lo_9[3];
  assign mux_cond_16 = dividendMSB_lo_3[3];
  assign mux_cond_17 = dividendMSB_hi_22[2];
  assign mux_cond_18 = divisorMSB_hi_6[3];
  assign mux_cond_19 = dividendMSB_lo_23[2];
  assign mux_cond_20 = divisorMSB_hi_26[2];
  assign mux_cond_21 = dividendMSB_hi_6[3];
  assign mux_cond_22 = divisorMSB_lo_19[3];
  assign mux_cond_23 = divisorMSB_lo_17[2];
  assign mux_cond_24 = dividendMSB_lo_3[2];
  assign mux_cond_25 = divisorMSB_hi_29;
  assign mux_cond_26 = dividendMSB_lo_17[2];
  assign mux_cond_27 = dividendMSB_lo_25[3];
  assign mux_cond_28 = divisorMSB_hi_7;
  assign mux_cond_29 = dividendMSB_hi_29;
  assign mux_cond_30 = divisorMSB_lo_9[2];
  assign mux_cond_31 = dividendMSB_hi_9;
  assign mux_cond_32 = divisorMSB_hi_28[2];
  assign mux_cond_33 = divisorMSB_hi_25;
  assign mux_cond_34 = divisorMSB_lo_25[2];
  assign mux_cond_35 = divisorMSB_hi_11;
  assign mux_cond_36 = divisorMSB_lo_23[2];
  assign mux_cond_37 = dividendMSB_hi_1;
  assign mux_cond_38 = dividendMSB_lo_9[2];
  assign mux_cond_39 = divisorMSB_hi_17;
  assign mux_cond_40 = dividendMSB_lo_17[3];
  assign mux_cond_41 = divisorMSB_lo_11[2];
  assign mux_cond_42 = divisorMSB_hi_15;
  assign mux_cond_43 = divisorMSB_hi_14[3];
  assign mux_cond_44 = divisor[63];
  assign mux_cond_45 = divisorMSB_hi_6[2];
  assign mux_cond_46 = divisorMSB_hi_8[3];
  assign mux_cond_47 = divisorMSB_hi_20[3];
  assign mux_cond_48 = dividendMSB_hi_28[2];
  assign mux_cond_49 = unrolls_less;
  assign mux_cond_50 = divisorMSB_hi_8[2];
  assign mux_cond_51 = divisorMSB_hi_23;
  assign mux_cond_52 = dividendMSB_lo_23[3];
  assign mux_cond_53 = divisorMSB_hi_22[3];
  assign mux_cond_54 = divisorMSB_lo_3[2];
  assign mux_cond_55 = divisorMSB_lo_25[3];
  assign mux_cond_56 = divisorMSB_lo_23[3];
  assign mux_cond_57 = divisorMSB_hi_27;
  assign mux_cond_58 = divisorMSB_hi_12[2];
  assign mux_cond_59 = dividendMSB_lo_11[3];
  assign mux_cond_60 = divisorMSB_lo_3[3];
  assign mux_cond_61 = dividendMSB_hi_21;
  assign mux_cond_62 = dividendMSB_hi_12[3];
  assign mux_cond_63 = dividendMSB_hi_14[3];
  assign mux_cond_64 = divisorMSB_hi_20[2];
  assign mux_cond_65 = dividendMSB_lo_5[2];
  assign mux_cond_66 = dividendMSB_hi_17;
  assign mux_cond_67 = dividendMSB_hi_8[2];
  assign mux_cond_68 = remainder[63];
  assign mux_cond_69 = dividendMSB_hi_12[2];
  assign mux_cond_70 = divisorMSB_hi_22[2];
  assign mux_cond_71 = dividendMSB_hi_19;
  assign mux_cond_72 = dividendMSB_hi_5;
  assign mux_cond_73 = loOut[31];
  assign mux_cond_74 = dividendMSB_hi_14[2];
  assign mux_cond_75 = divisorMSB_hi_12[3];
  assign mux_cond_76 = divisorMSB_hi_5;
  assign mux_cond_77 = divisorMSB_lo_11[3];
  assign mux_cond_78 = divisorMSB_lo_5[3];
  assign mux_cond_79 = dividendMSB_lo_5[3];
  assign mux_cond_80 = dividendMSB_hi_26[3];
  assign mux_cond_81 = dividendMSB_hi_15;
  assign mux_cond_82 = dividendMSB_hi_25;
  assign mux_cond_83 = divisorMSB_hi_13;
  assign mux_cond_84 = dividendMSB_hi_3;
  assign mux_cond_85 = dividendMSB_hi_23;
  assign mux_cond_86 = dividendMSB_lo_9[3];
  assign mux_cond_87 = divisorMSB_lo_17[3];
  assign mux_cond_88 = dividendMSB_hi_22[3];
  assign mux_cond_89 = dividendMSB_hi_6[2];
  assign mux_cond_90 = dividendMSB_hi_11;
  assign mux_cond_91 = divisorMSB_hi_19;
  assign mux_cond_92 = dividendMSB_lo_11[2];
  assign mux_cond_93 = divisorMSB_hi_9;
  assign mux_cond_94 = dividendMSB_lo_25[2];
  assign mux_cond_95 = divisorMSB_hi_1;
  assign mux_cond_96 = dividendMSB_hi_20[3];
  assign mux_cond_97 = dividendMSB_hi_26[2];
  assign isHi_shl = {isHi, 4'h0};
  assign isHi_pad = {15'h0,isHi_shl};
  assign neg_out_shl = {neg_out, 12'h0};
  assign neg_out_pad = {7'h0,neg_out_shl};
  assign req_dw_shl = {req_dw, 4'h0};
  assign req_dw_pad = {15'h0,req_dw_shl};
  assign state_shl = {state, 8'h0};
  assign state_pad = {9'h0,state_shl};
  assign resHi_shl = {resHi, 1'h0};
  assign resHi_pad = {18'h0,resHi_shl};
  assign mux_cond_0_shl = {mux_cond_0, 12'h0};
  assign mux_cond_0_pad = {7'h0,mux_cond_0_shl};
  assign mux_cond_1_shl = {mux_cond_1, 1'h0};
  assign mux_cond_1_pad = {18'h0,mux_cond_1_shl};
  assign mux_cond_2_shl = mux_cond_2;
  assign mux_cond_2_pad = {19'h0,mux_cond_2_shl};
  assign mux_cond_3_shl = {mux_cond_3, 12'h0};
  assign mux_cond_3_pad = {7'h0,mux_cond_3_shl};
  assign mux_cond_4_shl = {mux_cond_4, 15'h0};
  assign mux_cond_4_pad = {4'h0,mux_cond_4_shl};
  assign mux_cond_5_shl = {mux_cond_5, 11'h0};
  assign mux_cond_5_pad = {8'h0,mux_cond_5_shl};
  assign mux_cond_6_shl = {mux_cond_6, 7'h0};
  assign mux_cond_6_pad = {12'h0,mux_cond_6_shl};
  assign mux_cond_7_shl = {mux_cond_7, 17'h0};
  assign mux_cond_7_pad = {2'h0,mux_cond_7_shl};
  assign mux_cond_8_shl = {mux_cond_8, 11'h0};
  assign mux_cond_8_pad = {8'h0,mux_cond_8_shl};
  assign mux_cond_9_shl = {mux_cond_9, 15'h0};
  assign mux_cond_9_pad = {4'h0,mux_cond_9_shl};
  assign mux_cond_10_shl = {mux_cond_10, 13'h0};
  assign mux_cond_10_pad = {6'h0,mux_cond_10_shl};
  assign mux_cond_11_shl = mux_cond_11;
  assign mux_cond_11_pad = {19'h0,mux_cond_11_shl};
  assign mux_cond_12_shl = {mux_cond_12, 7'h0};
  assign mux_cond_12_pad = {12'h0,mux_cond_12_shl};
  assign mux_cond_13_shl = {mux_cond_13, 13'h0};
  assign mux_cond_13_pad = {6'h0,mux_cond_13_shl};
  assign mux_cond_14_shl = mux_cond_14;
  assign mux_cond_14_pad = {19'h0,mux_cond_14_shl};
  assign mux_cond_15_shl = {mux_cond_15, 9'h0};
  assign mux_cond_15_pad = {10'h0,mux_cond_15_shl};
  assign mux_cond_16_shl = {mux_cond_16, 8'h0};
  assign mux_cond_16_pad = {11'h0,mux_cond_16_shl};
  assign mux_cond_17_shl = {mux_cond_17, 8'h0};
  assign mux_cond_17_pad = {11'h0,mux_cond_17_shl};
  assign mux_cond_18_shl = {mux_cond_18, 8'h0};
  assign mux_cond_18_pad = {11'h0,mux_cond_18_shl};
  assign mux_cond_19_shl = {mux_cond_19, 2'h0};
  assign mux_cond_19_pad = {17'h0,mux_cond_19_shl};
  assign mux_cond_20_shl = {mux_cond_20, 16'h0};
  assign mux_cond_20_pad = {3'h0,mux_cond_20_shl};
  assign mux_cond_21_shl = {mux_cond_21, 6'h0};
  assign mux_cond_21_pad = {13'h0,mux_cond_21_shl};
  assign mux_cond_22_shl = {mux_cond_22, 11'h0};
  assign mux_cond_22_pad = {8'h0,mux_cond_22_shl};
  assign mux_cond_23_shl = mux_cond_23;
  assign mux_cond_23_pad = {19'h0,mux_cond_23_shl};
  assign mux_cond_24_shl = {mux_cond_24, 6'h0};
  assign mux_cond_24_pad = {13'h0,mux_cond_24_shl};
  assign mux_cond_25_shl = {mux_cond_25, 12'h0};
  assign mux_cond_25_pad = {7'h0,mux_cond_25_shl};
  assign mux_cond_26_shl = {mux_cond_26, 4'h0};
  assign mux_cond_26_pad = {15'h0,mux_cond_26_shl};
  assign mux_cond_27_shl = {mux_cond_27, 11'h0};
  assign mux_cond_27_pad = {8'h0,mux_cond_27_shl};
  assign mux_cond_28_shl = {mux_cond_28, 6'h0};
  assign mux_cond_28_pad = {13'h0,mux_cond_28_shl};
  assign mux_cond_29_shl = {mux_cond_29, 12'h0};
  assign mux_cond_29_pad = {7'h0,mux_cond_29_shl};
  assign mux_cond_30_shl = {mux_cond_30, 1'h0};
  assign mux_cond_30_pad = {18'h0,mux_cond_30_shl};
  assign mux_cond_31_shl = {mux_cond_31, 11'h0};
  assign mux_cond_31_pad = {8'h0,mux_cond_31_shl};
  assign mux_cond_32_shl = {mux_cond_32, 6'h0};
  assign mux_cond_32_pad = {13'h0,mux_cond_32_shl};
  assign mux_cond_33_shl = {mux_cond_33, 5'h0};
  assign mux_cond_33_pad = {14'h0,mux_cond_33_shl};
  assign mux_cond_34_shl = {mux_cond_34, 18'h0};
  assign mux_cond_34_pad = {1'h0,mux_cond_34_shl};
  assign mux_cond_35_shl = {mux_cond_35, 12'h0};
  assign mux_cond_35_pad = {7'h0,mux_cond_35_shl};
  assign mux_cond_36_shl = mux_cond_36;
  assign mux_cond_36_pad = {19'h0,mux_cond_36_shl};
  assign mux_cond_37_shl = {mux_cond_37, 8'h0};
  assign mux_cond_37_pad = {11'h0,mux_cond_37_shl};
  assign mux_cond_38_shl = {mux_cond_38, 5'h0};
  assign mux_cond_38_pad = {14'h0,mux_cond_38_shl};
  assign mux_cond_39_shl = {mux_cond_39, 16'h0};
  assign mux_cond_39_pad = {3'h0,mux_cond_39_shl};
  assign mux_cond_40_shl = {mux_cond_40, 3'h0};
  assign mux_cond_40_pad = {16'h0,mux_cond_40_shl};
  assign mux_cond_41_shl = {mux_cond_41, 9'h0};
  assign mux_cond_41_pad = {10'h0,mux_cond_41_shl};
  assign mux_cond_42_shl = {mux_cond_42, 15'h0};
  assign mux_cond_42_pad = {4'h0,mux_cond_42_shl};
  assign mux_cond_43_shl = {mux_cond_43, 13'h0};
  assign mux_cond_43_pad = {6'h0,mux_cond_43_shl};
  assign mux_cond_44_shl = {mux_cond_44, 12'h0};
  assign mux_cond_44_pad = {7'h0,mux_cond_44_shl};
  assign mux_cond_45_shl = mux_cond_45;
  assign mux_cond_45_pad = {19'h0,mux_cond_45_shl};
  assign mux_cond_46_shl = {mux_cond_46, 3'h0};
  assign mux_cond_46_pad = {16'h0,mux_cond_46_shl};
  assign mux_cond_47_shl = {mux_cond_47, 14'h0};
  assign mux_cond_47_pad = {5'h0,mux_cond_47_shl};
  assign mux_cond_48_shl = {mux_cond_48, 16'h0};
  assign mux_cond_48_pad = {3'h0,mux_cond_48_shl};
  assign mux_cond_49_shl = {mux_cond_49, 18'h0};
  assign mux_cond_49_pad = {1'h0,mux_cond_49_shl};
  assign mux_cond_50_shl = mux_cond_50;
  assign mux_cond_50_pad = {19'h0,mux_cond_50_shl};
  assign mux_cond_51_shl = {mux_cond_51, 7'h0};
  assign mux_cond_51_pad = {12'h0,mux_cond_51_shl};
  assign mux_cond_52_shl = mux_cond_52;
  assign mux_cond_52_pad = {19'h0,mux_cond_52_shl};
  assign mux_cond_53_shl = {mux_cond_53, 19'h0};
  assign mux_cond_53_pad = mux_cond_53_shl;
  assign mux_cond_54_shl = {mux_cond_54, 10'h0};
  assign mux_cond_54_pad = {9'h0,mux_cond_54_shl};
  assign mux_cond_55_shl = {mux_cond_55, 13'h0};
  assign mux_cond_55_pad = {6'h0,mux_cond_55_shl};
  assign mux_cond_56_shl = {mux_cond_56, 9'h0};
  assign mux_cond_56_pad = {10'h0,mux_cond_56_shl};
  assign mux_cond_57_shl = {mux_cond_57, 6'h0};
  assign mux_cond_57_pad = {13'h0,mux_cond_57_shl};
  assign mux_cond_58_shl = {mux_cond_58, 17'h0};
  assign mux_cond_58_pad = {2'h0,mux_cond_58_shl};
  assign mux_cond_59_shl = {mux_cond_59, 19'h0};
  assign mux_cond_59_pad = mux_cond_59_shl;
  assign mux_cond_60_shl = {mux_cond_60, 3'h0};
  assign mux_cond_60_pad = {16'h0,mux_cond_60_shl};
  assign mux_cond_61_shl = {mux_cond_61, 14'h0};
  assign mux_cond_61_pad = {5'h0,mux_cond_61_shl};
  assign mux_cond_62_shl = {mux_cond_62, 4'h0};
  assign mux_cond_62_pad = {15'h0,mux_cond_62_shl};
  assign mux_cond_63_shl = mux_cond_63;
  assign mux_cond_63_pad = {19'h0,mux_cond_63_shl};
  assign mux_cond_64_shl = {mux_cond_64, 10'h0};
  assign mux_cond_64_pad = {9'h0,mux_cond_64_shl};
  assign mux_cond_65_shl = {mux_cond_65, 17'h0};
  assign mux_cond_65_pad = {2'h0,mux_cond_65_shl};
  assign mux_cond_66_shl = {mux_cond_66, 9'h0};
  assign mux_cond_66_pad = {10'h0,mux_cond_66_shl};
  assign mux_cond_67_shl = {mux_cond_67, 6'h0};
  assign mux_cond_67_pad = {13'h0,mux_cond_67_shl};
  assign mux_cond_68_shl = {mux_cond_68, 19'h0};
  assign mux_cond_68_pad = mux_cond_68_shl;
  assign mux_cond_69_shl = {mux_cond_69, 10'h0};
  assign mux_cond_69_pad = {9'h0,mux_cond_69_shl};
  assign mux_cond_70_shl = {mux_cond_70, 10'h0};
  assign mux_cond_70_pad = {9'h0,mux_cond_70_shl};
  assign mux_cond_71_shl = {mux_cond_71, 13'h0};
  assign mux_cond_71_pad = {6'h0,mux_cond_71_shl};
  assign mux_cond_72_shl = {mux_cond_72, 18'h0};
  assign mux_cond_72_pad = {1'h0,mux_cond_72_shl};
  assign mux_cond_73_shl = {mux_cond_73, 12'h0};
  assign mux_cond_73_pad = {7'h0,mux_cond_73_shl};
  assign mux_cond_74_shl = {mux_cond_74, 13'h0};
  assign mux_cond_74_pad = {6'h0,mux_cond_74_shl};
  assign mux_cond_75_shl = {mux_cond_75, 13'h0};
  assign mux_cond_75_pad = {6'h0,mux_cond_75_shl};
  assign mux_cond_76_shl = {mux_cond_76, 13'h0};
  assign mux_cond_76_pad = {6'h0,mux_cond_76_shl};
  assign mux_cond_77_shl = {mux_cond_77, 13'h0};
  assign mux_cond_77_pad = {6'h0,mux_cond_77_shl};
  assign mux_cond_78_shl = {mux_cond_78, 17'h0};
  assign mux_cond_78_pad = {2'h0,mux_cond_78_shl};
  assign mux_cond_79_shl = {mux_cond_79, 12'h0};
  assign mux_cond_79_pad = {7'h0,mux_cond_79_shl};
  assign mux_cond_80_shl = {mux_cond_80, 17'h0};
  assign mux_cond_80_pad = {2'h0,mux_cond_80_shl};
  assign mux_cond_81_shl = {mux_cond_81, 13'h0};
  assign mux_cond_81_pad = {6'h0,mux_cond_81_shl};
  assign mux_cond_82_shl = {mux_cond_82, 12'h0};
  assign mux_cond_82_pad = {7'h0,mux_cond_82_shl};
  assign mux_cond_83_shl = {mux_cond_83, 4'h0};
  assign mux_cond_83_pad = {15'h0,mux_cond_83_shl};
  assign mux_cond_84_shl = {mux_cond_84, 16'h0};
  assign mux_cond_84_pad = {3'h0,mux_cond_84_shl};
  assign mux_cond_85_shl = {mux_cond_85, 9'h0};
  assign mux_cond_85_pad = {10'h0,mux_cond_85_shl};
  assign mux_cond_86_shl = {mux_cond_86, 10'h0};
  assign mux_cond_86_pad = {9'h0,mux_cond_86_shl};
  assign mux_cond_87_shl = {mux_cond_87, 2'h0};
  assign mux_cond_87_pad = {17'h0,mux_cond_87_shl};
  assign mux_cond_88_shl = {mux_cond_88, 6'h0};
  assign mux_cond_88_pad = {13'h0,mux_cond_88_shl};
  assign mux_cond_89_shl = {mux_cond_89, 11'h0};
  assign mux_cond_89_pad = {8'h0,mux_cond_89_shl};
  assign mux_cond_90_shl = {mux_cond_90, 7'h0};
  assign mux_cond_90_pad = {12'h0,mux_cond_90_shl};
  assign mux_cond_91_shl = {mux_cond_91, 16'h0};
  assign mux_cond_91_pad = {3'h0,mux_cond_91_shl};
  assign mux_cond_92_shl = {mux_cond_92, 17'h0};
  assign mux_cond_92_pad = {2'h0,mux_cond_92_shl};
  assign mux_cond_93_shl = {mux_cond_93, 5'h0};
  assign mux_cond_93_pad = {14'h0,mux_cond_93_shl};
  assign mux_cond_94_shl = {mux_cond_94, 18'h0};
  assign mux_cond_94_pad = {1'h0,mux_cond_94_shl};
  assign mux_cond_95_shl = {mux_cond_95, 1'h0};
  assign mux_cond_95_pad = {18'h0,mux_cond_95_shl};
  assign mux_cond_96_shl = {mux_cond_96, 17'h0};
  assign mux_cond_96_pad = {2'h0,mux_cond_96_shl};
  assign mux_cond_97_shl = {mux_cond_97, 1'h0};
  assign mux_cond_97_pad = {18'h0,mux_cond_97_shl};
  assign MulDiv_xor64 = neg_out_pad ^ req_dw_pad;
  assign MulDiv_xor31 = isHi_pad ^ MulDiv_xor64;
  assign MulDiv_xor66 = resHi_pad ^ mux_cond_0_pad;
  assign MulDiv_xor32 = state_pad ^ MulDiv_xor66;
  assign MulDiv_xor15 = MulDiv_xor31 ^ MulDiv_xor32;
  assign MulDiv_xor68 = mux_cond_2_pad ^ mux_cond_3_pad;
  assign MulDiv_xor33 = mux_cond_1_pad ^ MulDiv_xor68;
  assign MulDiv_xor70 = mux_cond_5_pad ^ mux_cond_6_pad;
  assign MulDiv_xor34 = mux_cond_4_pad ^ MulDiv_xor70;
  assign MulDiv_xor16 = MulDiv_xor33 ^ MulDiv_xor34;
  assign MulDiv_xor7 = MulDiv_xor15 ^ MulDiv_xor16;
  assign MulDiv_xor72 = mux_cond_8_pad ^ mux_cond_9_pad;
  assign MulDiv_xor35 = mux_cond_7_pad ^ MulDiv_xor72;
  assign MulDiv_xor74 = mux_cond_11_pad ^ mux_cond_12_pad;
  assign MulDiv_xor36 = mux_cond_10_pad ^ MulDiv_xor74;
  assign MulDiv_xor17 = MulDiv_xor35 ^ MulDiv_xor36;
  assign MulDiv_xor76 = mux_cond_14_pad ^ mux_cond_15_pad;
  assign MulDiv_xor37 = mux_cond_13_pad ^ MulDiv_xor76;
  assign MulDiv_xor77 = mux_cond_16_pad ^ mux_cond_17_pad;
  assign MulDiv_xor78 = mux_cond_18_pad ^ mux_cond_19_pad;
  assign MulDiv_xor38 = MulDiv_xor77 ^ MulDiv_xor78;
  assign MulDiv_xor18 = MulDiv_xor37 ^ MulDiv_xor38;
  assign MulDiv_xor8 = MulDiv_xor17 ^ MulDiv_xor18;
  assign MulDiv_xor3 = MulDiv_xor7 ^ MulDiv_xor8;
  assign MulDiv_xor80 = mux_cond_21_pad ^ mux_cond_22_pad;
  assign MulDiv_xor39 = mux_cond_20_pad ^ MulDiv_xor80;
  assign MulDiv_xor82 = mux_cond_24_pad ^ mux_cond_25_pad;
  assign MulDiv_xor40 = mux_cond_23_pad ^ MulDiv_xor82;
  assign MulDiv_xor19 = MulDiv_xor39 ^ MulDiv_xor40;
  assign MulDiv_xor84 = mux_cond_27_pad ^ mux_cond_28_pad;
  assign MulDiv_xor41 = mux_cond_26_pad ^ MulDiv_xor84;
  assign MulDiv_xor85 = mux_cond_29_pad ^ mux_cond_30_pad;
  assign MulDiv_xor86 = mux_cond_31_pad ^ mux_cond_32_pad;
  assign MulDiv_xor42 = MulDiv_xor85 ^ MulDiv_xor86;
  assign MulDiv_xor20 = MulDiv_xor41 ^ MulDiv_xor42;
  assign MulDiv_xor9 = MulDiv_xor19 ^ MulDiv_xor20;
  assign MulDiv_xor88 = mux_cond_34_pad ^ mux_cond_35_pad;
  assign MulDiv_xor43 = mux_cond_33_pad ^ MulDiv_xor88;
  assign MulDiv_xor90 = mux_cond_37_pad ^ mux_cond_38_pad;
  assign MulDiv_xor44 = mux_cond_36_pad ^ MulDiv_xor90;
  assign MulDiv_xor21 = MulDiv_xor43 ^ MulDiv_xor44;
  assign MulDiv_xor92 = mux_cond_40_pad ^ mux_cond_41_pad;
  assign MulDiv_xor45 = mux_cond_39_pad ^ MulDiv_xor92;
  assign MulDiv_xor93 = mux_cond_42_pad ^ mux_cond_43_pad;
  assign MulDiv_xor94 = mux_cond_44_pad ^ mux_cond_45_pad;
  assign MulDiv_xor46 = MulDiv_xor93 ^ MulDiv_xor94;
  assign MulDiv_xor22 = MulDiv_xor45 ^ MulDiv_xor46;
  assign MulDiv_xor10 = MulDiv_xor21 ^ MulDiv_xor22;
  assign MulDiv_xor4 = MulDiv_xor9 ^ MulDiv_xor10;
  assign MulDiv_xor1 = MulDiv_xor3 ^ MulDiv_xor4;
  assign MulDiv_xor96 = mux_cond_47_pad ^ mux_cond_48_pad;
  assign MulDiv_xor47 = mux_cond_46_pad ^ MulDiv_xor96;
  assign MulDiv_xor98 = mux_cond_50_pad ^ mux_cond_51_pad;
  assign MulDiv_xor48 = mux_cond_49_pad ^ MulDiv_xor98;
  assign MulDiv_xor23 = MulDiv_xor47 ^ MulDiv_xor48;
  assign MulDiv_xor100 = mux_cond_53_pad ^ mux_cond_54_pad;
  assign MulDiv_xor49 = mux_cond_52_pad ^ MulDiv_xor100;
  assign MulDiv_xor101 = mux_cond_55_pad ^ mux_cond_56_pad;
  assign MulDiv_xor102 = mux_cond_57_pad ^ mux_cond_58_pad;
  assign MulDiv_xor50 = MulDiv_xor101 ^ MulDiv_xor102;
  assign MulDiv_xor24 = MulDiv_xor49 ^ MulDiv_xor50;
  assign MulDiv_xor11 = MulDiv_xor23 ^ MulDiv_xor24;
  assign MulDiv_xor104 = mux_cond_60_pad ^ mux_cond_61_pad;
  assign MulDiv_xor51 = mux_cond_59_pad ^ MulDiv_xor104;
  assign MulDiv_xor106 = mux_cond_63_pad ^ mux_cond_64_pad;
  assign MulDiv_xor52 = mux_cond_62_pad ^ MulDiv_xor106;
  assign MulDiv_xor25 = MulDiv_xor51 ^ MulDiv_xor52;
  assign MulDiv_xor108 = mux_cond_66_pad ^ mux_cond_67_pad;
  assign MulDiv_xor53 = mux_cond_65_pad ^ MulDiv_xor108;
  assign MulDiv_xor109 = mux_cond_68_pad ^ mux_cond_69_pad;
  assign MulDiv_xor110 = mux_cond_70_pad ^ mux_cond_71_pad;
  assign MulDiv_xor54 = MulDiv_xor109 ^ MulDiv_xor110;
  assign MulDiv_xor26 = MulDiv_xor53 ^ MulDiv_xor54;
  assign MulDiv_xor12 = MulDiv_xor25 ^ MulDiv_xor26;
  assign MulDiv_xor5 = MulDiv_xor11 ^ MulDiv_xor12;
  assign MulDiv_xor112 = mux_cond_73_pad ^ mux_cond_74_pad;
  assign MulDiv_xor55 = mux_cond_72_pad ^ MulDiv_xor112;
  assign MulDiv_xor114 = mux_cond_76_pad ^ mux_cond_77_pad;
  assign MulDiv_xor56 = mux_cond_75_pad ^ MulDiv_xor114;
  assign MulDiv_xor27 = MulDiv_xor55 ^ MulDiv_xor56;
  assign MulDiv_xor116 = mux_cond_79_pad ^ mux_cond_80_pad;
  assign MulDiv_xor57 = mux_cond_78_pad ^ MulDiv_xor116;
  assign MulDiv_xor117 = mux_cond_81_pad ^ mux_cond_82_pad;
  assign MulDiv_xor118 = mux_cond_83_pad ^ mux_cond_84_pad;
  assign MulDiv_xor58 = MulDiv_xor117 ^ MulDiv_xor118;
  assign MulDiv_xor28 = MulDiv_xor57 ^ MulDiv_xor58;
  assign MulDiv_xor13 = MulDiv_xor27 ^ MulDiv_xor28;
  assign MulDiv_xor120 = mux_cond_86_pad ^ mux_cond_87_pad;
  assign MulDiv_xor59 = mux_cond_85_pad ^ MulDiv_xor120;
  assign MulDiv_xor122 = mux_cond_89_pad ^ mux_cond_90_pad;
  assign MulDiv_xor60 = mux_cond_88_pad ^ MulDiv_xor122;
  assign MulDiv_xor29 = MulDiv_xor59 ^ MulDiv_xor60;
  assign MulDiv_xor124 = mux_cond_92_pad ^ mux_cond_93_pad;
  assign MulDiv_xor61 = mux_cond_91_pad ^ MulDiv_xor124;
  assign MulDiv_xor125 = mux_cond_94_pad ^ mux_cond_95_pad;
  assign MulDiv_xor126 = mux_cond_96_pad ^ mux_cond_97_pad;
  assign MulDiv_xor62 = MulDiv_xor125 ^ MulDiv_xor126;
  assign MulDiv_xor30 = MulDiv_xor61 ^ MulDiv_xor62;
  assign MulDiv_xor14 = MulDiv_xor29 ^ MulDiv_xor30;
  assign MulDiv_xor6 = MulDiv_xor13 ^ MulDiv_xor14;
  assign MulDiv_xor2 = MulDiv_xor5 ^ MulDiv_xor6;
  assign MulDiv_xor0 = MulDiv_xor1 ^ MulDiv_xor2;
  assign io_covSum = MulDiv_covSum;
  assign metaAssert = 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  req_dw = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  req_tag = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  count = _RAND_3[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  neg_out = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  isHi = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  resHi = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {3{`RANDOM}};
  divisor = _RAND_7[64:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {5{`RANDOM}};
  remainder = _RAND_8[129:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  MulDiv_state = _RAND_9[19:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1048576; initvar = initvar+1)
    MulDiv_cov[initvar] = _RAND_10[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  MulDiv_covSum = _RAND_11[29:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      state <= 3'h0;
    end else if (reset) begin
      state <= 3'h0;
    end else if (_T_36) begin
      if (cmdMul) begin
        state <= 3'h2;
      end else if (_state_T_1) begin
        state <= 3'h1;
      end else begin
        state <= 3'h3;
      end
    end else if (_T_35) begin
      state <= 3'h0;
    end else if (_T_30) begin
      if (_T_31) begin
        if (neg_out) begin
          state <= 3'h5;
        end else begin
          state <= 3'h7;
        end
      end else if (_T_27) begin
        if (_T_29) begin
          state <= 3'h6;
        end else if (_T_26) begin
          state <= 3'h7;
        end else if (_T_23) begin
          state <= 3'h3;
        end
      end else if (_T_26) begin
        state <= 3'h7;
      end else if (_T_23) begin
        state <= 3'h3;
      end
    end else if (_T_27) begin
      if (_T_29) begin
        state <= 3'h6;
      end else if (_T_26) begin
        state <= 3'h7;
      end else if (_T_23) begin
        state <= 3'h3;
      end
    end else if (_T_26) begin
      state <= 3'h7;
    end else if (_T_23) begin
      state <= 3'h3;
    end
    if (metaReset) begin
      req_dw <= 1'h0;
    end else if (_T_36) begin
      req_dw <= io_req_bits_dw;
    end
    if (metaReset) begin
      req_tag <= 5'h0;
    end else if (_T_36) begin
      req_tag <= io_req_bits_tag;
    end
    if (metaReset) begin
      count <= 7'h0;
    end else if (_T_36) begin
      count <= {{4'd0}, _count_T_8};
    end else if (_T_30) begin
      if (eOut_1) begin
        count <= {{1'd0}, eOutPos};
      end else begin
        count <= _count_T_1;
      end
    end else if (_T_27) begin
      count <= _count_T_1;
    end
    if (metaReset) begin
      neg_out <= 1'h0;
    end else if (_T_36) begin
      if (cmdHi) begin
        neg_out <= lhs_sign;
      end else begin
        neg_out <= _neg_out_T;
      end
    end else if (_T_30) begin
      if (_T_33) begin
        neg_out <= 1'h0;
      end
    end
    if (metaReset) begin
      isHi <= 1'h0;
    end else if (_T_36) begin
      isHi <= cmdHi;
    end
    if (metaReset) begin
      resHi <= 1'h0;
    end else if (_T_36) begin
      resHi <= 1'h0;
    end else if (_T_30) begin
      if (_T_31) begin
        resHi <= isHi;
      end else if (_T_27) begin
        if (_T_29) begin
          resHi <= isHi;
        end else if (_T_26) begin
          resHi <= 1'h0;
        end
      end else if (_T_26) begin
        resHi <= 1'h0;
      end
    end else if (_T_27) begin
      if (_T_29) begin
        resHi <= isHi;
      end else if (_T_26) begin
        resHi <= 1'h0;
      end
    end else if (_T_26) begin
      resHi <= 1'h0;
    end
    if (metaReset) begin
      divisor <= 65'h0;
    end else if (_T_36) begin
      divisor <= _divisor_T;
    end else if (_T_23) begin
      if (divisor[63]) begin
        divisor <= subtractor;
      end
    end
    if (metaReset) begin
      remainder <= 130'h0;
    end else if (_T_36) begin
      remainder <= {{66'd0}, lhs_in};
    end else if (_T_30) begin
      remainder <= {{1'd0}, _GEN_16};
    end else if (_T_27) begin
      remainder <= _remainder_T;
    end else if (_T_26) begin
      remainder <= {{66'd0}, negated_remainder};
    end else if (_T_23) begin
      if (remainder[63]) begin
        remainder <= {{66'd0}, negated_remainder};
      end
    end
    MulDiv_state <= MulDiv_xor0;
    if (!(MulDiv_cov_read_data)) begin
      MulDiv_covSum <= MulDiv_covSum + 1'h1;
    end
  end
  always @(posedge clock) begin
    if(MulDiv_cov_write_en & MulDiv_cov_write_mask) begin
      MulDiv_cov[MulDiv_cov_write_addr] <= MulDiv_cov_write_data; // @[Coverage map for MulDiv]
    end
  end
endmodule
module PlusArgTimeout(
  input         clock,
  input         reset,
  input  [31:0] io_count,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 62:19]
  wire  _T; // @[PlusArg.scala 63:13]
  wire  _T_1; // @[PlusArg.scala 64:22]
  wire  _T_3; // @[PlusArg.scala 64:12]
  wire [29:0] PlusArgTimeout_covSum;
  wire  stopEn0;
  wire  plusarg_reader_metaAssert_wire;
  wire  PlusArgTimeout_or0;
  reg  PlusArgTimeout_metaAssert;
  reg [31:0] _RAND_0;
//  plusarg_reader #(.FORMAT("max_core_cycles=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 62:19]
//    .out(plusarg_reader_out)
//  );
  assign _T = plusarg_reader_out > 32'h0; // @[PlusArg.scala 63:13]
  assign _T_1 = io_count < plusarg_reader_out; // @[PlusArg.scala 64:22]
  assign _T_3 = _T_1 | reset; // @[PlusArg.scala 64:12]
  assign PlusArgTimeout_covSum = 30'h0;
  assign io_covSum = PlusArgTimeout_covSum;
  assign stopEn0 = _T & ~_T_3;
//  assign plusarg_reader_metaAssert_wire = plusarg_reader_metaAssert;
  assign PlusArgTimeout_or0 = stopEn0 | plusarg_reader_metaAssert_wire;
  assign metaAssert = PlusArgTimeout_metaAssert;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  PlusArgTimeout_metaAssert = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T & ~_T_3) begin
          $fwrite(32'h80000002,"Assertion failed: Timeout exceeded: Kill the emulation after INT rdtime cycles. Off if 0.\n    at PlusArg.scala:64 assert (io.count < max, s\"Timeout exceeded: $docstring\")\n"); // @[PlusArg.scala 64:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T & ~_T_3) begin
          $fatal; // @[PlusArg.scala 64:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    if (metaReset) begin
      PlusArgTimeout_metaAssert <= 1'h0;
    end else begin
      PlusArgTimeout_metaAssert <= PlusArgTimeout_metaAssert | PlusArgTimeout_or0;
    end
  end
endmodule
module OptimizationBarrier(
  input  [19:0] io_x_ppn,
  input         io_x_u,
  input         io_x_ae,
  input         io_x_sw,
  input         io_x_sx,
  input         io_x_sr,
  input         io_x_pw,
  input         io_x_px,
  input         io_x_pr,
  input         io_x_ppp,
  input         io_x_pal,
  input         io_x_paa,
  input         io_x_eff,
  input         io_x_c,
  output [19:0] io_y_ppn,
  output        io_y_u,
  output        io_y_ae,
  output        io_y_sw,
  output        io_y_sx,
  output        io_y_sr,
  output        io_y_pw,
  output        io_y_px,
  output        io_y_pr,
  output        io_y_ppp,
  output        io_y_pal,
  output        io_y_paa,
  output        io_y_eff,
  output        io_y_c,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire [29:0] OptimizationBarrier_covSum;
  assign io_y_ppn = io_x_ppn; // @[package.scala 263:12]
  assign io_y_u = io_x_u; // @[package.scala 263:12]
  assign io_y_ae = io_x_ae; // @[package.scala 263:12]
  assign io_y_sw = io_x_sw; // @[package.scala 263:12]
  assign io_y_sx = io_x_sx; // @[package.scala 263:12]
  assign io_y_sr = io_x_sr; // @[package.scala 263:12]
  assign io_y_pw = io_x_pw; // @[package.scala 263:12]
  assign io_y_px = io_x_px; // @[package.scala 263:12]
  assign io_y_pr = io_x_pr; // @[package.scala 263:12]
  assign io_y_ppp = io_x_ppp; // @[package.scala 263:12]
  assign io_y_pal = io_x_pal; // @[package.scala 263:12]
  assign io_y_paa = io_x_paa; // @[package.scala 263:12]
  assign io_y_eff = io_x_eff; // @[package.scala 263:12]
  assign io_y_c = io_x_c; // @[package.scala 263:12]
  assign OptimizationBarrier_covSum = 30'h0;
  assign io_covSum = OptimizationBarrier_covSum;
  assign metaAssert = 1'h0;
endmodule
module PMPChecker(
  input  [1:0]  io_prv,
  input         io_pmp_0_cfg_l,
  input  [1:0]  io_pmp_0_cfg_a,
  input         io_pmp_0_cfg_x,
  input         io_pmp_0_cfg_w,
  input         io_pmp_0_cfg_r,
  input  [29:0] io_pmp_0_addr,
  input  [31:0] io_pmp_0_mask,
  input         io_pmp_1_cfg_l,
  input  [1:0]  io_pmp_1_cfg_a,
  input         io_pmp_1_cfg_x,
  input         io_pmp_1_cfg_w,
  input         io_pmp_1_cfg_r,
  input  [29:0] io_pmp_1_addr,
  input  [31:0] io_pmp_1_mask,
  input         io_pmp_2_cfg_l,
  input  [1:0]  io_pmp_2_cfg_a,
  input         io_pmp_2_cfg_x,
  input         io_pmp_2_cfg_w,
  input         io_pmp_2_cfg_r,
  input  [29:0] io_pmp_2_addr,
  input  [31:0] io_pmp_2_mask,
  input         io_pmp_3_cfg_l,
  input  [1:0]  io_pmp_3_cfg_a,
  input         io_pmp_3_cfg_x,
  input         io_pmp_3_cfg_w,
  input         io_pmp_3_cfg_r,
  input  [29:0] io_pmp_3_addr,
  input  [31:0] io_pmp_3_mask,
  input         io_pmp_4_cfg_l,
  input  [1:0]  io_pmp_4_cfg_a,
  input         io_pmp_4_cfg_x,
  input         io_pmp_4_cfg_w,
  input         io_pmp_4_cfg_r,
  input  [29:0] io_pmp_4_addr,
  input  [31:0] io_pmp_4_mask,
  input         io_pmp_5_cfg_l,
  input  [1:0]  io_pmp_5_cfg_a,
  input         io_pmp_5_cfg_x,
  input         io_pmp_5_cfg_w,
  input         io_pmp_5_cfg_r,
  input  [29:0] io_pmp_5_addr,
  input  [31:0] io_pmp_5_mask,
  input         io_pmp_6_cfg_l,
  input  [1:0]  io_pmp_6_cfg_a,
  input         io_pmp_6_cfg_x,
  input         io_pmp_6_cfg_w,
  input         io_pmp_6_cfg_r,
  input  [29:0] io_pmp_6_addr,
  input  [31:0] io_pmp_6_mask,
  input         io_pmp_7_cfg_l,
  input  [1:0]  io_pmp_7_cfg_a,
  input         io_pmp_7_cfg_x,
  input         io_pmp_7_cfg_w,
  input         io_pmp_7_cfg_r,
  input  [29:0] io_pmp_7_addr,
  input  [31:0] io_pmp_7_mask,
  input  [31:0] io_addr,
  input  [1:0]  io_size,
  output        io_r,
  output        io_w,
  output        io_x,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  default_; // @[PMP.scala 157:56]
  wire [5:0] _res_hit_lsbMask_T_1; // @[package.scala 234:77]
  wire [31:0] _GEN_0; // @[PMP.scala 70:26]
  wire [31:0] res_hit_lsbMask; // @[PMP.scala 70:26]
  wire [31:0] _res_hit_msbMatch_T_1; // @[PMP.scala 62:36]
  wire [31:0] _res_hit_msbMatch_T_3; // @[PMP.scala 62:48]
  wire [28:0] _res_hit_msbMatch_T_5; // @[PMP.scala 71:53]
  wire [28:0] _res_hit_msbMatch_T_7; // @[PMP.scala 65:47]
  wire [28:0] _res_hit_msbMatch_T_9; // @[PMP.scala 65:52]
  wire  res_hit_msbMatch; // @[PMP.scala 65:58]
  wire [2:0] _res_hit_lsbMatch_T_5; // @[PMP.scala 72:55]
  wire [2:0] _res_hit_lsbMatch_T_7; // @[PMP.scala 65:47]
  wire [2:0] _res_hit_lsbMatch_T_9; // @[PMP.scala 65:52]
  wire  res_hit_lsbMatch; // @[PMP.scala 65:58]
  wire  _res_hit_T_1; // @[PMP.scala 73:16]
  wire [31:0] _res_hit_msbsLess_T_1; // @[PMP.scala 62:36]
  wire [31:0] _res_hit_msbsLess_T_3; // @[PMP.scala 62:48]
  wire [28:0] _res_hit_msbsLess_T_5; // @[PMP.scala 82:52]
  wire  res_hit_msbsLess; // @[PMP.scala 82:39]
  wire [28:0] _res_hit_msbsEqual_T_6; // @[PMP.scala 83:41]
  wire  res_hit_msbsEqual; // @[PMP.scala 83:69]
  wire [2:0] _res_hit_lsbsLess_T_1; // @[PMP.scala 84:42]
  wire [2:0] _res_hit_lsbsLess_T_6; // @[PMP.scala 84:64]
  wire  res_hit_lsbsLess; // @[PMP.scala 84:53]
  wire  _res_hit_T_7; // @[PMP.scala 85:30]
  wire  _res_hit_T_8; // @[PMP.scala 85:16]
  wire  res_hit_msbsLess_1; // @[PMP.scala 82:39]
  wire  res_hit_msbsEqual_1; // @[PMP.scala 83:69]
  wire  res_hit_lsbsLess_1; // @[PMP.scala 84:53]
  wire  _res_hit_T_10; // @[PMP.scala 85:30]
  wire  _res_hit_T_11; // @[PMP.scala 85:16]
  wire  _res_hit_T_12; // @[PMP.scala 96:48]
  wire  _res_hit_T_13; // @[PMP.scala 134:61]
  wire  res_hit; // @[PMP.scala 134:8]
  wire  res_ignore; // @[PMP.scala 165:26]
  wire [2:0] _res_aligned_straddlesLowerBound_T_15; // @[PMP.scala 125:123]
  wire  _res_aligned_straddlesLowerBound_T_16; // @[PMP.scala 125:145]
  wire  res_aligned_straddlesLowerBound; // @[PMP.scala 125:88]
  wire [2:0] _res_aligned_straddlesUpperBound_T_15; // @[PMP.scala 126:113]
  wire  _res_aligned_straddlesUpperBound_T_16; // @[PMP.scala 126:146]
  wire  res_aligned_straddlesUpperBound; // @[PMP.scala 126:83]
  wire  _res_aligned_rangeAligned_T; // @[PMP.scala 127:46]
  wire  res_aligned_rangeAligned; // @[PMP.scala 127:24]
  wire [2:0] _res_aligned_pow2Aligned_T_2; // @[PMP.scala 128:32]
  wire  res_aligned_pow2Aligned; // @[PMP.scala 128:57]
  wire  res_aligned; // @[PMP.scala 129:8]
  wire  _res_cur_cfg_r_T; // @[PMP.scala 183:40]
  wire  res_cur_cfg_r; // @[PMP.scala 183:26]
  wire  _res_cur_cfg_w_T; // @[PMP.scala 184:40]
  wire  res_cur_cfg_w; // @[PMP.scala 184:26]
  wire  _res_cur_cfg_x_T; // @[PMP.scala 185:40]
  wire  res_cur_cfg_x; // @[PMP.scala 185:26]
  wire  _res_T_44_cfg_x; // @[PMP.scala 186:8]
  wire  _res_T_44_cfg_w; // @[PMP.scala 186:8]
  wire  _res_T_44_cfg_r; // @[PMP.scala 186:8]
  wire [31:0] res_hit_lsbMask_1; // @[PMP.scala 70:26]
  wire [28:0] _res_hit_msbMatch_T_19; // @[PMP.scala 65:52]
  wire  res_hit_msbMatch_1; // @[PMP.scala 65:58]
  wire [2:0] _res_hit_lsbMatch_T_17; // @[PMP.scala 65:47]
  wire [2:0] _res_hit_lsbMatch_T_19; // @[PMP.scala 65:52]
  wire  res_hit_lsbMatch_1; // @[PMP.scala 65:58]
  wire  _res_hit_T_15; // @[PMP.scala 73:16]
  wire [31:0] _res_hit_msbsLess_T_13; // @[PMP.scala 62:36]
  wire [31:0] _res_hit_msbsLess_T_15; // @[PMP.scala 62:48]
  wire [28:0] _res_hit_msbsLess_T_17; // @[PMP.scala 82:52]
  wire  res_hit_msbsLess_2; // @[PMP.scala 82:39]
  wire [28:0] _res_hit_msbsEqual_T_20; // @[PMP.scala 83:41]
  wire  res_hit_msbsEqual_2; // @[PMP.scala 83:69]
  wire [2:0] _res_hit_lsbsLess_T_20; // @[PMP.scala 84:64]
  wire  res_hit_lsbsLess_2; // @[PMP.scala 84:53]
  wire  _res_hit_T_21; // @[PMP.scala 85:30]
  wire  _res_hit_T_22; // @[PMP.scala 85:16]
  wire  res_hit_lsbsLess_3; // @[PMP.scala 84:53]
  wire  _res_hit_T_24; // @[PMP.scala 85:30]
  wire  _res_hit_T_25; // @[PMP.scala 85:16]
  wire  _res_hit_T_26; // @[PMP.scala 96:48]
  wire  _res_hit_T_27; // @[PMP.scala 134:61]
  wire  res_hit_1; // @[PMP.scala 134:8]
  wire  res_ignore_1; // @[PMP.scala 165:26]
  wire [2:0] _res_aligned_straddlesLowerBound_T_32; // @[PMP.scala 125:123]
  wire  _res_aligned_straddlesLowerBound_T_33; // @[PMP.scala 125:145]
  wire  res_aligned_straddlesLowerBound_1; // @[PMP.scala 125:88]
  wire [2:0] _res_aligned_straddlesUpperBound_T_32; // @[PMP.scala 126:113]
  wire  _res_aligned_straddlesUpperBound_T_33; // @[PMP.scala 126:146]
  wire  res_aligned_straddlesUpperBound_1; // @[PMP.scala 126:83]
  wire  _res_aligned_rangeAligned_T_1; // @[PMP.scala 127:46]
  wire  res_aligned_rangeAligned_1; // @[PMP.scala 127:24]
  wire [2:0] _res_aligned_pow2Aligned_T_5; // @[PMP.scala 128:32]
  wire  res_aligned_pow2Aligned_1; // @[PMP.scala 128:57]
  wire  res_aligned_1; // @[PMP.scala 129:8]
  wire  _res_cur_cfg_r_T_2; // @[PMP.scala 183:40]
  wire  res_cur_1_cfg_r; // @[PMP.scala 183:26]
  wire  _res_cur_cfg_w_T_2; // @[PMP.scala 184:40]
  wire  res_cur_1_cfg_w; // @[PMP.scala 184:26]
  wire  _res_cur_cfg_x_T_2; // @[PMP.scala 185:40]
  wire  res_cur_1_cfg_x; // @[PMP.scala 185:26]
  wire  _res_T_89_cfg_x; // @[PMP.scala 186:8]
  wire  _res_T_89_cfg_w; // @[PMP.scala 186:8]
  wire  _res_T_89_cfg_r; // @[PMP.scala 186:8]
  wire [31:0] res_hit_lsbMask_2; // @[PMP.scala 70:26]
  wire [28:0] _res_hit_msbMatch_T_29; // @[PMP.scala 65:52]
  wire  res_hit_msbMatch_2; // @[PMP.scala 65:58]
  wire [2:0] _res_hit_lsbMatch_T_27; // @[PMP.scala 65:47]
  wire [2:0] _res_hit_lsbMatch_T_29; // @[PMP.scala 65:52]
  wire  res_hit_lsbMatch_2; // @[PMP.scala 65:58]
  wire  _res_hit_T_29; // @[PMP.scala 73:16]
  wire [31:0] _res_hit_msbsLess_T_25; // @[PMP.scala 62:36]
  wire [31:0] _res_hit_msbsLess_T_27; // @[PMP.scala 62:48]
  wire [28:0] _res_hit_msbsLess_T_29; // @[PMP.scala 82:52]
  wire  res_hit_msbsLess_4; // @[PMP.scala 82:39]
  wire [28:0] _res_hit_msbsEqual_T_34; // @[PMP.scala 83:41]
  wire  res_hit_msbsEqual_4; // @[PMP.scala 83:69]
  wire [2:0] _res_hit_lsbsLess_T_34; // @[PMP.scala 84:64]
  wire  res_hit_lsbsLess_4; // @[PMP.scala 84:53]
  wire  _res_hit_T_35; // @[PMP.scala 85:30]
  wire  _res_hit_T_36; // @[PMP.scala 85:16]
  wire  res_hit_lsbsLess_5; // @[PMP.scala 84:53]
  wire  _res_hit_T_38; // @[PMP.scala 85:30]
  wire  _res_hit_T_39; // @[PMP.scala 85:16]
  wire  _res_hit_T_40; // @[PMP.scala 96:48]
  wire  _res_hit_T_41; // @[PMP.scala 134:61]
  wire  res_hit_2; // @[PMP.scala 134:8]
  wire  res_ignore_2; // @[PMP.scala 165:26]
  wire [2:0] _res_aligned_straddlesLowerBound_T_49; // @[PMP.scala 125:123]
  wire  _res_aligned_straddlesLowerBound_T_50; // @[PMP.scala 125:145]
  wire  res_aligned_straddlesLowerBound_2; // @[PMP.scala 125:88]
  wire [2:0] _res_aligned_straddlesUpperBound_T_49; // @[PMP.scala 126:113]
  wire  _res_aligned_straddlesUpperBound_T_50; // @[PMP.scala 126:146]
  wire  res_aligned_straddlesUpperBound_2; // @[PMP.scala 126:83]
  wire  _res_aligned_rangeAligned_T_2; // @[PMP.scala 127:46]
  wire  res_aligned_rangeAligned_2; // @[PMP.scala 127:24]
  wire [2:0] _res_aligned_pow2Aligned_T_8; // @[PMP.scala 128:32]
  wire  res_aligned_pow2Aligned_2; // @[PMP.scala 128:57]
  wire  res_aligned_2; // @[PMP.scala 129:8]
  wire  _res_cur_cfg_r_T_4; // @[PMP.scala 183:40]
  wire  res_cur_2_cfg_r; // @[PMP.scala 183:26]
  wire  _res_cur_cfg_w_T_4; // @[PMP.scala 184:40]
  wire  res_cur_2_cfg_w; // @[PMP.scala 184:26]
  wire  _res_cur_cfg_x_T_4; // @[PMP.scala 185:40]
  wire  res_cur_2_cfg_x; // @[PMP.scala 185:26]
  wire  _res_T_134_cfg_x; // @[PMP.scala 186:8]
  wire  _res_T_134_cfg_w; // @[PMP.scala 186:8]
  wire  _res_T_134_cfg_r; // @[PMP.scala 186:8]
  wire [31:0] res_hit_lsbMask_3; // @[PMP.scala 70:26]
  wire [28:0] _res_hit_msbMatch_T_39; // @[PMP.scala 65:52]
  wire  res_hit_msbMatch_3; // @[PMP.scala 65:58]
  wire [2:0] _res_hit_lsbMatch_T_37; // @[PMP.scala 65:47]
  wire [2:0] _res_hit_lsbMatch_T_39; // @[PMP.scala 65:52]
  wire  res_hit_lsbMatch_3; // @[PMP.scala 65:58]
  wire  _res_hit_T_43; // @[PMP.scala 73:16]
  wire [31:0] _res_hit_msbsLess_T_37; // @[PMP.scala 62:36]
  wire [31:0] _res_hit_msbsLess_T_39; // @[PMP.scala 62:48]
  wire [28:0] _res_hit_msbsLess_T_41; // @[PMP.scala 82:52]
  wire  res_hit_msbsLess_6; // @[PMP.scala 82:39]
  wire [28:0] _res_hit_msbsEqual_T_48; // @[PMP.scala 83:41]
  wire  res_hit_msbsEqual_6; // @[PMP.scala 83:69]
  wire [2:0] _res_hit_lsbsLess_T_48; // @[PMP.scala 84:64]
  wire  res_hit_lsbsLess_6; // @[PMP.scala 84:53]
  wire  _res_hit_T_49; // @[PMP.scala 85:30]
  wire  _res_hit_T_50; // @[PMP.scala 85:16]
  wire  res_hit_lsbsLess_7; // @[PMP.scala 84:53]
  wire  _res_hit_T_52; // @[PMP.scala 85:30]
  wire  _res_hit_T_53; // @[PMP.scala 85:16]
  wire  _res_hit_T_54; // @[PMP.scala 96:48]
  wire  _res_hit_T_55; // @[PMP.scala 134:61]
  wire  res_hit_3; // @[PMP.scala 134:8]
  wire  res_ignore_3; // @[PMP.scala 165:26]
  wire [2:0] _res_aligned_straddlesLowerBound_T_66; // @[PMP.scala 125:123]
  wire  _res_aligned_straddlesLowerBound_T_67; // @[PMP.scala 125:145]
  wire  res_aligned_straddlesLowerBound_3; // @[PMP.scala 125:88]
  wire [2:0] _res_aligned_straddlesUpperBound_T_66; // @[PMP.scala 126:113]
  wire  _res_aligned_straddlesUpperBound_T_67; // @[PMP.scala 126:146]
  wire  res_aligned_straddlesUpperBound_3; // @[PMP.scala 126:83]
  wire  _res_aligned_rangeAligned_T_3; // @[PMP.scala 127:46]
  wire  res_aligned_rangeAligned_3; // @[PMP.scala 127:24]
  wire [2:0] _res_aligned_pow2Aligned_T_11; // @[PMP.scala 128:32]
  wire  res_aligned_pow2Aligned_3; // @[PMP.scala 128:57]
  wire  res_aligned_3; // @[PMP.scala 129:8]
  wire  _res_cur_cfg_r_T_6; // @[PMP.scala 183:40]
  wire  res_cur_3_cfg_r; // @[PMP.scala 183:26]
  wire  _res_cur_cfg_w_T_6; // @[PMP.scala 184:40]
  wire  res_cur_3_cfg_w; // @[PMP.scala 184:26]
  wire  _res_cur_cfg_x_T_6; // @[PMP.scala 185:40]
  wire  res_cur_3_cfg_x; // @[PMP.scala 185:26]
  wire  _res_T_179_cfg_x; // @[PMP.scala 186:8]
  wire  _res_T_179_cfg_w; // @[PMP.scala 186:8]
  wire  _res_T_179_cfg_r; // @[PMP.scala 186:8]
  wire [31:0] res_hit_lsbMask_4; // @[PMP.scala 70:26]
  wire [28:0] _res_hit_msbMatch_T_49; // @[PMP.scala 65:52]
  wire  res_hit_msbMatch_4; // @[PMP.scala 65:58]
  wire [2:0] _res_hit_lsbMatch_T_47; // @[PMP.scala 65:47]
  wire [2:0] _res_hit_lsbMatch_T_49; // @[PMP.scala 65:52]
  wire  res_hit_lsbMatch_4; // @[PMP.scala 65:58]
  wire  _res_hit_T_57; // @[PMP.scala 73:16]
  wire [31:0] _res_hit_msbsLess_T_49; // @[PMP.scala 62:36]
  wire [31:0] _res_hit_msbsLess_T_51; // @[PMP.scala 62:48]
  wire [28:0] _res_hit_msbsLess_T_53; // @[PMP.scala 82:52]
  wire  res_hit_msbsLess_8; // @[PMP.scala 82:39]
  wire [28:0] _res_hit_msbsEqual_T_62; // @[PMP.scala 83:41]
  wire  res_hit_msbsEqual_8; // @[PMP.scala 83:69]
  wire [2:0] _res_hit_lsbsLess_T_62; // @[PMP.scala 84:64]
  wire  res_hit_lsbsLess_8; // @[PMP.scala 84:53]
  wire  _res_hit_T_63; // @[PMP.scala 85:30]
  wire  _res_hit_T_64; // @[PMP.scala 85:16]
  wire  res_hit_lsbsLess_9; // @[PMP.scala 84:53]
  wire  _res_hit_T_66; // @[PMP.scala 85:30]
  wire  _res_hit_T_67; // @[PMP.scala 85:16]
  wire  _res_hit_T_68; // @[PMP.scala 96:48]
  wire  _res_hit_T_69; // @[PMP.scala 134:61]
  wire  res_hit_4; // @[PMP.scala 134:8]
  wire  res_ignore_4; // @[PMP.scala 165:26]
  wire [2:0] _res_aligned_straddlesLowerBound_T_83; // @[PMP.scala 125:123]
  wire  _res_aligned_straddlesLowerBound_T_84; // @[PMP.scala 125:145]
  wire  res_aligned_straddlesLowerBound_4; // @[PMP.scala 125:88]
  wire [2:0] _res_aligned_straddlesUpperBound_T_83; // @[PMP.scala 126:113]
  wire  _res_aligned_straddlesUpperBound_T_84; // @[PMP.scala 126:146]
  wire  res_aligned_straddlesUpperBound_4; // @[PMP.scala 126:83]
  wire  _res_aligned_rangeAligned_T_4; // @[PMP.scala 127:46]
  wire  res_aligned_rangeAligned_4; // @[PMP.scala 127:24]
  wire [2:0] _res_aligned_pow2Aligned_T_14; // @[PMP.scala 128:32]
  wire  res_aligned_pow2Aligned_4; // @[PMP.scala 128:57]
  wire  res_aligned_4; // @[PMP.scala 129:8]
  wire  _res_cur_cfg_r_T_8; // @[PMP.scala 183:40]
  wire  res_cur_4_cfg_r; // @[PMP.scala 183:26]
  wire  _res_cur_cfg_w_T_8; // @[PMP.scala 184:40]
  wire  res_cur_4_cfg_w; // @[PMP.scala 184:26]
  wire  _res_cur_cfg_x_T_8; // @[PMP.scala 185:40]
  wire  res_cur_4_cfg_x; // @[PMP.scala 185:26]
  wire  _res_T_224_cfg_x; // @[PMP.scala 186:8]
  wire  _res_T_224_cfg_w; // @[PMP.scala 186:8]
  wire  _res_T_224_cfg_r; // @[PMP.scala 186:8]
  wire [31:0] res_hit_lsbMask_5; // @[PMP.scala 70:26]
  wire [28:0] _res_hit_msbMatch_T_59; // @[PMP.scala 65:52]
  wire  res_hit_msbMatch_5; // @[PMP.scala 65:58]
  wire [2:0] _res_hit_lsbMatch_T_57; // @[PMP.scala 65:47]
  wire [2:0] _res_hit_lsbMatch_T_59; // @[PMP.scala 65:52]
  wire  res_hit_lsbMatch_5; // @[PMP.scala 65:58]
  wire  _res_hit_T_71; // @[PMP.scala 73:16]
  wire [31:0] _res_hit_msbsLess_T_61; // @[PMP.scala 62:36]
  wire [31:0] _res_hit_msbsLess_T_63; // @[PMP.scala 62:48]
  wire [28:0] _res_hit_msbsLess_T_65; // @[PMP.scala 82:52]
  wire  res_hit_msbsLess_10; // @[PMP.scala 82:39]
  wire [28:0] _res_hit_msbsEqual_T_76; // @[PMP.scala 83:41]
  wire  res_hit_msbsEqual_10; // @[PMP.scala 83:69]
  wire [2:0] _res_hit_lsbsLess_T_76; // @[PMP.scala 84:64]
  wire  res_hit_lsbsLess_10; // @[PMP.scala 84:53]
  wire  _res_hit_T_77; // @[PMP.scala 85:30]
  wire  _res_hit_T_78; // @[PMP.scala 85:16]
  wire  res_hit_lsbsLess_11; // @[PMP.scala 84:53]
  wire  _res_hit_T_80; // @[PMP.scala 85:30]
  wire  _res_hit_T_81; // @[PMP.scala 85:16]
  wire  _res_hit_T_82; // @[PMP.scala 96:48]
  wire  _res_hit_T_83; // @[PMP.scala 134:61]
  wire  res_hit_5; // @[PMP.scala 134:8]
  wire  res_ignore_5; // @[PMP.scala 165:26]
  wire [2:0] _res_aligned_straddlesLowerBound_T_100; // @[PMP.scala 125:123]
  wire  _res_aligned_straddlesLowerBound_T_101; // @[PMP.scala 125:145]
  wire  res_aligned_straddlesLowerBound_5; // @[PMP.scala 125:88]
  wire [2:0] _res_aligned_straddlesUpperBound_T_100; // @[PMP.scala 126:113]
  wire  _res_aligned_straddlesUpperBound_T_101; // @[PMP.scala 126:146]
  wire  res_aligned_straddlesUpperBound_5; // @[PMP.scala 126:83]
  wire  _res_aligned_rangeAligned_T_5; // @[PMP.scala 127:46]
  wire  res_aligned_rangeAligned_5; // @[PMP.scala 127:24]
  wire [2:0] _res_aligned_pow2Aligned_T_17; // @[PMP.scala 128:32]
  wire  res_aligned_pow2Aligned_5; // @[PMP.scala 128:57]
  wire  res_aligned_5; // @[PMP.scala 129:8]
  wire  _res_cur_cfg_r_T_10; // @[PMP.scala 183:40]
  wire  res_cur_5_cfg_r; // @[PMP.scala 183:26]
  wire  _res_cur_cfg_w_T_10; // @[PMP.scala 184:40]
  wire  res_cur_5_cfg_w; // @[PMP.scala 184:26]
  wire  _res_cur_cfg_x_T_10; // @[PMP.scala 185:40]
  wire  res_cur_5_cfg_x; // @[PMP.scala 185:26]
  wire  _res_T_269_cfg_x; // @[PMP.scala 186:8]
  wire  _res_T_269_cfg_w; // @[PMP.scala 186:8]
  wire  _res_T_269_cfg_r; // @[PMP.scala 186:8]
  wire [31:0] res_hit_lsbMask_6; // @[PMP.scala 70:26]
  wire [28:0] _res_hit_msbMatch_T_69; // @[PMP.scala 65:52]
  wire  res_hit_msbMatch_6; // @[PMP.scala 65:58]
  wire [2:0] _res_hit_lsbMatch_T_67; // @[PMP.scala 65:47]
  wire [2:0] _res_hit_lsbMatch_T_69; // @[PMP.scala 65:52]
  wire  res_hit_lsbMatch_6; // @[PMP.scala 65:58]
  wire  _res_hit_T_85; // @[PMP.scala 73:16]
  wire [31:0] _res_hit_msbsLess_T_73; // @[PMP.scala 62:36]
  wire [31:0] _res_hit_msbsLess_T_75; // @[PMP.scala 62:48]
  wire [28:0] _res_hit_msbsLess_T_77; // @[PMP.scala 82:52]
  wire  res_hit_msbsLess_12; // @[PMP.scala 82:39]
  wire [28:0] _res_hit_msbsEqual_T_90; // @[PMP.scala 83:41]
  wire  res_hit_msbsEqual_12; // @[PMP.scala 83:69]
  wire [2:0] _res_hit_lsbsLess_T_90; // @[PMP.scala 84:64]
  wire  res_hit_lsbsLess_12; // @[PMP.scala 84:53]
  wire  _res_hit_T_91; // @[PMP.scala 85:30]
  wire  _res_hit_T_92; // @[PMP.scala 85:16]
  wire  res_hit_lsbsLess_13; // @[PMP.scala 84:53]
  wire  _res_hit_T_94; // @[PMP.scala 85:30]
  wire  _res_hit_T_95; // @[PMP.scala 85:16]
  wire  _res_hit_T_96; // @[PMP.scala 96:48]
  wire  _res_hit_T_97; // @[PMP.scala 134:61]
  wire  res_hit_6; // @[PMP.scala 134:8]
  wire  res_ignore_6; // @[PMP.scala 165:26]
  wire [2:0] _res_aligned_straddlesLowerBound_T_117; // @[PMP.scala 125:123]
  wire  _res_aligned_straddlesLowerBound_T_118; // @[PMP.scala 125:145]
  wire  res_aligned_straddlesLowerBound_6; // @[PMP.scala 125:88]
  wire [2:0] _res_aligned_straddlesUpperBound_T_117; // @[PMP.scala 126:113]
  wire  _res_aligned_straddlesUpperBound_T_118; // @[PMP.scala 126:146]
  wire  res_aligned_straddlesUpperBound_6; // @[PMP.scala 126:83]
  wire  _res_aligned_rangeAligned_T_6; // @[PMP.scala 127:46]
  wire  res_aligned_rangeAligned_6; // @[PMP.scala 127:24]
  wire [2:0] _res_aligned_pow2Aligned_T_20; // @[PMP.scala 128:32]
  wire  res_aligned_pow2Aligned_6; // @[PMP.scala 128:57]
  wire  res_aligned_6; // @[PMP.scala 129:8]
  wire  _res_cur_cfg_r_T_12; // @[PMP.scala 183:40]
  wire  res_cur_6_cfg_r; // @[PMP.scala 183:26]
  wire  _res_cur_cfg_w_T_12; // @[PMP.scala 184:40]
  wire  res_cur_6_cfg_w; // @[PMP.scala 184:26]
  wire  _res_cur_cfg_x_T_12; // @[PMP.scala 185:40]
  wire  res_cur_6_cfg_x; // @[PMP.scala 185:26]
  wire  _res_T_314_cfg_x; // @[PMP.scala 186:8]
  wire  _res_T_314_cfg_w; // @[PMP.scala 186:8]
  wire  _res_T_314_cfg_r; // @[PMP.scala 186:8]
  wire [31:0] res_hit_lsbMask_7; // @[PMP.scala 70:26]
  wire [28:0] _res_hit_msbMatch_T_79; // @[PMP.scala 65:52]
  wire  res_hit_msbMatch_7; // @[PMP.scala 65:58]
  wire [2:0] _res_hit_lsbMatch_T_77; // @[PMP.scala 65:47]
  wire [2:0] _res_hit_lsbMatch_T_79; // @[PMP.scala 65:52]
  wire  res_hit_lsbMatch_7; // @[PMP.scala 65:58]
  wire  _res_hit_T_99; // @[PMP.scala 73:16]
  wire  res_hit_lsbsLess_15; // @[PMP.scala 84:53]
  wire  _res_hit_T_108; // @[PMP.scala 85:30]
  wire  _res_hit_T_109; // @[PMP.scala 85:16]
  wire  _res_hit_T_111; // @[PMP.scala 134:61]
  wire  res_hit_7; // @[PMP.scala 134:8]
  wire  res_ignore_7; // @[PMP.scala 165:26]
  wire [2:0] _res_aligned_straddlesUpperBound_T_134; // @[PMP.scala 126:113]
  wire  _res_aligned_straddlesUpperBound_T_135; // @[PMP.scala 126:146]
  wire  res_aligned_straddlesUpperBound_7; // @[PMP.scala 126:83]
  wire  res_aligned_rangeAligned_7; // @[PMP.scala 127:24]
  wire [2:0] _res_aligned_pow2Aligned_T_23; // @[PMP.scala 128:32]
  wire  res_aligned_pow2Aligned_7; // @[PMP.scala 128:57]
  wire  res_aligned_7; // @[PMP.scala 129:8]
  wire  _res_cur_cfg_r_T_14; // @[PMP.scala 183:40]
  wire  res_cur_7_cfg_r; // @[PMP.scala 183:26]
  wire  _res_cur_cfg_w_T_14; // @[PMP.scala 184:40]
  wire  res_cur_7_cfg_w; // @[PMP.scala 184:26]
  wire  _res_cur_cfg_x_T_14; // @[PMP.scala 185:40]
  wire  res_cur_7_cfg_x; // @[PMP.scala 185:26]
  wire [29:0] PMPChecker_covSum;
  assign default_ = io_prv > 2'h1; // @[PMP.scala 157:56]
  assign _res_hit_lsbMask_T_1 = 6'h7 << io_size; // @[package.scala 234:77]
  assign _GEN_0 = {{29'd0}, ~_res_hit_lsbMask_T_1[2:0]}; // @[PMP.scala 70:26]
  assign res_hit_lsbMask = io_pmp_7_mask | _GEN_0; // @[PMP.scala 70:26]
  assign _res_hit_msbMatch_T_1 = {io_pmp_7_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _res_hit_msbMatch_T_3 = ~_res_hit_msbMatch_T_1 | 32'h3; // @[PMP.scala 62:48]
  assign _res_hit_msbMatch_T_5 = ~_res_hit_msbMatch_T_3[31:3]; // @[PMP.scala 71:53]
  assign _res_hit_msbMatch_T_7 = io_addr[31:3] ^ _res_hit_msbMatch_T_5; // @[PMP.scala 65:47]
  assign _res_hit_msbMatch_T_9 = _res_hit_msbMatch_T_7 & ~io_pmp_7_mask[31:3]; // @[PMP.scala 65:52]
  assign res_hit_msbMatch = _res_hit_msbMatch_T_9 == 29'h0; // @[PMP.scala 65:58]
  assign _res_hit_lsbMatch_T_5 = ~_res_hit_msbMatch_T_3[2:0]; // @[PMP.scala 72:55]
  assign _res_hit_lsbMatch_T_7 = io_addr[2:0] ^ _res_hit_lsbMatch_T_5; // @[PMP.scala 65:47]
  assign _res_hit_lsbMatch_T_9 = _res_hit_lsbMatch_T_7 & ~res_hit_lsbMask[2:0]; // @[PMP.scala 65:52]
  assign res_hit_lsbMatch = _res_hit_lsbMatch_T_9 == 3'h0; // @[PMP.scala 65:58]
  assign _res_hit_T_1 = res_hit_msbMatch & res_hit_lsbMatch; // @[PMP.scala 73:16]
  assign _res_hit_msbsLess_T_1 = {io_pmp_6_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _res_hit_msbsLess_T_3 = ~_res_hit_msbsLess_T_1 | 32'h3; // @[PMP.scala 62:48]
  assign _res_hit_msbsLess_T_5 = ~_res_hit_msbsLess_T_3[31:3]; // @[PMP.scala 82:52]
  assign res_hit_msbsLess = io_addr[31:3] < _res_hit_msbsLess_T_5; // @[PMP.scala 82:39]
  assign _res_hit_msbsEqual_T_6 = io_addr[31:3] ^ _res_hit_msbsLess_T_5; // @[PMP.scala 83:41]
  assign res_hit_msbsEqual = _res_hit_msbsEqual_T_6 == 29'h0; // @[PMP.scala 83:69]
  assign _res_hit_lsbsLess_T_1 = io_addr[2:0] | ~_res_hit_lsbMask_T_1[2:0]; // @[PMP.scala 84:42]
  assign _res_hit_lsbsLess_T_6 = ~_res_hit_msbsLess_T_3[2:0]; // @[PMP.scala 84:64]
  assign res_hit_lsbsLess = _res_hit_lsbsLess_T_1 < _res_hit_lsbsLess_T_6; // @[PMP.scala 84:53]
  assign _res_hit_T_7 = res_hit_msbsEqual & res_hit_lsbsLess; // @[PMP.scala 85:30]
  assign _res_hit_T_8 = res_hit_msbsLess | _res_hit_T_7; // @[PMP.scala 85:16]
  assign res_hit_msbsLess_1 = io_addr[31:3] < _res_hit_msbMatch_T_5; // @[PMP.scala 82:39]
  assign res_hit_msbsEqual_1 = _res_hit_msbMatch_T_7 == 29'h0; // @[PMP.scala 83:69]
  assign res_hit_lsbsLess_1 = io_addr[2:0] < _res_hit_lsbMatch_T_5; // @[PMP.scala 84:53]
  assign _res_hit_T_10 = res_hit_msbsEqual_1 & res_hit_lsbsLess_1; // @[PMP.scala 85:30]
  assign _res_hit_T_11 = res_hit_msbsLess_1 | _res_hit_T_10; // @[PMP.scala 85:16]
  assign _res_hit_T_12 = ~_res_hit_T_8 & _res_hit_T_11; // @[PMP.scala 96:48]
  assign _res_hit_T_13 = io_pmp_7_cfg_a[0] & _res_hit_T_12; // @[PMP.scala 134:61]
  assign res_hit = io_pmp_7_cfg_a[1] ? _res_hit_T_1 : _res_hit_T_13; // @[PMP.scala 134:8]
  assign res_ignore = default_ & ~io_pmp_7_cfg_l; // @[PMP.scala 165:26]
  assign _res_aligned_straddlesLowerBound_T_15 = _res_hit_lsbsLess_T_6 & ~io_addr[2:0]; // @[PMP.scala 125:123]
  assign _res_aligned_straddlesLowerBound_T_16 = _res_aligned_straddlesLowerBound_T_15 != 3'h0; // @[PMP.scala 125:145]
  assign res_aligned_straddlesLowerBound = res_hit_msbsEqual & _res_aligned_straddlesLowerBound_T_16; // @[PMP.scala 125:88]
  assign _res_aligned_straddlesUpperBound_T_15 = _res_hit_lsbMatch_T_5 & _res_hit_lsbsLess_T_1; // @[PMP.scala 126:113]
  assign _res_aligned_straddlesUpperBound_T_16 = _res_aligned_straddlesUpperBound_T_15 != 3'h0; // @[PMP.scala 126:146]
  assign res_aligned_straddlesUpperBound = res_hit_msbsEqual_1 & _res_aligned_straddlesUpperBound_T_16; // @[PMP.scala 126:83]
  assign _res_aligned_rangeAligned_T = res_aligned_straddlesLowerBound | res_aligned_straddlesUpperBound; // @[PMP.scala 127:46]
  assign res_aligned_rangeAligned = ~_res_aligned_rangeAligned_T; // @[PMP.scala 127:24]
  assign _res_aligned_pow2Aligned_T_2 = ~_res_hit_lsbMask_T_1[2:0] & ~io_pmp_7_mask[2:0]; // @[PMP.scala 128:32]
  assign res_aligned_pow2Aligned = _res_aligned_pow2Aligned_T_2 == 3'h0; // @[PMP.scala 128:57]
  assign res_aligned = io_pmp_7_cfg_a[1] ? res_aligned_pow2Aligned : res_aligned_rangeAligned; // @[PMP.scala 129:8]
  assign _res_cur_cfg_r_T = io_pmp_7_cfg_r | res_ignore; // @[PMP.scala 183:40]
  assign res_cur_cfg_r = res_aligned & _res_cur_cfg_r_T; // @[PMP.scala 183:26]
  assign _res_cur_cfg_w_T = io_pmp_7_cfg_w | res_ignore; // @[PMP.scala 184:40]
  assign res_cur_cfg_w = res_aligned & _res_cur_cfg_w_T; // @[PMP.scala 184:26]
  assign _res_cur_cfg_x_T = io_pmp_7_cfg_x | res_ignore; // @[PMP.scala 185:40]
  assign res_cur_cfg_x = res_aligned & _res_cur_cfg_x_T; // @[PMP.scala 185:26]
  assign _res_T_44_cfg_x = res_hit ? res_cur_cfg_x : default_; // @[PMP.scala 186:8]
  assign _res_T_44_cfg_w = res_hit ? res_cur_cfg_w : default_; // @[PMP.scala 186:8]
  assign _res_T_44_cfg_r = res_hit ? res_cur_cfg_r : default_; // @[PMP.scala 186:8]
  assign res_hit_lsbMask_1 = io_pmp_6_mask | _GEN_0; // @[PMP.scala 70:26]
  assign _res_hit_msbMatch_T_19 = _res_hit_msbsEqual_T_6 & ~io_pmp_6_mask[31:3]; // @[PMP.scala 65:52]
  assign res_hit_msbMatch_1 = _res_hit_msbMatch_T_19 == 29'h0; // @[PMP.scala 65:58]
  assign _res_hit_lsbMatch_T_17 = io_addr[2:0] ^ _res_hit_lsbsLess_T_6; // @[PMP.scala 65:47]
  assign _res_hit_lsbMatch_T_19 = _res_hit_lsbMatch_T_17 & ~res_hit_lsbMask_1[2:0]; // @[PMP.scala 65:52]
  assign res_hit_lsbMatch_1 = _res_hit_lsbMatch_T_19 == 3'h0; // @[PMP.scala 65:58]
  assign _res_hit_T_15 = res_hit_msbMatch_1 & res_hit_lsbMatch_1; // @[PMP.scala 73:16]
  assign _res_hit_msbsLess_T_13 = {io_pmp_5_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _res_hit_msbsLess_T_15 = ~_res_hit_msbsLess_T_13 | 32'h3; // @[PMP.scala 62:48]
  assign _res_hit_msbsLess_T_17 = ~_res_hit_msbsLess_T_15[31:3]; // @[PMP.scala 82:52]
  assign res_hit_msbsLess_2 = io_addr[31:3] < _res_hit_msbsLess_T_17; // @[PMP.scala 82:39]
  assign _res_hit_msbsEqual_T_20 = io_addr[31:3] ^ _res_hit_msbsLess_T_17; // @[PMP.scala 83:41]
  assign res_hit_msbsEqual_2 = _res_hit_msbsEqual_T_20 == 29'h0; // @[PMP.scala 83:69]
  assign _res_hit_lsbsLess_T_20 = ~_res_hit_msbsLess_T_15[2:0]; // @[PMP.scala 84:64]
  assign res_hit_lsbsLess_2 = _res_hit_lsbsLess_T_1 < _res_hit_lsbsLess_T_20; // @[PMP.scala 84:53]
  assign _res_hit_T_21 = res_hit_msbsEqual_2 & res_hit_lsbsLess_2; // @[PMP.scala 85:30]
  assign _res_hit_T_22 = res_hit_msbsLess_2 | _res_hit_T_21; // @[PMP.scala 85:16]
  assign res_hit_lsbsLess_3 = io_addr[2:0] < _res_hit_lsbsLess_T_6; // @[PMP.scala 84:53]
  assign _res_hit_T_24 = res_hit_msbsEqual & res_hit_lsbsLess_3; // @[PMP.scala 85:30]
  assign _res_hit_T_25 = res_hit_msbsLess | _res_hit_T_24; // @[PMP.scala 85:16]
  assign _res_hit_T_26 = ~_res_hit_T_22 & _res_hit_T_25; // @[PMP.scala 96:48]
  assign _res_hit_T_27 = io_pmp_6_cfg_a[0] & _res_hit_T_26; // @[PMP.scala 134:61]
  assign res_hit_1 = io_pmp_6_cfg_a[1] ? _res_hit_T_15 : _res_hit_T_27; // @[PMP.scala 134:8]
  assign res_ignore_1 = default_ & ~io_pmp_6_cfg_l; // @[PMP.scala 165:26]
  assign _res_aligned_straddlesLowerBound_T_32 = _res_hit_lsbsLess_T_20 & ~io_addr[2:0]; // @[PMP.scala 125:123]
  assign _res_aligned_straddlesLowerBound_T_33 = _res_aligned_straddlesLowerBound_T_32 != 3'h0; // @[PMP.scala 125:145]
  assign res_aligned_straddlesLowerBound_1 = res_hit_msbsEqual_2 & _res_aligned_straddlesLowerBound_T_33; // @[PMP.scala 125:88]
  assign _res_aligned_straddlesUpperBound_T_32 = _res_hit_lsbsLess_T_6 & _res_hit_lsbsLess_T_1; // @[PMP.scala 126:113]
  assign _res_aligned_straddlesUpperBound_T_33 = _res_aligned_straddlesUpperBound_T_32 != 3'h0; // @[PMP.scala 126:146]
  assign res_aligned_straddlesUpperBound_1 = res_hit_msbsEqual & _res_aligned_straddlesUpperBound_T_33; // @[PMP.scala 126:83]
  assign _res_aligned_rangeAligned_T_1 = res_aligned_straddlesLowerBound_1 | res_aligned_straddlesUpperBound_1; // @[PMP.scala 127:46]
  assign res_aligned_rangeAligned_1 = ~_res_aligned_rangeAligned_T_1; // @[PMP.scala 127:24]
  assign _res_aligned_pow2Aligned_T_5 = ~_res_hit_lsbMask_T_1[2:0] & ~io_pmp_6_mask[2:0]; // @[PMP.scala 128:32]
  assign res_aligned_pow2Aligned_1 = _res_aligned_pow2Aligned_T_5 == 3'h0; // @[PMP.scala 128:57]
  assign res_aligned_1 = io_pmp_6_cfg_a[1] ? res_aligned_pow2Aligned_1 : res_aligned_rangeAligned_1; // @[PMP.scala 129:8]
  assign _res_cur_cfg_r_T_2 = io_pmp_6_cfg_r | res_ignore_1; // @[PMP.scala 183:40]
  assign res_cur_1_cfg_r = res_aligned_1 & _res_cur_cfg_r_T_2; // @[PMP.scala 183:26]
  assign _res_cur_cfg_w_T_2 = io_pmp_6_cfg_w | res_ignore_1; // @[PMP.scala 184:40]
  assign res_cur_1_cfg_w = res_aligned_1 & _res_cur_cfg_w_T_2; // @[PMP.scala 184:26]
  assign _res_cur_cfg_x_T_2 = io_pmp_6_cfg_x | res_ignore_1; // @[PMP.scala 185:40]
  assign res_cur_1_cfg_x = res_aligned_1 & _res_cur_cfg_x_T_2; // @[PMP.scala 185:26]
  assign _res_T_89_cfg_x = res_hit_1 ? res_cur_1_cfg_x : _res_T_44_cfg_x; // @[PMP.scala 186:8]
  assign _res_T_89_cfg_w = res_hit_1 ? res_cur_1_cfg_w : _res_T_44_cfg_w; // @[PMP.scala 186:8]
  assign _res_T_89_cfg_r = res_hit_1 ? res_cur_1_cfg_r : _res_T_44_cfg_r; // @[PMP.scala 186:8]
  assign res_hit_lsbMask_2 = io_pmp_5_mask | _GEN_0; // @[PMP.scala 70:26]
  assign _res_hit_msbMatch_T_29 = _res_hit_msbsEqual_T_20 & ~io_pmp_5_mask[31:3]; // @[PMP.scala 65:52]
  assign res_hit_msbMatch_2 = _res_hit_msbMatch_T_29 == 29'h0; // @[PMP.scala 65:58]
  assign _res_hit_lsbMatch_T_27 = io_addr[2:0] ^ _res_hit_lsbsLess_T_20; // @[PMP.scala 65:47]
  assign _res_hit_lsbMatch_T_29 = _res_hit_lsbMatch_T_27 & ~res_hit_lsbMask_2[2:0]; // @[PMP.scala 65:52]
  assign res_hit_lsbMatch_2 = _res_hit_lsbMatch_T_29 == 3'h0; // @[PMP.scala 65:58]
  assign _res_hit_T_29 = res_hit_msbMatch_2 & res_hit_lsbMatch_2; // @[PMP.scala 73:16]
  assign _res_hit_msbsLess_T_25 = {io_pmp_4_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _res_hit_msbsLess_T_27 = ~_res_hit_msbsLess_T_25 | 32'h3; // @[PMP.scala 62:48]
  assign _res_hit_msbsLess_T_29 = ~_res_hit_msbsLess_T_27[31:3]; // @[PMP.scala 82:52]
  assign res_hit_msbsLess_4 = io_addr[31:3] < _res_hit_msbsLess_T_29; // @[PMP.scala 82:39]
  assign _res_hit_msbsEqual_T_34 = io_addr[31:3] ^ _res_hit_msbsLess_T_29; // @[PMP.scala 83:41]
  assign res_hit_msbsEqual_4 = _res_hit_msbsEqual_T_34 == 29'h0; // @[PMP.scala 83:69]
  assign _res_hit_lsbsLess_T_34 = ~_res_hit_msbsLess_T_27[2:0]; // @[PMP.scala 84:64]
  assign res_hit_lsbsLess_4 = _res_hit_lsbsLess_T_1 < _res_hit_lsbsLess_T_34; // @[PMP.scala 84:53]
  assign _res_hit_T_35 = res_hit_msbsEqual_4 & res_hit_lsbsLess_4; // @[PMP.scala 85:30]
  assign _res_hit_T_36 = res_hit_msbsLess_4 | _res_hit_T_35; // @[PMP.scala 85:16]
  assign res_hit_lsbsLess_5 = io_addr[2:0] < _res_hit_lsbsLess_T_20; // @[PMP.scala 84:53]
  assign _res_hit_T_38 = res_hit_msbsEqual_2 & res_hit_lsbsLess_5; // @[PMP.scala 85:30]
  assign _res_hit_T_39 = res_hit_msbsLess_2 | _res_hit_T_38; // @[PMP.scala 85:16]
  assign _res_hit_T_40 = ~_res_hit_T_36 & _res_hit_T_39; // @[PMP.scala 96:48]
  assign _res_hit_T_41 = io_pmp_5_cfg_a[0] & _res_hit_T_40; // @[PMP.scala 134:61]
  assign res_hit_2 = io_pmp_5_cfg_a[1] ? _res_hit_T_29 : _res_hit_T_41; // @[PMP.scala 134:8]
  assign res_ignore_2 = default_ & ~io_pmp_5_cfg_l; // @[PMP.scala 165:26]
  assign _res_aligned_straddlesLowerBound_T_49 = _res_hit_lsbsLess_T_34 & ~io_addr[2:0]; // @[PMP.scala 125:123]
  assign _res_aligned_straddlesLowerBound_T_50 = _res_aligned_straddlesLowerBound_T_49 != 3'h0; // @[PMP.scala 125:145]
  assign res_aligned_straddlesLowerBound_2 = res_hit_msbsEqual_4 & _res_aligned_straddlesLowerBound_T_50; // @[PMP.scala 125:88]
  assign _res_aligned_straddlesUpperBound_T_49 = _res_hit_lsbsLess_T_20 & _res_hit_lsbsLess_T_1; // @[PMP.scala 126:113]
  assign _res_aligned_straddlesUpperBound_T_50 = _res_aligned_straddlesUpperBound_T_49 != 3'h0; // @[PMP.scala 126:146]
  assign res_aligned_straddlesUpperBound_2 = res_hit_msbsEqual_2 & _res_aligned_straddlesUpperBound_T_50; // @[PMP.scala 126:83]
  assign _res_aligned_rangeAligned_T_2 = res_aligned_straddlesLowerBound_2 | res_aligned_straddlesUpperBound_2; // @[PMP.scala 127:46]
  assign res_aligned_rangeAligned_2 = ~_res_aligned_rangeAligned_T_2; // @[PMP.scala 127:24]
  assign _res_aligned_pow2Aligned_T_8 = ~_res_hit_lsbMask_T_1[2:0] & ~io_pmp_5_mask[2:0]; // @[PMP.scala 128:32]
  assign res_aligned_pow2Aligned_2 = _res_aligned_pow2Aligned_T_8 == 3'h0; // @[PMP.scala 128:57]
  assign res_aligned_2 = io_pmp_5_cfg_a[1] ? res_aligned_pow2Aligned_2 : res_aligned_rangeAligned_2; // @[PMP.scala 129:8]
  assign _res_cur_cfg_r_T_4 = io_pmp_5_cfg_r | res_ignore_2; // @[PMP.scala 183:40]
  assign res_cur_2_cfg_r = res_aligned_2 & _res_cur_cfg_r_T_4; // @[PMP.scala 183:26]
  assign _res_cur_cfg_w_T_4 = io_pmp_5_cfg_w | res_ignore_2; // @[PMP.scala 184:40]
  assign res_cur_2_cfg_w = res_aligned_2 & _res_cur_cfg_w_T_4; // @[PMP.scala 184:26]
  assign _res_cur_cfg_x_T_4 = io_pmp_5_cfg_x | res_ignore_2; // @[PMP.scala 185:40]
  assign res_cur_2_cfg_x = res_aligned_2 & _res_cur_cfg_x_T_4; // @[PMP.scala 185:26]
  assign _res_T_134_cfg_x = res_hit_2 ? res_cur_2_cfg_x : _res_T_89_cfg_x; // @[PMP.scala 186:8]
  assign _res_T_134_cfg_w = res_hit_2 ? res_cur_2_cfg_w : _res_T_89_cfg_w; // @[PMP.scala 186:8]
  assign _res_T_134_cfg_r = res_hit_2 ? res_cur_2_cfg_r : _res_T_89_cfg_r; // @[PMP.scala 186:8]
  assign res_hit_lsbMask_3 = io_pmp_4_mask | _GEN_0; // @[PMP.scala 70:26]
  assign _res_hit_msbMatch_T_39 = _res_hit_msbsEqual_T_34 & ~io_pmp_4_mask[31:3]; // @[PMP.scala 65:52]
  assign res_hit_msbMatch_3 = _res_hit_msbMatch_T_39 == 29'h0; // @[PMP.scala 65:58]
  assign _res_hit_lsbMatch_T_37 = io_addr[2:0] ^ _res_hit_lsbsLess_T_34; // @[PMP.scala 65:47]
  assign _res_hit_lsbMatch_T_39 = _res_hit_lsbMatch_T_37 & ~res_hit_lsbMask_3[2:0]; // @[PMP.scala 65:52]
  assign res_hit_lsbMatch_3 = _res_hit_lsbMatch_T_39 == 3'h0; // @[PMP.scala 65:58]
  assign _res_hit_T_43 = res_hit_msbMatch_3 & res_hit_lsbMatch_3; // @[PMP.scala 73:16]
  assign _res_hit_msbsLess_T_37 = {io_pmp_3_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _res_hit_msbsLess_T_39 = ~_res_hit_msbsLess_T_37 | 32'h3; // @[PMP.scala 62:48]
  assign _res_hit_msbsLess_T_41 = ~_res_hit_msbsLess_T_39[31:3]; // @[PMP.scala 82:52]
  assign res_hit_msbsLess_6 = io_addr[31:3] < _res_hit_msbsLess_T_41; // @[PMP.scala 82:39]
  assign _res_hit_msbsEqual_T_48 = io_addr[31:3] ^ _res_hit_msbsLess_T_41; // @[PMP.scala 83:41]
  assign res_hit_msbsEqual_6 = _res_hit_msbsEqual_T_48 == 29'h0; // @[PMP.scala 83:69]
  assign _res_hit_lsbsLess_T_48 = ~_res_hit_msbsLess_T_39[2:0]; // @[PMP.scala 84:64]
  assign res_hit_lsbsLess_6 = _res_hit_lsbsLess_T_1 < _res_hit_lsbsLess_T_48; // @[PMP.scala 84:53]
  assign _res_hit_T_49 = res_hit_msbsEqual_6 & res_hit_lsbsLess_6; // @[PMP.scala 85:30]
  assign _res_hit_T_50 = res_hit_msbsLess_6 | _res_hit_T_49; // @[PMP.scala 85:16]
  assign res_hit_lsbsLess_7 = io_addr[2:0] < _res_hit_lsbsLess_T_34; // @[PMP.scala 84:53]
  assign _res_hit_T_52 = res_hit_msbsEqual_4 & res_hit_lsbsLess_7; // @[PMP.scala 85:30]
  assign _res_hit_T_53 = res_hit_msbsLess_4 | _res_hit_T_52; // @[PMP.scala 85:16]
  assign _res_hit_T_54 = ~_res_hit_T_50 & _res_hit_T_53; // @[PMP.scala 96:48]
  assign _res_hit_T_55 = io_pmp_4_cfg_a[0] & _res_hit_T_54; // @[PMP.scala 134:61]
  assign res_hit_3 = io_pmp_4_cfg_a[1] ? _res_hit_T_43 : _res_hit_T_55; // @[PMP.scala 134:8]
  assign res_ignore_3 = default_ & ~io_pmp_4_cfg_l; // @[PMP.scala 165:26]
  assign _res_aligned_straddlesLowerBound_T_66 = _res_hit_lsbsLess_T_48 & ~io_addr[2:0]; // @[PMP.scala 125:123]
  assign _res_aligned_straddlesLowerBound_T_67 = _res_aligned_straddlesLowerBound_T_66 != 3'h0; // @[PMP.scala 125:145]
  assign res_aligned_straddlesLowerBound_3 = res_hit_msbsEqual_6 & _res_aligned_straddlesLowerBound_T_67; // @[PMP.scala 125:88]
  assign _res_aligned_straddlesUpperBound_T_66 = _res_hit_lsbsLess_T_34 & _res_hit_lsbsLess_T_1; // @[PMP.scala 126:113]
  assign _res_aligned_straddlesUpperBound_T_67 = _res_aligned_straddlesUpperBound_T_66 != 3'h0; // @[PMP.scala 126:146]
  assign res_aligned_straddlesUpperBound_3 = res_hit_msbsEqual_4 & _res_aligned_straddlesUpperBound_T_67; // @[PMP.scala 126:83]
  assign _res_aligned_rangeAligned_T_3 = res_aligned_straddlesLowerBound_3 | res_aligned_straddlesUpperBound_3; // @[PMP.scala 127:46]
  assign res_aligned_rangeAligned_3 = ~_res_aligned_rangeAligned_T_3; // @[PMP.scala 127:24]
  assign _res_aligned_pow2Aligned_T_11 = ~_res_hit_lsbMask_T_1[2:0] & ~io_pmp_4_mask[2:0]; // @[PMP.scala 128:32]
  assign res_aligned_pow2Aligned_3 = _res_aligned_pow2Aligned_T_11 == 3'h0; // @[PMP.scala 128:57]
  assign res_aligned_3 = io_pmp_4_cfg_a[1] ? res_aligned_pow2Aligned_3 : res_aligned_rangeAligned_3; // @[PMP.scala 129:8]
  assign _res_cur_cfg_r_T_6 = io_pmp_4_cfg_r | res_ignore_3; // @[PMP.scala 183:40]
  assign res_cur_3_cfg_r = res_aligned_3 & _res_cur_cfg_r_T_6; // @[PMP.scala 183:26]
  assign _res_cur_cfg_w_T_6 = io_pmp_4_cfg_w | res_ignore_3; // @[PMP.scala 184:40]
  assign res_cur_3_cfg_w = res_aligned_3 & _res_cur_cfg_w_T_6; // @[PMP.scala 184:26]
  assign _res_cur_cfg_x_T_6 = io_pmp_4_cfg_x | res_ignore_3; // @[PMP.scala 185:40]
  assign res_cur_3_cfg_x = res_aligned_3 & _res_cur_cfg_x_T_6; // @[PMP.scala 185:26]
  assign _res_T_179_cfg_x = res_hit_3 ? res_cur_3_cfg_x : _res_T_134_cfg_x; // @[PMP.scala 186:8]
  assign _res_T_179_cfg_w = res_hit_3 ? res_cur_3_cfg_w : _res_T_134_cfg_w; // @[PMP.scala 186:8]
  assign _res_T_179_cfg_r = res_hit_3 ? res_cur_3_cfg_r : _res_T_134_cfg_r; // @[PMP.scala 186:8]
  assign res_hit_lsbMask_4 = io_pmp_3_mask | _GEN_0; // @[PMP.scala 70:26]
  assign _res_hit_msbMatch_T_49 = _res_hit_msbsEqual_T_48 & ~io_pmp_3_mask[31:3]; // @[PMP.scala 65:52]
  assign res_hit_msbMatch_4 = _res_hit_msbMatch_T_49 == 29'h0; // @[PMP.scala 65:58]
  assign _res_hit_lsbMatch_T_47 = io_addr[2:0] ^ _res_hit_lsbsLess_T_48; // @[PMP.scala 65:47]
  assign _res_hit_lsbMatch_T_49 = _res_hit_lsbMatch_T_47 & ~res_hit_lsbMask_4[2:0]; // @[PMP.scala 65:52]
  assign res_hit_lsbMatch_4 = _res_hit_lsbMatch_T_49 == 3'h0; // @[PMP.scala 65:58]
  assign _res_hit_T_57 = res_hit_msbMatch_4 & res_hit_lsbMatch_4; // @[PMP.scala 73:16]
  assign _res_hit_msbsLess_T_49 = {io_pmp_2_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _res_hit_msbsLess_T_51 = ~_res_hit_msbsLess_T_49 | 32'h3; // @[PMP.scala 62:48]
  assign _res_hit_msbsLess_T_53 = ~_res_hit_msbsLess_T_51[31:3]; // @[PMP.scala 82:52]
  assign res_hit_msbsLess_8 = io_addr[31:3] < _res_hit_msbsLess_T_53; // @[PMP.scala 82:39]
  assign _res_hit_msbsEqual_T_62 = io_addr[31:3] ^ _res_hit_msbsLess_T_53; // @[PMP.scala 83:41]
  assign res_hit_msbsEqual_8 = _res_hit_msbsEqual_T_62 == 29'h0; // @[PMP.scala 83:69]
  assign _res_hit_lsbsLess_T_62 = ~_res_hit_msbsLess_T_51[2:0]; // @[PMP.scala 84:64]
  assign res_hit_lsbsLess_8 = _res_hit_lsbsLess_T_1 < _res_hit_lsbsLess_T_62; // @[PMP.scala 84:53]
  assign _res_hit_T_63 = res_hit_msbsEqual_8 & res_hit_lsbsLess_8; // @[PMP.scala 85:30]
  assign _res_hit_T_64 = res_hit_msbsLess_8 | _res_hit_T_63; // @[PMP.scala 85:16]
  assign res_hit_lsbsLess_9 = io_addr[2:0] < _res_hit_lsbsLess_T_48; // @[PMP.scala 84:53]
  assign _res_hit_T_66 = res_hit_msbsEqual_6 & res_hit_lsbsLess_9; // @[PMP.scala 85:30]
  assign _res_hit_T_67 = res_hit_msbsLess_6 | _res_hit_T_66; // @[PMP.scala 85:16]
  assign _res_hit_T_68 = ~_res_hit_T_64 & _res_hit_T_67; // @[PMP.scala 96:48]
  assign _res_hit_T_69 = io_pmp_3_cfg_a[0] & _res_hit_T_68; // @[PMP.scala 134:61]
  assign res_hit_4 = io_pmp_3_cfg_a[1] ? _res_hit_T_57 : _res_hit_T_69; // @[PMP.scala 134:8]
  assign res_ignore_4 = default_ & ~io_pmp_3_cfg_l; // @[PMP.scala 165:26]
  assign _res_aligned_straddlesLowerBound_T_83 = _res_hit_lsbsLess_T_62 & ~io_addr[2:0]; // @[PMP.scala 125:123]
  assign _res_aligned_straddlesLowerBound_T_84 = _res_aligned_straddlesLowerBound_T_83 != 3'h0; // @[PMP.scala 125:145]
  assign res_aligned_straddlesLowerBound_4 = res_hit_msbsEqual_8 & _res_aligned_straddlesLowerBound_T_84; // @[PMP.scala 125:88]
  assign _res_aligned_straddlesUpperBound_T_83 = _res_hit_lsbsLess_T_48 & _res_hit_lsbsLess_T_1; // @[PMP.scala 126:113]
  assign _res_aligned_straddlesUpperBound_T_84 = _res_aligned_straddlesUpperBound_T_83 != 3'h0; // @[PMP.scala 126:146]
  assign res_aligned_straddlesUpperBound_4 = res_hit_msbsEqual_6 & _res_aligned_straddlesUpperBound_T_84; // @[PMP.scala 126:83]
  assign _res_aligned_rangeAligned_T_4 = res_aligned_straddlesLowerBound_4 | res_aligned_straddlesUpperBound_4; // @[PMP.scala 127:46]
  assign res_aligned_rangeAligned_4 = ~_res_aligned_rangeAligned_T_4; // @[PMP.scala 127:24]
  assign _res_aligned_pow2Aligned_T_14 = ~_res_hit_lsbMask_T_1[2:0] & ~io_pmp_3_mask[2:0]; // @[PMP.scala 128:32]
  assign res_aligned_pow2Aligned_4 = _res_aligned_pow2Aligned_T_14 == 3'h0; // @[PMP.scala 128:57]
  assign res_aligned_4 = io_pmp_3_cfg_a[1] ? res_aligned_pow2Aligned_4 : res_aligned_rangeAligned_4; // @[PMP.scala 129:8]
  assign _res_cur_cfg_r_T_8 = io_pmp_3_cfg_r | res_ignore_4; // @[PMP.scala 183:40]
  assign res_cur_4_cfg_r = res_aligned_4 & _res_cur_cfg_r_T_8; // @[PMP.scala 183:26]
  assign _res_cur_cfg_w_T_8 = io_pmp_3_cfg_w | res_ignore_4; // @[PMP.scala 184:40]
  assign res_cur_4_cfg_w = res_aligned_4 & _res_cur_cfg_w_T_8; // @[PMP.scala 184:26]
  assign _res_cur_cfg_x_T_8 = io_pmp_3_cfg_x | res_ignore_4; // @[PMP.scala 185:40]
  assign res_cur_4_cfg_x = res_aligned_4 & _res_cur_cfg_x_T_8; // @[PMP.scala 185:26]
  assign _res_T_224_cfg_x = res_hit_4 ? res_cur_4_cfg_x : _res_T_179_cfg_x; // @[PMP.scala 186:8]
  assign _res_T_224_cfg_w = res_hit_4 ? res_cur_4_cfg_w : _res_T_179_cfg_w; // @[PMP.scala 186:8]
  assign _res_T_224_cfg_r = res_hit_4 ? res_cur_4_cfg_r : _res_T_179_cfg_r; // @[PMP.scala 186:8]
  assign res_hit_lsbMask_5 = io_pmp_2_mask | _GEN_0; // @[PMP.scala 70:26]
  assign _res_hit_msbMatch_T_59 = _res_hit_msbsEqual_T_62 & ~io_pmp_2_mask[31:3]; // @[PMP.scala 65:52]
  assign res_hit_msbMatch_5 = _res_hit_msbMatch_T_59 == 29'h0; // @[PMP.scala 65:58]
  assign _res_hit_lsbMatch_T_57 = io_addr[2:0] ^ _res_hit_lsbsLess_T_62; // @[PMP.scala 65:47]
  assign _res_hit_lsbMatch_T_59 = _res_hit_lsbMatch_T_57 & ~res_hit_lsbMask_5[2:0]; // @[PMP.scala 65:52]
  assign res_hit_lsbMatch_5 = _res_hit_lsbMatch_T_59 == 3'h0; // @[PMP.scala 65:58]
  assign _res_hit_T_71 = res_hit_msbMatch_5 & res_hit_lsbMatch_5; // @[PMP.scala 73:16]
  assign _res_hit_msbsLess_T_61 = {io_pmp_1_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _res_hit_msbsLess_T_63 = ~_res_hit_msbsLess_T_61 | 32'h3; // @[PMP.scala 62:48]
  assign _res_hit_msbsLess_T_65 = ~_res_hit_msbsLess_T_63[31:3]; // @[PMP.scala 82:52]
  assign res_hit_msbsLess_10 = io_addr[31:3] < _res_hit_msbsLess_T_65; // @[PMP.scala 82:39]
  assign _res_hit_msbsEqual_T_76 = io_addr[31:3] ^ _res_hit_msbsLess_T_65; // @[PMP.scala 83:41]
  assign res_hit_msbsEqual_10 = _res_hit_msbsEqual_T_76 == 29'h0; // @[PMP.scala 83:69]
  assign _res_hit_lsbsLess_T_76 = ~_res_hit_msbsLess_T_63[2:0]; // @[PMP.scala 84:64]
  assign res_hit_lsbsLess_10 = _res_hit_lsbsLess_T_1 < _res_hit_lsbsLess_T_76; // @[PMP.scala 84:53]
  assign _res_hit_T_77 = res_hit_msbsEqual_10 & res_hit_lsbsLess_10; // @[PMP.scala 85:30]
  assign _res_hit_T_78 = res_hit_msbsLess_10 | _res_hit_T_77; // @[PMP.scala 85:16]
  assign res_hit_lsbsLess_11 = io_addr[2:0] < _res_hit_lsbsLess_T_62; // @[PMP.scala 84:53]
  assign _res_hit_T_80 = res_hit_msbsEqual_8 & res_hit_lsbsLess_11; // @[PMP.scala 85:30]
  assign _res_hit_T_81 = res_hit_msbsLess_8 | _res_hit_T_80; // @[PMP.scala 85:16]
  assign _res_hit_T_82 = ~_res_hit_T_78 & _res_hit_T_81; // @[PMP.scala 96:48]
  assign _res_hit_T_83 = io_pmp_2_cfg_a[0] & _res_hit_T_82; // @[PMP.scala 134:61]
  assign res_hit_5 = io_pmp_2_cfg_a[1] ? _res_hit_T_71 : _res_hit_T_83; // @[PMP.scala 134:8]
  assign res_ignore_5 = default_ & ~io_pmp_2_cfg_l; // @[PMP.scala 165:26]
  assign _res_aligned_straddlesLowerBound_T_100 = _res_hit_lsbsLess_T_76 & ~io_addr[2:0]; // @[PMP.scala 125:123]
  assign _res_aligned_straddlesLowerBound_T_101 = _res_aligned_straddlesLowerBound_T_100 != 3'h0; // @[PMP.scala 125:145]
  assign res_aligned_straddlesLowerBound_5 = res_hit_msbsEqual_10 & _res_aligned_straddlesLowerBound_T_101; // @[PMP.scala 125:88]
  assign _res_aligned_straddlesUpperBound_T_100 = _res_hit_lsbsLess_T_62 & _res_hit_lsbsLess_T_1; // @[PMP.scala 126:113]
  assign _res_aligned_straddlesUpperBound_T_101 = _res_aligned_straddlesUpperBound_T_100 != 3'h0; // @[PMP.scala 126:146]
  assign res_aligned_straddlesUpperBound_5 = res_hit_msbsEqual_8 & _res_aligned_straddlesUpperBound_T_101; // @[PMP.scala 126:83]
  assign _res_aligned_rangeAligned_T_5 = res_aligned_straddlesLowerBound_5 | res_aligned_straddlesUpperBound_5; // @[PMP.scala 127:46]
  assign res_aligned_rangeAligned_5 = ~_res_aligned_rangeAligned_T_5; // @[PMP.scala 127:24]
  assign _res_aligned_pow2Aligned_T_17 = ~_res_hit_lsbMask_T_1[2:0] & ~io_pmp_2_mask[2:0]; // @[PMP.scala 128:32]
  assign res_aligned_pow2Aligned_5 = _res_aligned_pow2Aligned_T_17 == 3'h0; // @[PMP.scala 128:57]
  assign res_aligned_5 = io_pmp_2_cfg_a[1] ? res_aligned_pow2Aligned_5 : res_aligned_rangeAligned_5; // @[PMP.scala 129:8]
  assign _res_cur_cfg_r_T_10 = io_pmp_2_cfg_r | res_ignore_5; // @[PMP.scala 183:40]
  assign res_cur_5_cfg_r = res_aligned_5 & _res_cur_cfg_r_T_10; // @[PMP.scala 183:26]
  assign _res_cur_cfg_w_T_10 = io_pmp_2_cfg_w | res_ignore_5; // @[PMP.scala 184:40]
  assign res_cur_5_cfg_w = res_aligned_5 & _res_cur_cfg_w_T_10; // @[PMP.scala 184:26]
  assign _res_cur_cfg_x_T_10 = io_pmp_2_cfg_x | res_ignore_5; // @[PMP.scala 185:40]
  assign res_cur_5_cfg_x = res_aligned_5 & _res_cur_cfg_x_T_10; // @[PMP.scala 185:26]
  assign _res_T_269_cfg_x = res_hit_5 ? res_cur_5_cfg_x : _res_T_224_cfg_x; // @[PMP.scala 186:8]
  assign _res_T_269_cfg_w = res_hit_5 ? res_cur_5_cfg_w : _res_T_224_cfg_w; // @[PMP.scala 186:8]
  assign _res_T_269_cfg_r = res_hit_5 ? res_cur_5_cfg_r : _res_T_224_cfg_r; // @[PMP.scala 186:8]
  assign res_hit_lsbMask_6 = io_pmp_1_mask | _GEN_0; // @[PMP.scala 70:26]
  assign _res_hit_msbMatch_T_69 = _res_hit_msbsEqual_T_76 & ~io_pmp_1_mask[31:3]; // @[PMP.scala 65:52]
  assign res_hit_msbMatch_6 = _res_hit_msbMatch_T_69 == 29'h0; // @[PMP.scala 65:58]
  assign _res_hit_lsbMatch_T_67 = io_addr[2:0] ^ _res_hit_lsbsLess_T_76; // @[PMP.scala 65:47]
  assign _res_hit_lsbMatch_T_69 = _res_hit_lsbMatch_T_67 & ~res_hit_lsbMask_6[2:0]; // @[PMP.scala 65:52]
  assign res_hit_lsbMatch_6 = _res_hit_lsbMatch_T_69 == 3'h0; // @[PMP.scala 65:58]
  assign _res_hit_T_85 = res_hit_msbMatch_6 & res_hit_lsbMatch_6; // @[PMP.scala 73:16]
  assign _res_hit_msbsLess_T_73 = {io_pmp_0_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _res_hit_msbsLess_T_75 = ~_res_hit_msbsLess_T_73 | 32'h3; // @[PMP.scala 62:48]
  assign _res_hit_msbsLess_T_77 = ~_res_hit_msbsLess_T_75[31:3]; // @[PMP.scala 82:52]
  assign res_hit_msbsLess_12 = io_addr[31:3] < _res_hit_msbsLess_T_77; // @[PMP.scala 82:39]
  assign _res_hit_msbsEqual_T_90 = io_addr[31:3] ^ _res_hit_msbsLess_T_77; // @[PMP.scala 83:41]
  assign res_hit_msbsEqual_12 = _res_hit_msbsEqual_T_90 == 29'h0; // @[PMP.scala 83:69]
  assign _res_hit_lsbsLess_T_90 = ~_res_hit_msbsLess_T_75[2:0]; // @[PMP.scala 84:64]
  assign res_hit_lsbsLess_12 = _res_hit_lsbsLess_T_1 < _res_hit_lsbsLess_T_90; // @[PMP.scala 84:53]
  assign _res_hit_T_91 = res_hit_msbsEqual_12 & res_hit_lsbsLess_12; // @[PMP.scala 85:30]
  assign _res_hit_T_92 = res_hit_msbsLess_12 | _res_hit_T_91; // @[PMP.scala 85:16]
  assign res_hit_lsbsLess_13 = io_addr[2:0] < _res_hit_lsbsLess_T_76; // @[PMP.scala 84:53]
  assign _res_hit_T_94 = res_hit_msbsEqual_10 & res_hit_lsbsLess_13; // @[PMP.scala 85:30]
  assign _res_hit_T_95 = res_hit_msbsLess_10 | _res_hit_T_94; // @[PMP.scala 85:16]
  assign _res_hit_T_96 = ~_res_hit_T_92 & _res_hit_T_95; // @[PMP.scala 96:48]
  assign _res_hit_T_97 = io_pmp_1_cfg_a[0] & _res_hit_T_96; // @[PMP.scala 134:61]
  assign res_hit_6 = io_pmp_1_cfg_a[1] ? _res_hit_T_85 : _res_hit_T_97; // @[PMP.scala 134:8]
  assign res_ignore_6 = default_ & ~io_pmp_1_cfg_l; // @[PMP.scala 165:26]
  assign _res_aligned_straddlesLowerBound_T_117 = _res_hit_lsbsLess_T_90 & ~io_addr[2:0]; // @[PMP.scala 125:123]
  assign _res_aligned_straddlesLowerBound_T_118 = _res_aligned_straddlesLowerBound_T_117 != 3'h0; // @[PMP.scala 125:145]
  assign res_aligned_straddlesLowerBound_6 = res_hit_msbsEqual_12 & _res_aligned_straddlesLowerBound_T_118; // @[PMP.scala 125:88]
  assign _res_aligned_straddlesUpperBound_T_117 = _res_hit_lsbsLess_T_76 & _res_hit_lsbsLess_T_1; // @[PMP.scala 126:113]
  assign _res_aligned_straddlesUpperBound_T_118 = _res_aligned_straddlesUpperBound_T_117 != 3'h0; // @[PMP.scala 126:146]
  assign res_aligned_straddlesUpperBound_6 = res_hit_msbsEqual_10 & _res_aligned_straddlesUpperBound_T_118; // @[PMP.scala 126:83]
  assign _res_aligned_rangeAligned_T_6 = res_aligned_straddlesLowerBound_6 | res_aligned_straddlesUpperBound_6; // @[PMP.scala 127:46]
  assign res_aligned_rangeAligned_6 = ~_res_aligned_rangeAligned_T_6; // @[PMP.scala 127:24]
  assign _res_aligned_pow2Aligned_T_20 = ~_res_hit_lsbMask_T_1[2:0] & ~io_pmp_1_mask[2:0]; // @[PMP.scala 128:32]
  assign res_aligned_pow2Aligned_6 = _res_aligned_pow2Aligned_T_20 == 3'h0; // @[PMP.scala 128:57]
  assign res_aligned_6 = io_pmp_1_cfg_a[1] ? res_aligned_pow2Aligned_6 : res_aligned_rangeAligned_6; // @[PMP.scala 129:8]
  assign _res_cur_cfg_r_T_12 = io_pmp_1_cfg_r | res_ignore_6; // @[PMP.scala 183:40]
  assign res_cur_6_cfg_r = res_aligned_6 & _res_cur_cfg_r_T_12; // @[PMP.scala 183:26]
  assign _res_cur_cfg_w_T_12 = io_pmp_1_cfg_w | res_ignore_6; // @[PMP.scala 184:40]
  assign res_cur_6_cfg_w = res_aligned_6 & _res_cur_cfg_w_T_12; // @[PMP.scala 184:26]
  assign _res_cur_cfg_x_T_12 = io_pmp_1_cfg_x | res_ignore_6; // @[PMP.scala 185:40]
  assign res_cur_6_cfg_x = res_aligned_6 & _res_cur_cfg_x_T_12; // @[PMP.scala 185:26]
  assign _res_T_314_cfg_x = res_hit_6 ? res_cur_6_cfg_x : _res_T_269_cfg_x; // @[PMP.scala 186:8]
  assign _res_T_314_cfg_w = res_hit_6 ? res_cur_6_cfg_w : _res_T_269_cfg_w; // @[PMP.scala 186:8]
  assign _res_T_314_cfg_r = res_hit_6 ? res_cur_6_cfg_r : _res_T_269_cfg_r; // @[PMP.scala 186:8]
  assign res_hit_lsbMask_7 = io_pmp_0_mask | _GEN_0; // @[PMP.scala 70:26]
  assign _res_hit_msbMatch_T_79 = _res_hit_msbsEqual_T_90 & ~io_pmp_0_mask[31:3]; // @[PMP.scala 65:52]
  assign res_hit_msbMatch_7 = _res_hit_msbMatch_T_79 == 29'h0; // @[PMP.scala 65:58]
  assign _res_hit_lsbMatch_T_77 = io_addr[2:0] ^ _res_hit_lsbsLess_T_90; // @[PMP.scala 65:47]
  assign _res_hit_lsbMatch_T_79 = _res_hit_lsbMatch_T_77 & ~res_hit_lsbMask_7[2:0]; // @[PMP.scala 65:52]
  assign res_hit_lsbMatch_7 = _res_hit_lsbMatch_T_79 == 3'h0; // @[PMP.scala 65:58]
  assign _res_hit_T_99 = res_hit_msbMatch_7 & res_hit_lsbMatch_7; // @[PMP.scala 73:16]
  assign res_hit_lsbsLess_15 = io_addr[2:0] < _res_hit_lsbsLess_T_90; // @[PMP.scala 84:53]
  assign _res_hit_T_108 = res_hit_msbsEqual_12 & res_hit_lsbsLess_15; // @[PMP.scala 85:30]
  assign _res_hit_T_109 = res_hit_msbsLess_12 | _res_hit_T_108; // @[PMP.scala 85:16]
  assign _res_hit_T_111 = io_pmp_0_cfg_a[0] & _res_hit_T_109; // @[PMP.scala 134:61]
  assign res_hit_7 = io_pmp_0_cfg_a[1] ? _res_hit_T_99 : _res_hit_T_111; // @[PMP.scala 134:8]
  assign res_ignore_7 = default_ & ~io_pmp_0_cfg_l; // @[PMP.scala 165:26]
  assign _res_aligned_straddlesUpperBound_T_134 = _res_hit_lsbsLess_T_90 & _res_hit_lsbsLess_T_1; // @[PMP.scala 126:113]
  assign _res_aligned_straddlesUpperBound_T_135 = _res_aligned_straddlesUpperBound_T_134 != 3'h0; // @[PMP.scala 126:146]
  assign res_aligned_straddlesUpperBound_7 = res_hit_msbsEqual_12 & _res_aligned_straddlesUpperBound_T_135; // @[PMP.scala 126:83]
  assign res_aligned_rangeAligned_7 = ~res_aligned_straddlesUpperBound_7; // @[PMP.scala 127:24]
  assign _res_aligned_pow2Aligned_T_23 = ~_res_hit_lsbMask_T_1[2:0] & ~io_pmp_0_mask[2:0]; // @[PMP.scala 128:32]
  assign res_aligned_pow2Aligned_7 = _res_aligned_pow2Aligned_T_23 == 3'h0; // @[PMP.scala 128:57]
  assign res_aligned_7 = io_pmp_0_cfg_a[1] ? res_aligned_pow2Aligned_7 : res_aligned_rangeAligned_7; // @[PMP.scala 129:8]
  assign _res_cur_cfg_r_T_14 = io_pmp_0_cfg_r | res_ignore_7; // @[PMP.scala 183:40]
  assign res_cur_7_cfg_r = res_aligned_7 & _res_cur_cfg_r_T_14; // @[PMP.scala 183:26]
  assign _res_cur_cfg_w_T_14 = io_pmp_0_cfg_w | res_ignore_7; // @[PMP.scala 184:40]
  assign res_cur_7_cfg_w = res_aligned_7 & _res_cur_cfg_w_T_14; // @[PMP.scala 184:26]
  assign _res_cur_cfg_x_T_14 = io_pmp_0_cfg_x | res_ignore_7; // @[PMP.scala 185:40]
  assign res_cur_7_cfg_x = res_aligned_7 & _res_cur_cfg_x_T_14; // @[PMP.scala 185:26]
  assign io_r = res_hit_7 ? res_cur_7_cfg_r : _res_T_314_cfg_r; // @[PMP.scala 189:8]
  assign io_w = res_hit_7 ? res_cur_7_cfg_w : _res_T_314_cfg_w; // @[PMP.scala 190:8]
  assign io_x = res_hit_7 ? res_cur_7_cfg_x : _res_T_314_cfg_x; // @[PMP.scala 191:8]
  assign PMPChecker_covSum = 30'h0;
  assign io_covSum = PMPChecker_covSum;
  assign metaAssert = 1'h0;
endmodule
module PMPChecker_2(
  input  [1:0]  io_prv,
  input         io_pmp_0_cfg_l,
  input  [1:0]  io_pmp_0_cfg_a,
  input         io_pmp_0_cfg_x,
  input         io_pmp_0_cfg_w,
  input         io_pmp_0_cfg_r,
  input  [29:0] io_pmp_0_addr,
  input  [31:0] io_pmp_0_mask,
  input         io_pmp_1_cfg_l,
  input  [1:0]  io_pmp_1_cfg_a,
  input         io_pmp_1_cfg_x,
  input         io_pmp_1_cfg_w,
  input         io_pmp_1_cfg_r,
  input  [29:0] io_pmp_1_addr,
  input  [31:0] io_pmp_1_mask,
  input         io_pmp_2_cfg_l,
  input  [1:0]  io_pmp_2_cfg_a,
  input         io_pmp_2_cfg_x,
  input         io_pmp_2_cfg_w,
  input         io_pmp_2_cfg_r,
  input  [29:0] io_pmp_2_addr,
  input  [31:0] io_pmp_2_mask,
  input         io_pmp_3_cfg_l,
  input  [1:0]  io_pmp_3_cfg_a,
  input         io_pmp_3_cfg_x,
  input         io_pmp_3_cfg_w,
  input         io_pmp_3_cfg_r,
  input  [29:0] io_pmp_3_addr,
  input  [31:0] io_pmp_3_mask,
  input         io_pmp_4_cfg_l,
  input  [1:0]  io_pmp_4_cfg_a,
  input         io_pmp_4_cfg_x,
  input         io_pmp_4_cfg_w,
  input         io_pmp_4_cfg_r,
  input  [29:0] io_pmp_4_addr,
  input  [31:0] io_pmp_4_mask,
  input         io_pmp_5_cfg_l,
  input  [1:0]  io_pmp_5_cfg_a,
  input         io_pmp_5_cfg_x,
  input         io_pmp_5_cfg_w,
  input         io_pmp_5_cfg_r,
  input  [29:0] io_pmp_5_addr,
  input  [31:0] io_pmp_5_mask,
  input         io_pmp_6_cfg_l,
  input  [1:0]  io_pmp_6_cfg_a,
  input         io_pmp_6_cfg_x,
  input         io_pmp_6_cfg_w,
  input         io_pmp_6_cfg_r,
  input  [29:0] io_pmp_6_addr,
  input  [31:0] io_pmp_6_mask,
  input         io_pmp_7_cfg_l,
  input  [1:0]  io_pmp_7_cfg_a,
  input         io_pmp_7_cfg_x,
  input         io_pmp_7_cfg_w,
  input         io_pmp_7_cfg_r,
  input  [29:0] io_pmp_7_addr,
  input  [31:0] io_pmp_7_mask,
  input  [31:0] io_addr,
  output        io_r,
  output        io_w,
  output        io_x,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  default_; // @[PMP.scala 157:56]
  wire [31:0] _res_hit_T_1; // @[PMP.scala 62:36]
  wire [31:0] _res_hit_T_3; // @[PMP.scala 62:48]
  wire [31:0] _res_hit_T_5; // @[PMP.scala 65:47]
  wire [31:0] _res_hit_T_7; // @[PMP.scala 65:52]
  wire  _res_hit_T_8; // @[PMP.scala 65:58]
  wire [31:0] _res_hit_T_14; // @[PMP.scala 62:36]
  wire [31:0] _res_hit_T_16; // @[PMP.scala 62:48]
  wire  _res_hit_T_18; // @[PMP.scala 79:9]
  wire  _res_hit_T_24; // @[PMP.scala 79:9]
  wire  _res_hit_T_25; // @[PMP.scala 96:48]
  wire  _res_hit_T_26; // @[PMP.scala 134:61]
  wire  res_hit; // @[PMP.scala 134:8]
  wire  res_ignore; // @[PMP.scala 165:26]
  wire  res_cur_cfg_r; // @[PMP.scala 183:40]
  wire  res_cur_cfg_w; // @[PMP.scala 184:40]
  wire  res_cur_cfg_x; // @[PMP.scala 185:40]
  wire  _res_T_44_cfg_x; // @[PMP.scala 186:8]
  wire  _res_T_44_cfg_w; // @[PMP.scala 186:8]
  wire  _res_T_44_cfg_r; // @[PMP.scala 186:8]
  wire [31:0] _res_hit_T_32; // @[PMP.scala 65:47]
  wire [31:0] _res_hit_T_34; // @[PMP.scala 65:52]
  wire  _res_hit_T_35; // @[PMP.scala 65:58]
  wire [31:0] _res_hit_T_41; // @[PMP.scala 62:36]
  wire [31:0] _res_hit_T_43; // @[PMP.scala 62:48]
  wire  _res_hit_T_45; // @[PMP.scala 79:9]
  wire  _res_hit_T_52; // @[PMP.scala 96:48]
  wire  _res_hit_T_53; // @[PMP.scala 134:61]
  wire  res_hit_1; // @[PMP.scala 134:8]
  wire  res_ignore_1; // @[PMP.scala 165:26]
  wire  res_cur_1_cfg_r; // @[PMP.scala 183:40]
  wire  res_cur_1_cfg_w; // @[PMP.scala 184:40]
  wire  res_cur_1_cfg_x; // @[PMP.scala 185:40]
  wire  _res_T_89_cfg_x; // @[PMP.scala 186:8]
  wire  _res_T_89_cfg_w; // @[PMP.scala 186:8]
  wire  _res_T_89_cfg_r; // @[PMP.scala 186:8]
  wire [31:0] _res_hit_T_59; // @[PMP.scala 65:47]
  wire [31:0] _res_hit_T_61; // @[PMP.scala 65:52]
  wire  _res_hit_T_62; // @[PMP.scala 65:58]
  wire [31:0] _res_hit_T_68; // @[PMP.scala 62:36]
  wire [31:0] _res_hit_T_70; // @[PMP.scala 62:48]
  wire  _res_hit_T_72; // @[PMP.scala 79:9]
  wire  _res_hit_T_79; // @[PMP.scala 96:48]
  wire  _res_hit_T_80; // @[PMP.scala 134:61]
  wire  res_hit_2; // @[PMP.scala 134:8]
  wire  res_ignore_2; // @[PMP.scala 165:26]
  wire  res_cur_2_cfg_r; // @[PMP.scala 183:40]
  wire  res_cur_2_cfg_w; // @[PMP.scala 184:40]
  wire  res_cur_2_cfg_x; // @[PMP.scala 185:40]
  wire  _res_T_134_cfg_x; // @[PMP.scala 186:8]
  wire  _res_T_134_cfg_w; // @[PMP.scala 186:8]
  wire  _res_T_134_cfg_r; // @[PMP.scala 186:8]
  wire [31:0] _res_hit_T_86; // @[PMP.scala 65:47]
  wire [31:0] _res_hit_T_88; // @[PMP.scala 65:52]
  wire  _res_hit_T_89; // @[PMP.scala 65:58]
  wire [31:0] _res_hit_T_95; // @[PMP.scala 62:36]
  wire [31:0] _res_hit_T_97; // @[PMP.scala 62:48]
  wire  _res_hit_T_99; // @[PMP.scala 79:9]
  wire  _res_hit_T_106; // @[PMP.scala 96:48]
  wire  _res_hit_T_107; // @[PMP.scala 134:61]
  wire  res_hit_3; // @[PMP.scala 134:8]
  wire  res_ignore_3; // @[PMP.scala 165:26]
  wire  res_cur_3_cfg_r; // @[PMP.scala 183:40]
  wire  res_cur_3_cfg_w; // @[PMP.scala 184:40]
  wire  res_cur_3_cfg_x; // @[PMP.scala 185:40]
  wire  _res_T_179_cfg_x; // @[PMP.scala 186:8]
  wire  _res_T_179_cfg_w; // @[PMP.scala 186:8]
  wire  _res_T_179_cfg_r; // @[PMP.scala 186:8]
  wire [31:0] _res_hit_T_113; // @[PMP.scala 65:47]
  wire [31:0] _res_hit_T_115; // @[PMP.scala 65:52]
  wire  _res_hit_T_116; // @[PMP.scala 65:58]
  wire [31:0] _res_hit_T_122; // @[PMP.scala 62:36]
  wire [31:0] _res_hit_T_124; // @[PMP.scala 62:48]
  wire  _res_hit_T_126; // @[PMP.scala 79:9]
  wire  _res_hit_T_133; // @[PMP.scala 96:48]
  wire  _res_hit_T_134; // @[PMP.scala 134:61]
  wire  res_hit_4; // @[PMP.scala 134:8]
  wire  res_ignore_4; // @[PMP.scala 165:26]
  wire  res_cur_4_cfg_r; // @[PMP.scala 183:40]
  wire  res_cur_4_cfg_w; // @[PMP.scala 184:40]
  wire  res_cur_4_cfg_x; // @[PMP.scala 185:40]
  wire  _res_T_224_cfg_x; // @[PMP.scala 186:8]
  wire  _res_T_224_cfg_w; // @[PMP.scala 186:8]
  wire  _res_T_224_cfg_r; // @[PMP.scala 186:8]
  wire [31:0] _res_hit_T_140; // @[PMP.scala 65:47]
  wire [31:0] _res_hit_T_142; // @[PMP.scala 65:52]
  wire  _res_hit_T_143; // @[PMP.scala 65:58]
  wire [31:0] _res_hit_T_149; // @[PMP.scala 62:36]
  wire [31:0] _res_hit_T_151; // @[PMP.scala 62:48]
  wire  _res_hit_T_153; // @[PMP.scala 79:9]
  wire  _res_hit_T_160; // @[PMP.scala 96:48]
  wire  _res_hit_T_161; // @[PMP.scala 134:61]
  wire  res_hit_5; // @[PMP.scala 134:8]
  wire  res_ignore_5; // @[PMP.scala 165:26]
  wire  res_cur_5_cfg_r; // @[PMP.scala 183:40]
  wire  res_cur_5_cfg_w; // @[PMP.scala 184:40]
  wire  res_cur_5_cfg_x; // @[PMP.scala 185:40]
  wire  _res_T_269_cfg_x; // @[PMP.scala 186:8]
  wire  _res_T_269_cfg_w; // @[PMP.scala 186:8]
  wire  _res_T_269_cfg_r; // @[PMP.scala 186:8]
  wire [31:0] _res_hit_T_167; // @[PMP.scala 65:47]
  wire [31:0] _res_hit_T_169; // @[PMP.scala 65:52]
  wire  _res_hit_T_170; // @[PMP.scala 65:58]
  wire [31:0] _res_hit_T_176; // @[PMP.scala 62:36]
  wire [31:0] _res_hit_T_178; // @[PMP.scala 62:48]
  wire  _res_hit_T_180; // @[PMP.scala 79:9]
  wire  _res_hit_T_187; // @[PMP.scala 96:48]
  wire  _res_hit_T_188; // @[PMP.scala 134:61]
  wire  res_hit_6; // @[PMP.scala 134:8]
  wire  res_ignore_6; // @[PMP.scala 165:26]
  wire  res_cur_6_cfg_r; // @[PMP.scala 183:40]
  wire  res_cur_6_cfg_w; // @[PMP.scala 184:40]
  wire  res_cur_6_cfg_x; // @[PMP.scala 185:40]
  wire  _res_T_314_cfg_x; // @[PMP.scala 186:8]
  wire  _res_T_314_cfg_w; // @[PMP.scala 186:8]
  wire  _res_T_314_cfg_r; // @[PMP.scala 186:8]
  wire [31:0] _res_hit_T_194; // @[PMP.scala 65:47]
  wire [31:0] _res_hit_T_196; // @[PMP.scala 65:52]
  wire  _res_hit_T_197; // @[PMP.scala 65:58]
  wire  _res_hit_T_215; // @[PMP.scala 134:61]
  wire  res_hit_7; // @[PMP.scala 134:8]
  wire  res_ignore_7; // @[PMP.scala 165:26]
  wire  res_cur_7_cfg_r; // @[PMP.scala 183:40]
  wire  res_cur_7_cfg_w; // @[PMP.scala 184:40]
  wire  res_cur_7_cfg_x; // @[PMP.scala 185:40]
  wire [29:0] PMPChecker_2_covSum;
  assign default_ = io_prv > 2'h1; // @[PMP.scala 157:56]
  assign _res_hit_T_1 = {io_pmp_7_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _res_hit_T_3 = ~_res_hit_T_1 | 32'h3; // @[PMP.scala 62:48]
  assign _res_hit_T_5 = io_addr ^ ~_res_hit_T_3; // @[PMP.scala 65:47]
  assign _res_hit_T_7 = _res_hit_T_5 & ~io_pmp_7_mask; // @[PMP.scala 65:52]
  assign _res_hit_T_8 = _res_hit_T_7 == 32'h0; // @[PMP.scala 65:58]
  assign _res_hit_T_14 = {io_pmp_6_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _res_hit_T_16 = ~_res_hit_T_14 | 32'h3; // @[PMP.scala 62:48]
  assign _res_hit_T_18 = io_addr < ~_res_hit_T_16; // @[PMP.scala 79:9]
  assign _res_hit_T_24 = io_addr < ~_res_hit_T_3; // @[PMP.scala 79:9]
  assign _res_hit_T_25 = ~_res_hit_T_18 & _res_hit_T_24; // @[PMP.scala 96:48]
  assign _res_hit_T_26 = io_pmp_7_cfg_a[0] & _res_hit_T_25; // @[PMP.scala 134:61]
  assign res_hit = io_pmp_7_cfg_a[1] ? _res_hit_T_8 : _res_hit_T_26; // @[PMP.scala 134:8]
  assign res_ignore = default_ & ~io_pmp_7_cfg_l; // @[PMP.scala 165:26]
  assign res_cur_cfg_r = io_pmp_7_cfg_r | res_ignore; // @[PMP.scala 183:40]
  assign res_cur_cfg_w = io_pmp_7_cfg_w | res_ignore; // @[PMP.scala 184:40]
  assign res_cur_cfg_x = io_pmp_7_cfg_x | res_ignore; // @[PMP.scala 185:40]
  assign _res_T_44_cfg_x = res_hit ? res_cur_cfg_x : default_; // @[PMP.scala 186:8]
  assign _res_T_44_cfg_w = res_hit ? res_cur_cfg_w : default_; // @[PMP.scala 186:8]
  assign _res_T_44_cfg_r = res_hit ? res_cur_cfg_r : default_; // @[PMP.scala 186:8]
  assign _res_hit_T_32 = io_addr ^ ~_res_hit_T_16; // @[PMP.scala 65:47]
  assign _res_hit_T_34 = _res_hit_T_32 & ~io_pmp_6_mask; // @[PMP.scala 65:52]
  assign _res_hit_T_35 = _res_hit_T_34 == 32'h0; // @[PMP.scala 65:58]
  assign _res_hit_T_41 = {io_pmp_5_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _res_hit_T_43 = ~_res_hit_T_41 | 32'h3; // @[PMP.scala 62:48]
  assign _res_hit_T_45 = io_addr < ~_res_hit_T_43; // @[PMP.scala 79:9]
  assign _res_hit_T_52 = ~_res_hit_T_45 & _res_hit_T_18; // @[PMP.scala 96:48]
  assign _res_hit_T_53 = io_pmp_6_cfg_a[0] & _res_hit_T_52; // @[PMP.scala 134:61]
  assign res_hit_1 = io_pmp_6_cfg_a[1] ? _res_hit_T_35 : _res_hit_T_53; // @[PMP.scala 134:8]
  assign res_ignore_1 = default_ & ~io_pmp_6_cfg_l; // @[PMP.scala 165:26]
  assign res_cur_1_cfg_r = io_pmp_6_cfg_r | res_ignore_1; // @[PMP.scala 183:40]
  assign res_cur_1_cfg_w = io_pmp_6_cfg_w | res_ignore_1; // @[PMP.scala 184:40]
  assign res_cur_1_cfg_x = io_pmp_6_cfg_x | res_ignore_1; // @[PMP.scala 185:40]
  assign _res_T_89_cfg_x = res_hit_1 ? res_cur_1_cfg_x : _res_T_44_cfg_x; // @[PMP.scala 186:8]
  assign _res_T_89_cfg_w = res_hit_1 ? res_cur_1_cfg_w : _res_T_44_cfg_w; // @[PMP.scala 186:8]
  assign _res_T_89_cfg_r = res_hit_1 ? res_cur_1_cfg_r : _res_T_44_cfg_r; // @[PMP.scala 186:8]
  assign _res_hit_T_59 = io_addr ^ ~_res_hit_T_43; // @[PMP.scala 65:47]
  assign _res_hit_T_61 = _res_hit_T_59 & ~io_pmp_5_mask; // @[PMP.scala 65:52]
  assign _res_hit_T_62 = _res_hit_T_61 == 32'h0; // @[PMP.scala 65:58]
  assign _res_hit_T_68 = {io_pmp_4_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _res_hit_T_70 = ~_res_hit_T_68 | 32'h3; // @[PMP.scala 62:48]
  assign _res_hit_T_72 = io_addr < ~_res_hit_T_70; // @[PMP.scala 79:9]
  assign _res_hit_T_79 = ~_res_hit_T_72 & _res_hit_T_45; // @[PMP.scala 96:48]
  assign _res_hit_T_80 = io_pmp_5_cfg_a[0] & _res_hit_T_79; // @[PMP.scala 134:61]
  assign res_hit_2 = io_pmp_5_cfg_a[1] ? _res_hit_T_62 : _res_hit_T_80; // @[PMP.scala 134:8]
  assign res_ignore_2 = default_ & ~io_pmp_5_cfg_l; // @[PMP.scala 165:26]
  assign res_cur_2_cfg_r = io_pmp_5_cfg_r | res_ignore_2; // @[PMP.scala 183:40]
  assign res_cur_2_cfg_w = io_pmp_5_cfg_w | res_ignore_2; // @[PMP.scala 184:40]
  assign res_cur_2_cfg_x = io_pmp_5_cfg_x | res_ignore_2; // @[PMP.scala 185:40]
  assign _res_T_134_cfg_x = res_hit_2 ? res_cur_2_cfg_x : _res_T_89_cfg_x; // @[PMP.scala 186:8]
  assign _res_T_134_cfg_w = res_hit_2 ? res_cur_2_cfg_w : _res_T_89_cfg_w; // @[PMP.scala 186:8]
  assign _res_T_134_cfg_r = res_hit_2 ? res_cur_2_cfg_r : _res_T_89_cfg_r; // @[PMP.scala 186:8]
  assign _res_hit_T_86 = io_addr ^ ~_res_hit_T_70; // @[PMP.scala 65:47]
  assign _res_hit_T_88 = _res_hit_T_86 & ~io_pmp_4_mask; // @[PMP.scala 65:52]
  assign _res_hit_T_89 = _res_hit_T_88 == 32'h0; // @[PMP.scala 65:58]
  assign _res_hit_T_95 = {io_pmp_3_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _res_hit_T_97 = ~_res_hit_T_95 | 32'h3; // @[PMP.scala 62:48]
  assign _res_hit_T_99 = io_addr < ~_res_hit_T_97; // @[PMP.scala 79:9]
  assign _res_hit_T_106 = ~_res_hit_T_99 & _res_hit_T_72; // @[PMP.scala 96:48]
  assign _res_hit_T_107 = io_pmp_4_cfg_a[0] & _res_hit_T_106; // @[PMP.scala 134:61]
  assign res_hit_3 = io_pmp_4_cfg_a[1] ? _res_hit_T_89 : _res_hit_T_107; // @[PMP.scala 134:8]
  assign res_ignore_3 = default_ & ~io_pmp_4_cfg_l; // @[PMP.scala 165:26]
  assign res_cur_3_cfg_r = io_pmp_4_cfg_r | res_ignore_3; // @[PMP.scala 183:40]
  assign res_cur_3_cfg_w = io_pmp_4_cfg_w | res_ignore_3; // @[PMP.scala 184:40]
  assign res_cur_3_cfg_x = io_pmp_4_cfg_x | res_ignore_3; // @[PMP.scala 185:40]
  assign _res_T_179_cfg_x = res_hit_3 ? res_cur_3_cfg_x : _res_T_134_cfg_x; // @[PMP.scala 186:8]
  assign _res_T_179_cfg_w = res_hit_3 ? res_cur_3_cfg_w : _res_T_134_cfg_w; // @[PMP.scala 186:8]
  assign _res_T_179_cfg_r = res_hit_3 ? res_cur_3_cfg_r : _res_T_134_cfg_r; // @[PMP.scala 186:8]
  assign _res_hit_T_113 = io_addr ^ ~_res_hit_T_97; // @[PMP.scala 65:47]
  assign _res_hit_T_115 = _res_hit_T_113 & ~io_pmp_3_mask; // @[PMP.scala 65:52]
  assign _res_hit_T_116 = _res_hit_T_115 == 32'h0; // @[PMP.scala 65:58]
  assign _res_hit_T_122 = {io_pmp_2_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _res_hit_T_124 = ~_res_hit_T_122 | 32'h3; // @[PMP.scala 62:48]
  assign _res_hit_T_126 = io_addr < ~_res_hit_T_124; // @[PMP.scala 79:9]
  assign _res_hit_T_133 = ~_res_hit_T_126 & _res_hit_T_99; // @[PMP.scala 96:48]
  assign _res_hit_T_134 = io_pmp_3_cfg_a[0] & _res_hit_T_133; // @[PMP.scala 134:61]
  assign res_hit_4 = io_pmp_3_cfg_a[1] ? _res_hit_T_116 : _res_hit_T_134; // @[PMP.scala 134:8]
  assign res_ignore_4 = default_ & ~io_pmp_3_cfg_l; // @[PMP.scala 165:26]
  assign res_cur_4_cfg_r = io_pmp_3_cfg_r | res_ignore_4; // @[PMP.scala 183:40]
  assign res_cur_4_cfg_w = io_pmp_3_cfg_w | res_ignore_4; // @[PMP.scala 184:40]
  assign res_cur_4_cfg_x = io_pmp_3_cfg_x | res_ignore_4; // @[PMP.scala 185:40]
  assign _res_T_224_cfg_x = res_hit_4 ? res_cur_4_cfg_x : _res_T_179_cfg_x; // @[PMP.scala 186:8]
  assign _res_T_224_cfg_w = res_hit_4 ? res_cur_4_cfg_w : _res_T_179_cfg_w; // @[PMP.scala 186:8]
  assign _res_T_224_cfg_r = res_hit_4 ? res_cur_4_cfg_r : _res_T_179_cfg_r; // @[PMP.scala 186:8]
  assign _res_hit_T_140 = io_addr ^ ~_res_hit_T_124; // @[PMP.scala 65:47]
  assign _res_hit_T_142 = _res_hit_T_140 & ~io_pmp_2_mask; // @[PMP.scala 65:52]
  assign _res_hit_T_143 = _res_hit_T_142 == 32'h0; // @[PMP.scala 65:58]
  assign _res_hit_T_149 = {io_pmp_1_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _res_hit_T_151 = ~_res_hit_T_149 | 32'h3; // @[PMP.scala 62:48]
  assign _res_hit_T_153 = io_addr < ~_res_hit_T_151; // @[PMP.scala 79:9]
  assign _res_hit_T_160 = ~_res_hit_T_153 & _res_hit_T_126; // @[PMP.scala 96:48]
  assign _res_hit_T_161 = io_pmp_2_cfg_a[0] & _res_hit_T_160; // @[PMP.scala 134:61]
  assign res_hit_5 = io_pmp_2_cfg_a[1] ? _res_hit_T_143 : _res_hit_T_161; // @[PMP.scala 134:8]
  assign res_ignore_5 = default_ & ~io_pmp_2_cfg_l; // @[PMP.scala 165:26]
  assign res_cur_5_cfg_r = io_pmp_2_cfg_r | res_ignore_5; // @[PMP.scala 183:40]
  assign res_cur_5_cfg_w = io_pmp_2_cfg_w | res_ignore_5; // @[PMP.scala 184:40]
  assign res_cur_5_cfg_x = io_pmp_2_cfg_x | res_ignore_5; // @[PMP.scala 185:40]
  assign _res_T_269_cfg_x = res_hit_5 ? res_cur_5_cfg_x : _res_T_224_cfg_x; // @[PMP.scala 186:8]
  assign _res_T_269_cfg_w = res_hit_5 ? res_cur_5_cfg_w : _res_T_224_cfg_w; // @[PMP.scala 186:8]
  assign _res_T_269_cfg_r = res_hit_5 ? res_cur_5_cfg_r : _res_T_224_cfg_r; // @[PMP.scala 186:8]
  assign _res_hit_T_167 = io_addr ^ ~_res_hit_T_151; // @[PMP.scala 65:47]
  assign _res_hit_T_169 = _res_hit_T_167 & ~io_pmp_1_mask; // @[PMP.scala 65:52]
  assign _res_hit_T_170 = _res_hit_T_169 == 32'h0; // @[PMP.scala 65:58]
  assign _res_hit_T_176 = {io_pmp_0_addr, 2'h0}; // @[PMP.scala 62:36]
  assign _res_hit_T_178 = ~_res_hit_T_176 | 32'h3; // @[PMP.scala 62:48]
  assign _res_hit_T_180 = io_addr < ~_res_hit_T_178; // @[PMP.scala 79:9]
  assign _res_hit_T_187 = ~_res_hit_T_180 & _res_hit_T_153; // @[PMP.scala 96:48]
  assign _res_hit_T_188 = io_pmp_1_cfg_a[0] & _res_hit_T_187; // @[PMP.scala 134:61]
  assign res_hit_6 = io_pmp_1_cfg_a[1] ? _res_hit_T_170 : _res_hit_T_188; // @[PMP.scala 134:8]
  assign res_ignore_6 = default_ & ~io_pmp_1_cfg_l; // @[PMP.scala 165:26]
  assign res_cur_6_cfg_r = io_pmp_1_cfg_r | res_ignore_6; // @[PMP.scala 183:40]
  assign res_cur_6_cfg_w = io_pmp_1_cfg_w | res_ignore_6; // @[PMP.scala 184:40]
  assign res_cur_6_cfg_x = io_pmp_1_cfg_x | res_ignore_6; // @[PMP.scala 185:40]
  assign _res_T_314_cfg_x = res_hit_6 ? res_cur_6_cfg_x : _res_T_269_cfg_x; // @[PMP.scala 186:8]
  assign _res_T_314_cfg_w = res_hit_6 ? res_cur_6_cfg_w : _res_T_269_cfg_w; // @[PMP.scala 186:8]
  assign _res_T_314_cfg_r = res_hit_6 ? res_cur_6_cfg_r : _res_T_269_cfg_r; // @[PMP.scala 186:8]
  assign _res_hit_T_194 = io_addr ^ ~_res_hit_T_178; // @[PMP.scala 65:47]
  assign _res_hit_T_196 = _res_hit_T_194 & ~io_pmp_0_mask; // @[PMP.scala 65:52]
  assign _res_hit_T_197 = _res_hit_T_196 == 32'h0; // @[PMP.scala 65:58]
  assign _res_hit_T_215 = io_pmp_0_cfg_a[0] & _res_hit_T_180; // @[PMP.scala 134:61]
  assign res_hit_7 = io_pmp_0_cfg_a[1] ? _res_hit_T_197 : _res_hit_T_215; // @[PMP.scala 134:8]
  assign res_ignore_7 = default_ & ~io_pmp_0_cfg_l; // @[PMP.scala 165:26]
  assign res_cur_7_cfg_r = io_pmp_0_cfg_r | res_ignore_7; // @[PMP.scala 183:40]
  assign res_cur_7_cfg_w = io_pmp_0_cfg_w | res_ignore_7; // @[PMP.scala 184:40]
  assign res_cur_7_cfg_x = io_pmp_0_cfg_x | res_ignore_7; // @[PMP.scala 185:40]
  assign io_r = res_hit_7 ? res_cur_7_cfg_r : _res_T_314_cfg_r; // @[PMP.scala 189:8]
  assign io_w = res_hit_7 ? res_cur_7_cfg_w : _res_T_314_cfg_w; // @[PMP.scala 190:8]
  assign io_x = res_hit_7 ? res_cur_7_cfg_x : _res_T_314_cfg_x; // @[PMP.scala 191:8]
  assign PMPChecker_2_covSum = 30'h0;
  assign io_covSum = PMPChecker_2_covSum;
  assign metaAssert = 1'h0;
endmodule
module MulAddRecFNPipe(
  input         clock,
  input         reset,
  input         io_validin,
  input  [1:0]  io_op,
  input  [32:0] io_a,
  input  [32:0] io_b,
  input  [32:0] io_c,
  input  [2:0]  io_roundingMode,
  output [32:0] io_out,
  output [4:0]  io_exceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  wire [1:0] mulAddRecFNToRaw_preMul_io_op; // @[FPU.scala 648:41]
  wire [32:0] mulAddRecFNToRaw_preMul_io_a; // @[FPU.scala 648:41]
  wire [32:0] mulAddRecFNToRaw_preMul_io_b; // @[FPU.scala 648:41]
  wire [32:0] mulAddRecFNToRaw_preMul_io_c; // @[FPU.scala 648:41]
  wire [23:0] mulAddRecFNToRaw_preMul_io_mulAddA; // @[FPU.scala 648:41]
  wire [23:0] mulAddRecFNToRaw_preMul_io_mulAddB; // @[FPU.scala 648:41]
  wire [47:0] mulAddRecFNToRaw_preMul_io_mulAddC; // @[FPU.scala 648:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny; // @[FPU.scala 648:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB; // @[FPU.scala 648:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfA; // @[FPU.scala 648:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA; // @[FPU.scala 648:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfB; // @[FPU.scala 648:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB; // @[FPU.scala 648:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_signProd; // @[FPU.scala 648:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC; // @[FPU.scala 648:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfC; // @[FPU.scala 648:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC; // @[FPU.scala 648:41]
  wire [9:0] mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum; // @[FPU.scala 648:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags; // @[FPU.scala 648:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant; // @[FPU.scala 648:41]
  wire [4:0] mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist; // @[FPU.scala 648:41]
  wire [25:0] mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC; // @[FPU.scala 648:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC; // @[FPU.scala 648:41]
  wire [29:0] mulAddRecFNToRaw_preMul_io_covSum; // @[FPU.scala 648:41]
  wire  mulAddRecFNToRaw_preMul_metaAssert; // @[FPU.scala 648:41]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny; // @[FPU.scala 649:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB; // @[FPU.scala 649:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA; // @[FPU.scala 649:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA; // @[FPU.scala 649:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB; // @[FPU.scala 649:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB; // @[FPU.scala 649:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_signProd; // @[FPU.scala 649:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC; // @[FPU.scala 649:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC; // @[FPU.scala 649:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC; // @[FPU.scala 649:42]
  wire [9:0] mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum; // @[FPU.scala 649:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags; // @[FPU.scala 649:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant; // @[FPU.scala 649:42]
  wire [4:0] mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist; // @[FPU.scala 649:42]
  wire [25:0] mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC; // @[FPU.scala 649:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC; // @[FPU.scala 649:42]
  wire [48:0] mulAddRecFNToRaw_postMul_io_mulAddResult; // @[FPU.scala 649:42]
  wire [2:0] mulAddRecFNToRaw_postMul_io_roundingMode; // @[FPU.scala 649:42]
  wire  mulAddRecFNToRaw_postMul_io_invalidExc; // @[FPU.scala 649:42]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isNaN; // @[FPU.scala 649:42]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isInf; // @[FPU.scala 649:42]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isZero; // @[FPU.scala 649:42]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_sign; // @[FPU.scala 649:42]
  wire [9:0] mulAddRecFNToRaw_postMul_io_rawOut_sExp; // @[FPU.scala 649:42]
  wire [26:0] mulAddRecFNToRaw_postMul_io_rawOut_sig; // @[FPU.scala 649:42]
  wire [29:0] mulAddRecFNToRaw_postMul_io_covSum; // @[FPU.scala 649:42]
  wire  mulAddRecFNToRaw_postMul_metaAssert; // @[FPU.scala 649:42]
  wire  roundRawFNToRecFN_io_invalidExc; // @[FPU.scala 676:35]
  wire  roundRawFNToRecFN_io_infiniteExc; // @[FPU.scala 676:35]
  wire  roundRawFNToRecFN_io_in_isNaN; // @[FPU.scala 676:35]
  wire  roundRawFNToRecFN_io_in_isInf; // @[FPU.scala 676:35]
  wire  roundRawFNToRecFN_io_in_isZero; // @[FPU.scala 676:35]
  wire  roundRawFNToRecFN_io_in_sign; // @[FPU.scala 676:35]
  wire [9:0] roundRawFNToRecFN_io_in_sExp; // @[FPU.scala 676:35]
  wire [26:0] roundRawFNToRecFN_io_in_sig; // @[FPU.scala 676:35]
  wire [2:0] roundRawFNToRecFN_io_roundingMode; // @[FPU.scala 676:35]
  wire  roundRawFNToRecFN_io_detectTininess; // @[FPU.scala 676:35]
  wire [32:0] roundRawFNToRecFN_io_out; // @[FPU.scala 676:35]
  wire [4:0] roundRawFNToRecFN_io_exceptionFlags; // @[FPU.scala 676:35]
  wire [29:0] roundRawFNToRecFN_io_covSum; // @[FPU.scala 676:35]
  wire  roundRawFNToRecFN_metaAssert; // @[FPU.scala 676:35]
  wire [47:0] _mulAddResult_T; // @[FPU.scala 657:45]
  wire [48:0] mulAddResult; // @[FPU.scala 658:50]
  reg  mulAddRecFNToRaw_postMul_io_fromPreMul_b_isSigNaNAny; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  reg  mulAddRecFNToRaw_postMul_io_fromPreMul_b_isNaNAOrB; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  reg  mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfA; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg  mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroA; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg  mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfB; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg  mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroB; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg  mulAddRecFNToRaw_postMul_io_fromPreMul_b_signProd; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg  mulAddRecFNToRaw_postMul_io_fromPreMul_b_isNaNC; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7;
  reg  mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfC; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8;
  reg  mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroC; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  reg [9:0] mulAddRecFNToRaw_postMul_io_fromPreMul_b_sExpSum; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10;
  reg  mulAddRecFNToRaw_postMul_io_fromPreMul_b_doSubMags; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11;
  reg  mulAddRecFNToRaw_postMul_io_fromPreMul_b_CIsDominant; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12;
  reg [4:0] mulAddRecFNToRaw_postMul_io_fromPreMul_b_CDom_CAlignDist; // @[Reg.scala 15:16]
  reg [31:0] _RAND_13;
  reg [25:0] mulAddRecFNToRaw_postMul_io_fromPreMul_b_highAlignedSigC; // @[Reg.scala 15:16]
  reg [31:0] _RAND_14;
  reg  mulAddRecFNToRaw_postMul_io_fromPreMul_b_bit0AlignedSigC; // @[Reg.scala 15:16]
  reg [31:0] _RAND_15;
  reg [48:0] mulAddRecFNToRaw_postMul_io_mulAddResult_b; // @[Reg.scala 15:16]
  reg [63:0] _RAND_16;
  reg [2:0] mulAddRecFNToRaw_postMul_io_roundingMode_b; // @[Reg.scala 15:16]
  reg [31:0] _RAND_17;
  reg [2:0] roundingMode_stage0_b; // @[Reg.scala 15:16]
  reg [31:0] _RAND_18;
  reg  detectTininess_stage0_b; // @[Reg.scala 15:16]
  reg [31:0] _RAND_19;
  reg  valid_stage0_v; // @[Valid.scala 117:22]
  reg [31:0] _RAND_20;
  reg  roundRawFNToRecFN_io_invalidExc_b; // @[Reg.scala 15:16]
  reg [31:0] _RAND_21;
  reg  roundRawFNToRecFN_io_in_b_isNaN; // @[Reg.scala 15:16]
  reg [31:0] _RAND_22;
  reg  roundRawFNToRecFN_io_in_b_isInf; // @[Reg.scala 15:16]
  reg [31:0] _RAND_23;
  reg  roundRawFNToRecFN_io_in_b_isZero; // @[Reg.scala 15:16]
  reg [31:0] _RAND_24;
  reg  roundRawFNToRecFN_io_in_b_sign; // @[Reg.scala 15:16]
  reg [31:0] _RAND_25;
  reg [9:0] roundRawFNToRecFN_io_in_b_sExp; // @[Reg.scala 15:16]
  reg [31:0] _RAND_26;
  reg [26:0] roundRawFNToRecFN_io_in_b_sig; // @[Reg.scala 15:16]
  reg [31:0] _RAND_27;
  reg [2:0] roundRawFNToRecFN_io_roundingMode_b; // @[Reg.scala 15:16]
  reg [31:0] _RAND_28;
  reg  roundRawFNToRecFN_io_detectTininess_b; // @[Reg.scala 15:16]
  reg [31:0] _RAND_29;
  reg  MulAddRecFNPipe_state; // @[Register tracking MulAddRecFNPipe state]
  reg [31:0] _RAND_30;
  reg  MulAddRecFNPipe_cov [0:1]; // @[Coverage map for MulAddRecFNPipe]
  reg [31:0] _RAND_31;
  wire  MulAddRecFNPipe_cov_read_data; // @[Coverage map for MulAddRecFNPipe]
  wire  MulAddRecFNPipe_cov_read_addr; // @[Coverage map for MulAddRecFNPipe]
  wire  MulAddRecFNPipe_cov_write_data; // @[Coverage map for MulAddRecFNPipe]
  wire  MulAddRecFNPipe_cov_write_addr; // @[Coverage map for MulAddRecFNPipe]
  wire  MulAddRecFNPipe_cov_write_mask; // @[Coverage map for MulAddRecFNPipe]
  wire  MulAddRecFNPipe_cov_write_en; // @[Coverage map for MulAddRecFNPipe]
  reg [29:0] MulAddRecFNPipe_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_32;
  wire  valid_stage0_v_shl;
  wire  valid_stage0_v_pad;
  wire [29:0] mulAddRecFNToRaw_preMul_sum;
  wire [29:0] mulAddRecFNToRaw_postMul_sum;
  wire [29:0] roundRawFNToRecFN_sum;
  wire  mulAddRecFNToRaw_preMul_metaAssert_wire;
  wire  mulAddRecFNToRaw_postMul_metaAssert_wire;
  wire  roundRawFNToRecFN_metaAssert_wire;
  wire  MulAddRecFNPipe_or2;
  wire  MulAddRecFNPipe_or0;
  reg  MulAddRecFNPipe_metaAssert;
  reg [31:0] _RAND_33;
  MulAddRecFNToRaw_preMul mulAddRecFNToRaw_preMul ( // @[FPU.scala 648:41]
    .io_op(mulAddRecFNToRaw_preMul_io_op),
    .io_a(mulAddRecFNToRaw_preMul_io_a),
    .io_b(mulAddRecFNToRaw_preMul_io_b),
    .io_c(mulAddRecFNToRaw_preMul_io_c),
    .io_mulAddA(mulAddRecFNToRaw_preMul_io_mulAddA),
    .io_mulAddB(mulAddRecFNToRaw_preMul_io_mulAddB),
    .io_mulAddC(mulAddRecFNToRaw_preMul_io_mulAddC),
    .io_toPostMul_isSigNaNAny(mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny),
    .io_toPostMul_isNaNAOrB(mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB),
    .io_toPostMul_isInfA(mulAddRecFNToRaw_preMul_io_toPostMul_isInfA),
    .io_toPostMul_isZeroA(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA),
    .io_toPostMul_isInfB(mulAddRecFNToRaw_preMul_io_toPostMul_isInfB),
    .io_toPostMul_isZeroB(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB),
    .io_toPostMul_signProd(mulAddRecFNToRaw_preMul_io_toPostMul_signProd),
    .io_toPostMul_isNaNC(mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC),
    .io_toPostMul_isInfC(mulAddRecFNToRaw_preMul_io_toPostMul_isInfC),
    .io_toPostMul_isZeroC(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC),
    .io_toPostMul_sExpSum(mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum),
    .io_toPostMul_doSubMags(mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags),
    .io_toPostMul_CIsDominant(mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant),
    .io_toPostMul_CDom_CAlignDist(mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist),
    .io_toPostMul_highAlignedSigC(mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC),
    .io_toPostMul_bit0AlignedSigC(mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC),
    .io_covSum(mulAddRecFNToRaw_preMul_io_covSum),
    .metaAssert(mulAddRecFNToRaw_preMul_metaAssert)
  );
  MulAddRecFNToRaw_postMul mulAddRecFNToRaw_postMul ( // @[FPU.scala 649:42]
    .io_fromPreMul_isSigNaNAny(mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny),
    .io_fromPreMul_isNaNAOrB(mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB),
    .io_fromPreMul_isInfA(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA),
    .io_fromPreMul_isZeroA(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA),
    .io_fromPreMul_isInfB(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB),
    .io_fromPreMul_isZeroB(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB),
    .io_fromPreMul_signProd(mulAddRecFNToRaw_postMul_io_fromPreMul_signProd),
    .io_fromPreMul_isNaNC(mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC),
    .io_fromPreMul_isInfC(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC),
    .io_fromPreMul_isZeroC(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC),
    .io_fromPreMul_sExpSum(mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum),
    .io_fromPreMul_doSubMags(mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags),
    .io_fromPreMul_CIsDominant(mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant),
    .io_fromPreMul_CDom_CAlignDist(mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist),
    .io_fromPreMul_highAlignedSigC(mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC),
    .io_fromPreMul_bit0AlignedSigC(mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC),
    .io_mulAddResult(mulAddRecFNToRaw_postMul_io_mulAddResult),
    .io_roundingMode(mulAddRecFNToRaw_postMul_io_roundingMode),
    .io_invalidExc(mulAddRecFNToRaw_postMul_io_invalidExc),
    .io_rawOut_isNaN(mulAddRecFNToRaw_postMul_io_rawOut_isNaN),
    .io_rawOut_isInf(mulAddRecFNToRaw_postMul_io_rawOut_isInf),
    .io_rawOut_isZero(mulAddRecFNToRaw_postMul_io_rawOut_isZero),
    .io_rawOut_sign(mulAddRecFNToRaw_postMul_io_rawOut_sign),
    .io_rawOut_sExp(mulAddRecFNToRaw_postMul_io_rawOut_sExp),
    .io_rawOut_sig(mulAddRecFNToRaw_postMul_io_rawOut_sig),
    .io_covSum(mulAddRecFNToRaw_postMul_io_covSum),
    .metaAssert(mulAddRecFNToRaw_postMul_metaAssert)
  );
  RoundRawFNToRecFN_2 roundRawFNToRecFN ( // @[FPU.scala 676:35]
    .io_invalidExc(roundRawFNToRecFN_io_invalidExc),
    .io_infiniteExc(roundRawFNToRecFN_io_infiniteExc),
    .io_in_isNaN(roundRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundRawFNToRecFN_io_in_sig),
    .io_roundingMode(roundRawFNToRecFN_io_roundingMode),
    .io_detectTininess(roundRawFNToRecFN_io_detectTininess),
    .io_out(roundRawFNToRecFN_io_out),
    .io_exceptionFlags(roundRawFNToRecFN_io_exceptionFlags),
    .io_covSum(roundRawFNToRecFN_io_covSum),
    .metaAssert(roundRawFNToRecFN_metaAssert)
  );
  assign _mulAddResult_T = mulAddRecFNToRaw_preMul_io_mulAddA * mulAddRecFNToRaw_preMul_io_mulAddB; // @[FPU.scala 657:45]
  assign mulAddResult = _mulAddResult_T + mulAddRecFNToRaw_preMul_io_mulAddC; // @[FPU.scala 658:50]
  assign io_out = roundRawFNToRecFN_io_out; // @[FPU.scala 687:23]
  assign io_exceptionFlags = roundRawFNToRecFN_io_exceptionFlags; // @[FPU.scala 688:23]
  assign mulAddRecFNToRaw_preMul_io_op = io_op; // @[FPU.scala 651:35]
  assign mulAddRecFNToRaw_preMul_io_a = io_a; // @[FPU.scala 652:35]
  assign mulAddRecFNToRaw_preMul_io_b = io_b; // @[FPU.scala 653:35]
  assign mulAddRecFNToRaw_preMul_io_c = io_c; // @[FPU.scala 654:35]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny = mulAddRecFNToRaw_postMul_io_fromPreMul_b_isSigNaNAny; // @[FPU.scala 666:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB = mulAddRecFNToRaw_postMul_io_fromPreMul_b_isNaNAOrB; // @[FPU.scala 666:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA = mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfA; // @[FPU.scala 666:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA = mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroA; // @[FPU.scala 666:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB = mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfB; // @[FPU.scala 666:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB = mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroB; // @[FPU.scala 666:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_signProd = mulAddRecFNToRaw_postMul_io_fromPreMul_b_signProd; // @[FPU.scala 666:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC = mulAddRecFNToRaw_postMul_io_fromPreMul_b_isNaNC; // @[FPU.scala 666:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC = mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfC; // @[FPU.scala 666:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC = mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroC; // @[FPU.scala 666:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum = mulAddRecFNToRaw_postMul_io_fromPreMul_b_sExpSum; // @[FPU.scala 666:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags = mulAddRecFNToRaw_postMul_io_fromPreMul_b_doSubMags; // @[FPU.scala 666:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant = mulAddRecFNToRaw_postMul_io_fromPreMul_b_CIsDominant; // @[FPU.scala 666:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist = mulAddRecFNToRaw_postMul_io_fromPreMul_b_CDom_CAlignDist; // @[FPU.scala 666:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC = mulAddRecFNToRaw_postMul_io_fromPreMul_b_highAlignedSigC; // @[FPU.scala 666:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC = mulAddRecFNToRaw_postMul_io_fromPreMul_b_bit0AlignedSigC; // @[FPU.scala 666:46]
  assign mulAddRecFNToRaw_postMul_io_mulAddResult = mulAddRecFNToRaw_postMul_io_mulAddResult_b; // @[FPU.scala 667:46]
  assign mulAddRecFNToRaw_postMul_io_roundingMode = mulAddRecFNToRaw_postMul_io_roundingMode_b; // @[FPU.scala 668:46]
  assign roundRawFNToRecFN_io_invalidExc = roundRawFNToRecFN_io_invalidExc_b; // @[FPU.scala 679:45]
  assign roundRawFNToRecFN_io_infiniteExc = 1'h0; // @[FPU.scala 685:38]
  assign roundRawFNToRecFN_io_in_isNaN = roundRawFNToRecFN_io_in_b_isNaN; // @[FPU.scala 680:45]
  assign roundRawFNToRecFN_io_in_isInf = roundRawFNToRecFN_io_in_b_isInf; // @[FPU.scala 680:45]
  assign roundRawFNToRecFN_io_in_isZero = roundRawFNToRecFN_io_in_b_isZero; // @[FPU.scala 680:45]
  assign roundRawFNToRecFN_io_in_sign = roundRawFNToRecFN_io_in_b_sign; // @[FPU.scala 680:45]
  assign roundRawFNToRecFN_io_in_sExp = roundRawFNToRecFN_io_in_b_sExp; // @[FPU.scala 680:45]
  assign roundRawFNToRecFN_io_in_sig = roundRawFNToRecFN_io_in_b_sig; // @[FPU.scala 680:45]
  assign roundRawFNToRecFN_io_roundingMode = roundRawFNToRecFN_io_roundingMode_b; // @[FPU.scala 681:45]
  assign roundRawFNToRecFN_io_detectTininess = roundRawFNToRecFN_io_detectTininess_b; // @[FPU.scala 682:45]
  assign MulAddRecFNPipe_cov_read_addr = MulAddRecFNPipe_state;
  assign MulAddRecFNPipe_cov_read_data = MulAddRecFNPipe_cov[MulAddRecFNPipe_cov_read_addr]; // @[Coverage map for MulAddRecFNPipe]
  assign MulAddRecFNPipe_cov_write_data = 1'h1;
  assign MulAddRecFNPipe_cov_write_addr = MulAddRecFNPipe_state;
  assign MulAddRecFNPipe_cov_write_mask = 1'h1;
  assign MulAddRecFNPipe_cov_write_en = 1'h1;
  assign valid_stage0_v_shl = valid_stage0_v;
  assign valid_stage0_v_pad = valid_stage0_v_shl;
  assign mulAddRecFNToRaw_preMul_sum = MulAddRecFNPipe_covSum + mulAddRecFNToRaw_preMul_io_covSum;
  assign mulAddRecFNToRaw_postMul_sum = mulAddRecFNToRaw_preMul_sum + mulAddRecFNToRaw_postMul_io_covSum;
  assign roundRawFNToRecFN_sum = mulAddRecFNToRaw_postMul_sum + roundRawFNToRecFN_io_covSum;
  assign io_covSum = roundRawFNToRecFN_sum;
  assign mulAddRecFNToRaw_preMul_metaAssert_wire = mulAddRecFNToRaw_preMul_metaAssert;
  assign mulAddRecFNToRaw_postMul_metaAssert_wire = mulAddRecFNToRaw_postMul_metaAssert;
  assign roundRawFNToRecFN_metaAssert_wire = roundRawFNToRecFN_metaAssert;
  assign MulAddRecFNPipe_or2 = mulAddRecFNToRaw_postMul_metaAssert_wire | roundRawFNToRecFN_metaAssert_wire;
  assign MulAddRecFNPipe_or0 = mulAddRecFNToRaw_preMul_metaAssert_wire | MulAddRecFNPipe_or2;
  assign metaAssert = MulAddRecFNPipe_metaAssert;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mulAddRecFNToRaw_postMul_io_fromPreMul_b_isSigNaNAny = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mulAddRecFNToRaw_postMul_io_fromPreMul_b_isNaNAOrB = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfA = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroA = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfB = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroB = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  mulAddRecFNToRaw_postMul_io_fromPreMul_b_signProd = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  mulAddRecFNToRaw_postMul_io_fromPreMul_b_isNaNC = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfC = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroC = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  mulAddRecFNToRaw_postMul_io_fromPreMul_b_sExpSum = _RAND_10[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  mulAddRecFNToRaw_postMul_io_fromPreMul_b_doSubMags = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  mulAddRecFNToRaw_postMul_io_fromPreMul_b_CIsDominant = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  mulAddRecFNToRaw_postMul_io_fromPreMul_b_CDom_CAlignDist = _RAND_13[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  mulAddRecFNToRaw_postMul_io_fromPreMul_b_highAlignedSigC = _RAND_14[25:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  mulAddRecFNToRaw_postMul_io_fromPreMul_b_bit0AlignedSigC = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {2{`RANDOM}};
  mulAddRecFNToRaw_postMul_io_mulAddResult_b = _RAND_16[48:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  mulAddRecFNToRaw_postMul_io_roundingMode_b = _RAND_17[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  roundingMode_stage0_b = _RAND_18[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  detectTininess_stage0_b = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  valid_stage0_v = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  roundRawFNToRecFN_io_invalidExc_b = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  roundRawFNToRecFN_io_in_b_isNaN = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  roundRawFNToRecFN_io_in_b_isInf = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  roundRawFNToRecFN_io_in_b_isZero = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  roundRawFNToRecFN_io_in_b_sign = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  roundRawFNToRecFN_io_in_b_sExp = _RAND_26[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  roundRawFNToRecFN_io_in_b_sig = _RAND_27[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  roundRawFNToRecFN_io_roundingMode_b = _RAND_28[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  roundRawFNToRecFN_io_detectTininess_b = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  MulAddRecFNPipe_state = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    MulAddRecFNPipe_cov[initvar] = _RAND_31[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  MulAddRecFNPipe_covSum = _RAND_32[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  MulAddRecFNPipe_metaAssert = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_isSigNaNAny <= 1'h0;
    end else if (io_validin) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_isSigNaNAny <= mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny;
    end
    if (metaReset) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_isNaNAOrB <= 1'h0;
    end else if (io_validin) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_isNaNAOrB <= mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB;
    end
    if (metaReset) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfA <= 1'h0;
    end else if (io_validin) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfA <= mulAddRecFNToRaw_preMul_io_toPostMul_isInfA;
    end
    if (metaReset) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroA <= 1'h0;
    end else if (io_validin) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroA <= mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA;
    end
    if (metaReset) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfB <= 1'h0;
    end else if (io_validin) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfB <= mulAddRecFNToRaw_preMul_io_toPostMul_isInfB;
    end
    if (metaReset) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroB <= 1'h0;
    end else if (io_validin) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroB <= mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB;
    end
    if (metaReset) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_signProd <= 1'h0;
    end else if (io_validin) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_signProd <= mulAddRecFNToRaw_preMul_io_toPostMul_signProd;
    end
    if (metaReset) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_isNaNC <= 1'h0;
    end else if (io_validin) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_isNaNC <= mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC;
    end
    if (metaReset) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfC <= 1'h0;
    end else if (io_validin) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfC <= mulAddRecFNToRaw_preMul_io_toPostMul_isInfC;
    end
    if (metaReset) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroC <= 1'h0;
    end else if (io_validin) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroC <= mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC;
    end
    if (metaReset) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_sExpSum <= 10'h0;
    end else if (io_validin) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_sExpSum <= mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum;
    end
    if (metaReset) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_doSubMags <= 1'h0;
    end else if (io_validin) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_doSubMags <= mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags;
    end
    if (metaReset) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_CIsDominant <= 1'h0;
    end else if (io_validin) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_CIsDominant <= mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant;
    end
    if (metaReset) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_CDom_CAlignDist <= 5'h0;
    end else if (io_validin) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_CDom_CAlignDist <= mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist;
    end
    if (metaReset) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_highAlignedSigC <= 26'h0;
    end else if (io_validin) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_highAlignedSigC <= mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC;
    end
    if (metaReset) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_bit0AlignedSigC <= 1'h0;
    end else if (io_validin) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_bit0AlignedSigC <= mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC;
    end
    if (metaReset) begin
      mulAddRecFNToRaw_postMul_io_mulAddResult_b <= 49'h0;
    end else if (io_validin) begin
      mulAddRecFNToRaw_postMul_io_mulAddResult_b <= mulAddResult;
    end
    if (metaReset) begin
      mulAddRecFNToRaw_postMul_io_roundingMode_b <= 3'h0;
    end else if (io_validin) begin
      mulAddRecFNToRaw_postMul_io_roundingMode_b <= io_roundingMode;
    end
    if (metaReset) begin
      roundingMode_stage0_b <= 3'h0;
    end else if (io_validin) begin
      roundingMode_stage0_b <= io_roundingMode;
    end
    if (metaReset) begin
      detectTininess_stage0_b <= 1'h0;
    end else begin
      detectTininess_stage0_b <= io_validin | detectTininess_stage0_b;
    end
    if (metaReset) begin
      valid_stage0_v <= 1'h0;
    end else if (reset) begin
      valid_stage0_v <= 1'h0;
    end else begin
      valid_stage0_v <= io_validin;
    end
    if (metaReset) begin
      roundRawFNToRecFN_io_invalidExc_b <= 1'h0;
    end else if (valid_stage0_v) begin
      roundRawFNToRecFN_io_invalidExc_b <= mulAddRecFNToRaw_postMul_io_invalidExc;
    end
    if (metaReset) begin
      roundRawFNToRecFN_io_in_b_isNaN <= 1'h0;
    end else if (valid_stage0_v) begin
      roundRawFNToRecFN_io_in_b_isNaN <= mulAddRecFNToRaw_postMul_io_rawOut_isNaN;
    end
    if (metaReset) begin
      roundRawFNToRecFN_io_in_b_isInf <= 1'h0;
    end else if (valid_stage0_v) begin
      roundRawFNToRecFN_io_in_b_isInf <= mulAddRecFNToRaw_postMul_io_rawOut_isInf;
    end
    if (metaReset) begin
      roundRawFNToRecFN_io_in_b_isZero <= 1'h0;
    end else if (valid_stage0_v) begin
      roundRawFNToRecFN_io_in_b_isZero <= mulAddRecFNToRaw_postMul_io_rawOut_isZero;
    end
    if (metaReset) begin
      roundRawFNToRecFN_io_in_b_sign <= 1'h0;
    end else if (valid_stage0_v) begin
      roundRawFNToRecFN_io_in_b_sign <= mulAddRecFNToRaw_postMul_io_rawOut_sign;
    end
    if (metaReset) begin
      roundRawFNToRecFN_io_in_b_sExp <= 10'h0;
    end else if (valid_stage0_v) begin
      roundRawFNToRecFN_io_in_b_sExp <= mulAddRecFNToRaw_postMul_io_rawOut_sExp;
    end
    if (metaReset) begin
      roundRawFNToRecFN_io_in_b_sig <= 27'h0;
    end else if (valid_stage0_v) begin
      roundRawFNToRecFN_io_in_b_sig <= mulAddRecFNToRaw_postMul_io_rawOut_sig;
    end
    if (metaReset) begin
      roundRawFNToRecFN_io_roundingMode_b <= 3'h0;
    end else if (valid_stage0_v) begin
      roundRawFNToRecFN_io_roundingMode_b <= roundingMode_stage0_b;
    end
    if (metaReset) begin
      roundRawFNToRecFN_io_detectTininess_b <= 1'h0;
    end else if (valid_stage0_v) begin
      roundRawFNToRecFN_io_detectTininess_b <= detectTininess_stage0_b;
    end
    MulAddRecFNPipe_state <= valid_stage0_v_pad;
    if (!(MulAddRecFNPipe_cov_read_data)) begin
      MulAddRecFNPipe_covSum <= MulAddRecFNPipe_covSum + 1'h1;
    end
    if (metaReset) begin
      MulAddRecFNPipe_metaAssert <= 1'h0;
    end else begin
      MulAddRecFNPipe_metaAssert <= MulAddRecFNPipe_metaAssert | MulAddRecFNPipe_or0;
    end
  end
  always @(posedge clock) begin
    if(MulAddRecFNPipe_cov_write_en & MulAddRecFNPipe_cov_write_mask) begin
      MulAddRecFNPipe_cov[MulAddRecFNPipe_cov_write_addr] <= MulAddRecFNPipe_cov_write_data; // @[Coverage map for MulAddRecFNPipe]
    end
  end
endmodule
module CompareRecFN(
  input  [64:0] io_a,
  input  [64:0] io_b,
  input         io_signaling,
  output        io_lt,
  output        io_eq,
  output [4:0]  io_exceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire [11:0] rawA_exp; // @[rawFloatFromRecFN.scala 50:21]
  wire  rawA_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  rawA_isSpecial; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawA__isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawA__isInf; // @[rawFloatFromRecFN.scala 56:33]
  wire  rawA__sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [12:0] rawA__sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire  rawA_out_sig_hi_lo; // @[rawFloatFromRecFN.scala 60:39]
  wire [51:0] rawA_out_sig_lo; // @[rawFloatFromRecFN.scala 60:51]
  wire [53:0] rawA__sig; // @[Cat.scala 30:58]
  wire [11:0] rawB_exp; // @[rawFloatFromRecFN.scala 50:21]
  wire  rawB_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  rawB_isSpecial; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawB__isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawB__isInf; // @[rawFloatFromRecFN.scala 56:33]
  wire  rawB__sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [12:0] rawB__sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire  rawB_out_sig_hi_lo; // @[rawFloatFromRecFN.scala 60:39]
  wire [51:0] rawB_out_sig_lo; // @[rawFloatFromRecFN.scala 60:51]
  wire [53:0] rawB__sig; // @[Cat.scala 30:58]
  wire  ordered; // @[CompareRecFN.scala 57:32]
  wire  bothInfs; // @[CompareRecFN.scala 58:33]
  wire  bothZeros; // @[CompareRecFN.scala 59:33]
  wire  eqExps; // @[CompareRecFN.scala 60:29]
  wire  _common_ltMags_T; // @[CompareRecFN.scala 62:20]
  wire  _common_ltMags_T_1; // @[CompareRecFN.scala 62:57]
  wire  _common_ltMags_T_2; // @[CompareRecFN.scala 62:44]
  wire  common_ltMags; // @[CompareRecFN.scala 62:33]
  wire  _common_eqMags_T; // @[CompareRecFN.scala 63:45]
  wire  common_eqMags; // @[CompareRecFN.scala 63:32]
  wire  _ordered_lt_T_2; // @[CompareRecFN.scala 67:25]
  wire  _ordered_lt_T_5; // @[CompareRecFN.scala 69:35]
  wire  _ordered_lt_T_7; // @[CompareRecFN.scala 69:54]
  wire  _ordered_lt_T_9; // @[CompareRecFN.scala 70:41]
  wire  _ordered_lt_T_10; // @[CompareRecFN.scala 69:74]
  wire  _ordered_lt_T_11; // @[CompareRecFN.scala 68:30]
  wire  _ordered_lt_T_12; // @[CompareRecFN.scala 67:41]
  wire  ordered_lt; // @[CompareRecFN.scala 66:21]
  wire  _ordered_eq_T; // @[CompareRecFN.scala 72:34]
  wire  _ordered_eq_T_1; // @[CompareRecFN.scala 72:62]
  wire  _ordered_eq_T_2; // @[CompareRecFN.scala 72:49]
  wire  ordered_eq; // @[CompareRecFN.scala 72:19]
  wire  _invalid_T_2; // @[common.scala 81:46]
  wire  _invalid_T_5; // @[common.scala 81:46]
  wire  _invalid_T_6; // @[CompareRecFN.scala 75:32]
  wire  _invalid_T_8; // @[CompareRecFN.scala 76:27]
  wire  invalid; // @[CompareRecFN.scala 75:58]
  wire [29:0] CompareRecFN_covSum;
  assign rawA_exp = io_a[63:52]; // @[rawFloatFromRecFN.scala 50:21]
  assign rawA_isZero = rawA_exp[11:9] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign rawA_isSpecial = rawA_exp[11:10] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawA__isNaN = rawA_isSpecial & rawA_exp[9]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawA__isInf = rawA_isSpecial & ~rawA_exp[9]; // @[rawFloatFromRecFN.scala 56:33]
  assign rawA__sign = io_a[64]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawA__sExp = {1'b0,$signed(rawA_exp)}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawA_out_sig_hi_lo = ~rawA_isZero; // @[rawFloatFromRecFN.scala 60:39]
  assign rawA_out_sig_lo = io_a[51:0]; // @[rawFloatFromRecFN.scala 60:51]
  assign rawA__sig = {1'h0,rawA_out_sig_hi_lo,rawA_out_sig_lo}; // @[Cat.scala 30:58]
  assign rawB_exp = io_b[63:52]; // @[rawFloatFromRecFN.scala 50:21]
  assign rawB_isZero = rawB_exp[11:9] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign rawB_isSpecial = rawB_exp[11:10] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawB__isNaN = rawB_isSpecial & rawB_exp[9]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawB__isInf = rawB_isSpecial & ~rawB_exp[9]; // @[rawFloatFromRecFN.scala 56:33]
  assign rawB__sign = io_b[64]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawB__sExp = {1'b0,$signed(rawB_exp)}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawB_out_sig_hi_lo = ~rawB_isZero; // @[rawFloatFromRecFN.scala 60:39]
  assign rawB_out_sig_lo = io_b[51:0]; // @[rawFloatFromRecFN.scala 60:51]
  assign rawB__sig = {1'h0,rawB_out_sig_hi_lo,rawB_out_sig_lo}; // @[Cat.scala 30:58]
  assign ordered = ~rawA__isNaN & ~rawB__isNaN; // @[CompareRecFN.scala 57:32]
  assign bothInfs = rawA__isInf & rawB__isInf; // @[CompareRecFN.scala 58:33]
  assign bothZeros = rawA_isZero & rawB_isZero; // @[CompareRecFN.scala 59:33]
  assign eqExps = $signed(rawA__sExp) == $signed(rawB__sExp); // @[CompareRecFN.scala 60:29]
  assign _common_ltMags_T = $signed(rawA__sExp) < $signed(rawB__sExp); // @[CompareRecFN.scala 62:20]
  assign _common_ltMags_T_1 = rawA__sig < rawB__sig; // @[CompareRecFN.scala 62:57]
  assign _common_ltMags_T_2 = eqExps & _common_ltMags_T_1; // @[CompareRecFN.scala 62:44]
  assign common_ltMags = _common_ltMags_T | _common_ltMags_T_2; // @[CompareRecFN.scala 62:33]
  assign _common_eqMags_T = rawA__sig == rawB__sig; // @[CompareRecFN.scala 63:45]
  assign common_eqMags = eqExps & _common_eqMags_T; // @[CompareRecFN.scala 63:32]
  assign _ordered_lt_T_2 = rawA__sign & ~rawB__sign; // @[CompareRecFN.scala 67:25]
  assign _ordered_lt_T_5 = rawA__sign & ~common_ltMags; // @[CompareRecFN.scala 69:35]
  assign _ordered_lt_T_7 = _ordered_lt_T_5 & ~common_eqMags; // @[CompareRecFN.scala 69:54]
  assign _ordered_lt_T_9 = ~rawB__sign & common_ltMags; // @[CompareRecFN.scala 70:41]
  assign _ordered_lt_T_10 = _ordered_lt_T_7 | _ordered_lt_T_9; // @[CompareRecFN.scala 69:74]
  assign _ordered_lt_T_11 = ~bothInfs & _ordered_lt_T_10; // @[CompareRecFN.scala 68:30]
  assign _ordered_lt_T_12 = _ordered_lt_T_2 | _ordered_lt_T_11; // @[CompareRecFN.scala 67:41]
  assign ordered_lt = ~bothZeros & _ordered_lt_T_12; // @[CompareRecFN.scala 66:21]
  assign _ordered_eq_T = rawA__sign == rawB__sign; // @[CompareRecFN.scala 72:34]
  assign _ordered_eq_T_1 = bothInfs | common_eqMags; // @[CompareRecFN.scala 72:62]
  assign _ordered_eq_T_2 = _ordered_eq_T & _ordered_eq_T_1; // @[CompareRecFN.scala 72:49]
  assign ordered_eq = bothZeros | _ordered_eq_T_2; // @[CompareRecFN.scala 72:19]
  assign _invalid_T_2 = rawA__isNaN & ~rawA__sig[51]; // @[common.scala 81:46]
  assign _invalid_T_5 = rawB__isNaN & ~rawB__sig[51]; // @[common.scala 81:46]
  assign _invalid_T_6 = _invalid_T_2 | _invalid_T_5; // @[CompareRecFN.scala 75:32]
  assign _invalid_T_8 = io_signaling & ~ordered; // @[CompareRecFN.scala 76:27]
  assign invalid = _invalid_T_6 | _invalid_T_8; // @[CompareRecFN.scala 75:58]
  assign io_lt = ordered & ordered_lt; // @[CompareRecFN.scala 78:11]
  assign io_eq = ordered & ordered_eq; // @[CompareRecFN.scala 79:11]
  assign io_exceptionFlags = {invalid,4'h0}; // @[CompareRecFN.scala 81:23]
  assign CompareRecFN_covSum = 30'h0;
  assign io_covSum = CompareRecFN_covSum;
  assign metaAssert = 1'h0;
endmodule
module RecFNToIN(
  input  [64:0] io_in,
  input  [2:0]  io_roundingMode,
  input         io_signedOut,
  output [63:0] io_out,
  output [2:0]  io_intExceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire [11:0] rawIn_exp; // @[rawFloatFromRecFN.scala 50:21]
  wire  rawIn_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  rawIn_isSpecial; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawIn__isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawIn__isInf; // @[rawFloatFromRecFN.scala 56:33]
  wire  rawIn__sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [12:0] rawIn__sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire  rawIn_out_sig_hi_lo; // @[rawFloatFromRecFN.scala 60:39]
  wire [51:0] rawIn_out_sig_lo; // @[rawFloatFromRecFN.scala 60:51]
  wire [53:0] rawIn__sig; // @[Cat.scala 30:58]
  wire  magGeOne; // @[RecFNToIN.scala 58:30]
  wire [10:0] posExp; // @[RecFNToIN.scala 59:28]
  wire  _magJustBelowOne_T_1; // @[RecFNToIN.scala 60:47]
  wire  magJustBelowOne; // @[RecFNToIN.scala 60:37]
  wire  roundingMode_near_even; // @[RecFNToIN.scala 64:53]
  wire  roundingMode_min; // @[RecFNToIN.scala 66:53]
  wire  roundingMode_max; // @[RecFNToIN.scala 67:53]
  wire  roundingMode_near_maxMag; // @[RecFNToIN.scala 68:53]
  wire  roundingMode_odd; // @[RecFNToIN.scala 69:53]
  wire [51:0] shiftedSig_lo; // @[RecFNToIN.scala 80:32]
  wire [52:0] _shiftedSig_T; // @[Cat.scala 30:58]
  wire [5:0] _shiftedSig_T_2; // @[RecFNToIN.scala 81:16]
  wire [115:0] _GEN_0; // @[RecFNToIN.scala 80:50]
  wire [115:0] shiftedSig; // @[RecFNToIN.scala 80:50]
  wire [64:0] alignedSig_hi; // @[RecFNToIN.scala 86:23]
  wire  alignedSig_lo; // @[RecFNToIN.scala 86:69]
  wire [65:0] alignedSig; // @[Cat.scala 30:58]
  wire [63:0] unroundedInt; // @[RecFNToIN.scala 87:54]
  wire  _common_inexact_T_1; // @[RecFNToIN.scala 89:57]
  wire  common_inexact; // @[RecFNToIN.scala 89:29]
  wire  _roundIncr_near_even_T_1; // @[RecFNToIN.scala 91:46]
  wire  _roundIncr_near_even_T_3; // @[RecFNToIN.scala 91:71]
  wire  _roundIncr_near_even_T_4; // @[RecFNToIN.scala 91:51]
  wire  _roundIncr_near_even_T_5; // @[RecFNToIN.scala 91:25]
  wire  _roundIncr_near_even_T_8; // @[RecFNToIN.scala 92:26]
  wire  roundIncr_near_even; // @[RecFNToIN.scala 91:78]
  wire  _roundIncr_near_maxMag_T_1; // @[RecFNToIN.scala 93:43]
  wire  roundIncr_near_maxMag; // @[RecFNToIN.scala 93:61]
  wire  _roundIncr_T; // @[RecFNToIN.scala 95:35]
  wire  _roundIncr_T_1; // @[RecFNToIN.scala 96:35]
  wire  _roundIncr_T_2; // @[RecFNToIN.scala 95:61]
  wire  _roundIncr_T_3; // @[RecFNToIN.scala 97:28]
  wire  _roundIncr_T_4; // @[RecFNToIN.scala 98:26]
  wire  _roundIncr_T_5; // @[RecFNToIN.scala 97:49]
  wire  _roundIncr_T_6; // @[RecFNToIN.scala 96:61]
  wire  _roundIncr_T_8; // @[RecFNToIN.scala 99:43]
  wire  _roundIncr_T_9; // @[RecFNToIN.scala 99:27]
  wire  roundIncr; // @[RecFNToIN.scala 98:46]
  wire [63:0] complUnroundedInt; // @[RecFNToIN.scala 100:32]
  wire  _roundedInt_T; // @[RecFNToIN.scala 102:23]
  wire [63:0] _roundedInt_T_2; // @[RecFNToIN.scala 103:31]
  wire [63:0] _roundedInt_T_3; // @[RecFNToIN.scala 102:12]
  wire  _roundedInt_T_4; // @[RecFNToIN.scala 105:31]
  wire [63:0] _GEN_1; // @[RecFNToIN.scala 105:11]
  wire [63:0] roundedInt; // @[RecFNToIN.scala 105:11]
  wire  magGeOne_atOverflowEdge; // @[RecFNToIN.scala 107:43]
  wire  _roundCarryBut2_T_1; // @[RecFNToIN.scala 110:56]
  wire  roundCarryBut2; // @[RecFNToIN.scala 110:61]
  wire  _common_overflow_T; // @[RecFNToIN.scala 113:21]
  wire  _common_overflow_T_2; // @[RecFNToIN.scala 117:60]
  wire  _common_overflow_T_3; // @[RecFNToIN.scala 117:64]
  wire  _common_overflow_T_4; // @[RecFNToIN.scala 116:49]
  wire  _common_overflow_T_5; // @[RecFNToIN.scala 119:38]
  wire  _common_overflow_T_6; // @[RecFNToIN.scala 119:62]
  wire  _common_overflow_T_7; // @[RecFNToIN.scala 118:49]
  wire  _common_overflow_T_8; // @[RecFNToIN.scala 115:24]
  wire  _common_overflow_T_10; // @[RecFNToIN.scala 122:50]
  wire  _common_overflow_T_11; // @[RecFNToIN.scala 123:57]
  wire  _common_overflow_T_12; // @[RecFNToIN.scala 121:32]
  wire  _common_overflow_T_13; // @[RecFNToIN.scala 114:20]
  wire  _common_overflow_T_14; // @[RecFNToIN.scala 113:40]
  wire  _common_overflow_T_16; // @[RecFNToIN.scala 125:27]
  wire  _common_overflow_T_17; // @[RecFNToIN.scala 125:41]
  wire  common_overflow; // @[RecFNToIN.scala 112:12]
  wire  invalidExc; // @[RecFNToIN.scala 130:34]
  wire  overflow; // @[RecFNToIN.scala 131:32]
  wire  _inexact_T_2; // @[RecFNToIN.scala 132:32]
  wire  inexact; // @[RecFNToIN.scala 132:52]
  wire  excSign; // @[RecFNToIN.scala 134:32]
  wire  _excOut_T; // @[RecFNToIN.scala 136:27]
  wire [63:0] _excOut_T_1; // @[RecFNToIN.scala 136:12]
  wire [62:0] _excOut_T_3; // @[RecFNToIN.scala 140:12]
  wire [63:0] _GEN_2; // @[RecFNToIN.scala 139:11]
  wire [63:0] excOut; // @[RecFNToIN.scala 139:11]
  wire  _io_out_T; // @[RecFNToIN.scala 142:30]
  wire [1:0] io_intExceptionFlags_hi; // @[Cat.scala 30:58]
  wire [29:0] RecFNToIN_covSum;
  assign rawIn_exp = io_in[63:52]; // @[rawFloatFromRecFN.scala 50:21]
  assign rawIn_isZero = rawIn_exp[11:9] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign rawIn_isSpecial = rawIn_exp[11:10] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawIn__isNaN = rawIn_isSpecial & rawIn_exp[9]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawIn__isInf = rawIn_isSpecial & ~rawIn_exp[9]; // @[rawFloatFromRecFN.scala 56:33]
  assign rawIn__sign = io_in[64]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawIn__sExp = {1'b0,$signed(rawIn_exp)}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawIn_out_sig_hi_lo = ~rawIn_isZero; // @[rawFloatFromRecFN.scala 60:39]
  assign rawIn_out_sig_lo = io_in[51:0]; // @[rawFloatFromRecFN.scala 60:51]
  assign rawIn__sig = {1'h0,rawIn_out_sig_hi_lo,rawIn_out_sig_lo}; // @[Cat.scala 30:58]
  assign magGeOne = rawIn__sExp[11]; // @[RecFNToIN.scala 58:30]
  assign posExp = rawIn__sExp[10:0]; // @[RecFNToIN.scala 59:28]
  assign _magJustBelowOne_T_1 = &posExp; // @[RecFNToIN.scala 60:47]
  assign magJustBelowOne = ~magGeOne & _magJustBelowOne_T_1; // @[RecFNToIN.scala 60:37]
  assign roundingMode_near_even = io_roundingMode == 3'h0; // @[RecFNToIN.scala 64:53]
  assign roundingMode_min = io_roundingMode == 3'h2; // @[RecFNToIN.scala 66:53]
  assign roundingMode_max = io_roundingMode == 3'h3; // @[RecFNToIN.scala 67:53]
  assign roundingMode_near_maxMag = io_roundingMode == 3'h4; // @[RecFNToIN.scala 68:53]
  assign roundingMode_odd = io_roundingMode == 3'h6; // @[RecFNToIN.scala 69:53]
  assign shiftedSig_lo = rawIn__sig[51:0]; // @[RecFNToIN.scala 80:32]
  assign _shiftedSig_T = {magGeOne,shiftedSig_lo}; // @[Cat.scala 30:58]
  assign _shiftedSig_T_2 = magGeOne ? rawIn__sExp[5:0] : 6'h0; // @[RecFNToIN.scala 81:16]
  assign _GEN_0 = {{63'd0}, _shiftedSig_T}; // @[RecFNToIN.scala 80:50]
  assign shiftedSig = _GEN_0 << _shiftedSig_T_2; // @[RecFNToIN.scala 80:50]
  assign alignedSig_hi = shiftedSig[115:51]; // @[RecFNToIN.scala 86:23]
  assign alignedSig_lo = |shiftedSig[50:0]; // @[RecFNToIN.scala 86:69]
  assign alignedSig = {alignedSig_hi,alignedSig_lo}; // @[Cat.scala 30:58]
  assign unroundedInt = alignedSig[65:2]; // @[RecFNToIN.scala 87:54]
  assign _common_inexact_T_1 = |alignedSig[1:0]; // @[RecFNToIN.scala 89:57]
  assign common_inexact = magGeOne ? _common_inexact_T_1 : rawIn_out_sig_hi_lo; // @[RecFNToIN.scala 89:29]
  assign _roundIncr_near_even_T_1 = &alignedSig[2:1]; // @[RecFNToIN.scala 91:46]
  assign _roundIncr_near_even_T_3 = &alignedSig[1:0]; // @[RecFNToIN.scala 91:71]
  assign _roundIncr_near_even_T_4 = _roundIncr_near_even_T_1 | _roundIncr_near_even_T_3; // @[RecFNToIN.scala 91:51]
  assign _roundIncr_near_even_T_5 = magGeOne & _roundIncr_near_even_T_4; // @[RecFNToIN.scala 91:25]
  assign _roundIncr_near_even_T_8 = magJustBelowOne & _common_inexact_T_1; // @[RecFNToIN.scala 92:26]
  assign roundIncr_near_even = _roundIncr_near_even_T_5 | _roundIncr_near_even_T_8; // @[RecFNToIN.scala 91:78]
  assign _roundIncr_near_maxMag_T_1 = magGeOne & alignedSig[1]; // @[RecFNToIN.scala 93:43]
  assign roundIncr_near_maxMag = _roundIncr_near_maxMag_T_1 | magJustBelowOne; // @[RecFNToIN.scala 93:61]
  assign _roundIncr_T = roundingMode_near_even & roundIncr_near_even; // @[RecFNToIN.scala 95:35]
  assign _roundIncr_T_1 = roundingMode_near_maxMag & roundIncr_near_maxMag; // @[RecFNToIN.scala 96:35]
  assign _roundIncr_T_2 = _roundIncr_T | _roundIncr_T_1; // @[RecFNToIN.scala 95:61]
  assign _roundIncr_T_3 = roundingMode_min | roundingMode_odd; // @[RecFNToIN.scala 97:28]
  assign _roundIncr_T_4 = rawIn__sign & common_inexact; // @[RecFNToIN.scala 98:26]
  assign _roundIncr_T_5 = _roundIncr_T_3 & _roundIncr_T_4; // @[RecFNToIN.scala 97:49]
  assign _roundIncr_T_6 = _roundIncr_T_2 | _roundIncr_T_5; // @[RecFNToIN.scala 96:61]
  assign _roundIncr_T_8 = ~rawIn__sign & common_inexact; // @[RecFNToIN.scala 99:43]
  assign _roundIncr_T_9 = roundingMode_max & _roundIncr_T_8; // @[RecFNToIN.scala 99:27]
  assign roundIncr = _roundIncr_T_6 | _roundIncr_T_9; // @[RecFNToIN.scala 98:46]
  assign complUnroundedInt = rawIn__sign ? ~unroundedInt : unroundedInt; // @[RecFNToIN.scala 100:32]
  assign _roundedInt_T = roundIncr ^ rawIn__sign; // @[RecFNToIN.scala 102:23]
  assign _roundedInt_T_2 = complUnroundedInt + 64'h1; // @[RecFNToIN.scala 103:31]
  assign _roundedInt_T_3 = _roundedInt_T ? _roundedInt_T_2 : complUnroundedInt; // @[RecFNToIN.scala 102:12]
  assign _roundedInt_T_4 = roundingMode_odd & common_inexact; // @[RecFNToIN.scala 105:31]
  assign _GEN_1 = {{63'd0}, _roundedInt_T_4}; // @[RecFNToIN.scala 105:11]
  assign roundedInt = _roundedInt_T_3 | _GEN_1; // @[RecFNToIN.scala 105:11]
  assign magGeOne_atOverflowEdge = posExp == 11'h3f; // @[RecFNToIN.scala 107:43]
  assign _roundCarryBut2_T_1 = &unroundedInt[61:0]; // @[RecFNToIN.scala 110:56]
  assign roundCarryBut2 = _roundCarryBut2_T_1 & roundIncr; // @[RecFNToIN.scala 110:61]
  assign _common_overflow_T = posExp >= 11'h40; // @[RecFNToIN.scala 113:21]
  assign _common_overflow_T_2 = |unroundedInt[62:0]; // @[RecFNToIN.scala 117:60]
  assign _common_overflow_T_3 = _common_overflow_T_2 | roundIncr; // @[RecFNToIN.scala 117:64]
  assign _common_overflow_T_4 = magGeOne_atOverflowEdge & _common_overflow_T_3; // @[RecFNToIN.scala 116:49]
  assign _common_overflow_T_5 = posExp == 11'h3e; // @[RecFNToIN.scala 119:38]
  assign _common_overflow_T_6 = _common_overflow_T_5 & roundCarryBut2; // @[RecFNToIN.scala 119:62]
  assign _common_overflow_T_7 = magGeOne_atOverflowEdge | _common_overflow_T_6; // @[RecFNToIN.scala 118:49]
  assign _common_overflow_T_8 = rawIn__sign ? _common_overflow_T_4 : _common_overflow_T_7; // @[RecFNToIN.scala 115:24]
  assign _common_overflow_T_10 = magGeOne_atOverflowEdge & unroundedInt[62]; // @[RecFNToIN.scala 122:50]
  assign _common_overflow_T_11 = _common_overflow_T_10 & roundCarryBut2; // @[RecFNToIN.scala 123:57]
  assign _common_overflow_T_12 = rawIn__sign | _common_overflow_T_11; // @[RecFNToIN.scala 121:32]
  assign _common_overflow_T_13 = io_signedOut ? _common_overflow_T_8 : _common_overflow_T_12; // @[RecFNToIN.scala 114:20]
  assign _common_overflow_T_14 = _common_overflow_T | _common_overflow_T_13; // @[RecFNToIN.scala 113:40]
  assign _common_overflow_T_16 = ~io_signedOut & rawIn__sign; // @[RecFNToIN.scala 125:27]
  assign _common_overflow_T_17 = _common_overflow_T_16 & roundIncr; // @[RecFNToIN.scala 125:41]
  assign common_overflow = magGeOne ? _common_overflow_T_14 : _common_overflow_T_17; // @[RecFNToIN.scala 112:12]
  assign invalidExc = rawIn__isNaN | rawIn__isInf; // @[RecFNToIN.scala 130:34]
  assign overflow = ~invalidExc & common_overflow; // @[RecFNToIN.scala 131:32]
  assign _inexact_T_2 = ~invalidExc & ~common_overflow; // @[RecFNToIN.scala 132:32]
  assign inexact = _inexact_T_2 & common_inexact; // @[RecFNToIN.scala 132:52]
  assign excSign = ~rawIn__isNaN & rawIn__sign; // @[RecFNToIN.scala 134:32]
  assign _excOut_T = io_signedOut == excSign; // @[RecFNToIN.scala 136:27]
  assign _excOut_T_1 = _excOut_T ? 64'h8000000000000000 : 64'h0; // @[RecFNToIN.scala 136:12]
  assign _excOut_T_3 = excSign ? 63'h0 : 63'h7fffffffffffffff; // @[RecFNToIN.scala 140:12]
  assign _GEN_2 = {{1'd0}, _excOut_T_3}; // @[RecFNToIN.scala 139:11]
  assign excOut = _excOut_T_1 | _GEN_2; // @[RecFNToIN.scala 139:11]
  assign _io_out_T = invalidExc | common_overflow; // @[RecFNToIN.scala 142:30]
  assign io_intExceptionFlags_hi = {invalidExc,overflow}; // @[Cat.scala 30:58]
  assign io_out = _io_out_T ? excOut : roundedInt; // @[RecFNToIN.scala 142:12]
  assign io_intExceptionFlags = {io_intExceptionFlags_hi,inexact}; // @[RecFNToIN.scala 143:26]
  assign RecFNToIN_covSum = 30'h0;
  assign io_covSum = RecFNToIN_covSum;
  assign metaAssert = 1'h0;
endmodule
module RecFNToIN_1(
  input  [64:0] io_in,
  input  [2:0]  io_roundingMode,
  input         io_signedOut,
  output [2:0]  io_intExceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire [11:0] rawIn_exp; // @[rawFloatFromRecFN.scala 50:21]
  wire  rawIn_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  rawIn_isSpecial; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawIn__isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawIn__isInf; // @[rawFloatFromRecFN.scala 56:33]
  wire  rawIn__sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [12:0] rawIn__sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire  rawIn_out_sig_hi_lo; // @[rawFloatFromRecFN.scala 60:39]
  wire [51:0] rawIn_out_sig_lo; // @[rawFloatFromRecFN.scala 60:51]
  wire [53:0] rawIn__sig; // @[Cat.scala 30:58]
  wire  magGeOne; // @[RecFNToIN.scala 58:30]
  wire [10:0] posExp; // @[RecFNToIN.scala 59:28]
  wire  _magJustBelowOne_T_1; // @[RecFNToIN.scala 60:47]
  wire  magJustBelowOne; // @[RecFNToIN.scala 60:37]
  wire  roundingMode_near_even; // @[RecFNToIN.scala 64:53]
  wire  roundingMode_min; // @[RecFNToIN.scala 66:53]
  wire  roundingMode_max; // @[RecFNToIN.scala 67:53]
  wire  roundingMode_near_maxMag; // @[RecFNToIN.scala 68:53]
  wire  roundingMode_odd; // @[RecFNToIN.scala 69:53]
  wire [51:0] shiftedSig_lo; // @[RecFNToIN.scala 80:32]
  wire [52:0] _shiftedSig_T; // @[Cat.scala 30:58]
  wire [4:0] _shiftedSig_T_2; // @[RecFNToIN.scala 81:16]
  wire [83:0] _GEN_0; // @[RecFNToIN.scala 80:50]
  wire [83:0] shiftedSig; // @[RecFNToIN.scala 80:50]
  wire [32:0] alignedSig_hi; // @[RecFNToIN.scala 86:23]
  wire  alignedSig_lo; // @[RecFNToIN.scala 86:69]
  wire [33:0] alignedSig; // @[Cat.scala 30:58]
  wire [31:0] unroundedInt; // @[RecFNToIN.scala 87:54]
  wire  _common_inexact_T_1; // @[RecFNToIN.scala 89:57]
  wire  common_inexact; // @[RecFNToIN.scala 89:29]
  wire  _roundIncr_near_even_T_1; // @[RecFNToIN.scala 91:46]
  wire  _roundIncr_near_even_T_3; // @[RecFNToIN.scala 91:71]
  wire  _roundIncr_near_even_T_4; // @[RecFNToIN.scala 91:51]
  wire  _roundIncr_near_even_T_5; // @[RecFNToIN.scala 91:25]
  wire  _roundIncr_near_even_T_8; // @[RecFNToIN.scala 92:26]
  wire  roundIncr_near_even; // @[RecFNToIN.scala 91:78]
  wire  _roundIncr_near_maxMag_T_1; // @[RecFNToIN.scala 93:43]
  wire  roundIncr_near_maxMag; // @[RecFNToIN.scala 93:61]
  wire  _roundIncr_T; // @[RecFNToIN.scala 95:35]
  wire  _roundIncr_T_1; // @[RecFNToIN.scala 96:35]
  wire  _roundIncr_T_2; // @[RecFNToIN.scala 95:61]
  wire  _roundIncr_T_3; // @[RecFNToIN.scala 97:28]
  wire  _roundIncr_T_4; // @[RecFNToIN.scala 98:26]
  wire  _roundIncr_T_5; // @[RecFNToIN.scala 97:49]
  wire  _roundIncr_T_6; // @[RecFNToIN.scala 96:61]
  wire  _roundIncr_T_8; // @[RecFNToIN.scala 99:43]
  wire  _roundIncr_T_9; // @[RecFNToIN.scala 99:27]
  wire  roundIncr; // @[RecFNToIN.scala 98:46]
  wire  magGeOne_atOverflowEdge; // @[RecFNToIN.scala 107:43]
  wire  _roundCarryBut2_T_1; // @[RecFNToIN.scala 110:56]
  wire  roundCarryBut2; // @[RecFNToIN.scala 110:61]
  wire  _common_overflow_T; // @[RecFNToIN.scala 113:21]
  wire  _common_overflow_T_2; // @[RecFNToIN.scala 117:60]
  wire  _common_overflow_T_3; // @[RecFNToIN.scala 117:64]
  wire  _common_overflow_T_4; // @[RecFNToIN.scala 116:49]
  wire  _common_overflow_T_5; // @[RecFNToIN.scala 119:38]
  wire  _common_overflow_T_6; // @[RecFNToIN.scala 119:62]
  wire  _common_overflow_T_7; // @[RecFNToIN.scala 118:49]
  wire  _common_overflow_T_8; // @[RecFNToIN.scala 115:24]
  wire  _common_overflow_T_10; // @[RecFNToIN.scala 122:50]
  wire  _common_overflow_T_11; // @[RecFNToIN.scala 123:57]
  wire  _common_overflow_T_12; // @[RecFNToIN.scala 121:32]
  wire  _common_overflow_T_13; // @[RecFNToIN.scala 114:20]
  wire  _common_overflow_T_14; // @[RecFNToIN.scala 113:40]
  wire  _common_overflow_T_16; // @[RecFNToIN.scala 125:27]
  wire  _common_overflow_T_17; // @[RecFNToIN.scala 125:41]
  wire  common_overflow; // @[RecFNToIN.scala 112:12]
  wire  invalidExc; // @[RecFNToIN.scala 130:34]
  wire  overflow; // @[RecFNToIN.scala 131:32]
  wire  _inexact_T_2; // @[RecFNToIN.scala 132:32]
  wire  inexact; // @[RecFNToIN.scala 132:52]
  wire [1:0] io_intExceptionFlags_hi; // @[Cat.scala 30:58]
  wire [29:0] RecFNToIN_1_covSum;
  assign rawIn_exp = io_in[63:52]; // @[rawFloatFromRecFN.scala 50:21]
  assign rawIn_isZero = rawIn_exp[11:9] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign rawIn_isSpecial = rawIn_exp[11:10] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawIn__isNaN = rawIn_isSpecial & rawIn_exp[9]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawIn__isInf = rawIn_isSpecial & ~rawIn_exp[9]; // @[rawFloatFromRecFN.scala 56:33]
  assign rawIn__sign = io_in[64]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawIn__sExp = {1'b0,$signed(rawIn_exp)}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawIn_out_sig_hi_lo = ~rawIn_isZero; // @[rawFloatFromRecFN.scala 60:39]
  assign rawIn_out_sig_lo = io_in[51:0]; // @[rawFloatFromRecFN.scala 60:51]
  assign rawIn__sig = {1'h0,rawIn_out_sig_hi_lo,rawIn_out_sig_lo}; // @[Cat.scala 30:58]
  assign magGeOne = rawIn__sExp[11]; // @[RecFNToIN.scala 58:30]
  assign posExp = rawIn__sExp[10:0]; // @[RecFNToIN.scala 59:28]
  assign _magJustBelowOne_T_1 = &posExp; // @[RecFNToIN.scala 60:47]
  assign magJustBelowOne = ~magGeOne & _magJustBelowOne_T_1; // @[RecFNToIN.scala 60:37]
  assign roundingMode_near_even = io_roundingMode == 3'h0; // @[RecFNToIN.scala 64:53]
  assign roundingMode_min = io_roundingMode == 3'h2; // @[RecFNToIN.scala 66:53]
  assign roundingMode_max = io_roundingMode == 3'h3; // @[RecFNToIN.scala 67:53]
  assign roundingMode_near_maxMag = io_roundingMode == 3'h4; // @[RecFNToIN.scala 68:53]
  assign roundingMode_odd = io_roundingMode == 3'h6; // @[RecFNToIN.scala 69:53]
  assign shiftedSig_lo = rawIn__sig[51:0]; // @[RecFNToIN.scala 80:32]
  assign _shiftedSig_T = {magGeOne,shiftedSig_lo}; // @[Cat.scala 30:58]
  assign _shiftedSig_T_2 = magGeOne ? rawIn__sExp[4:0] : 5'h0; // @[RecFNToIN.scala 81:16]
  assign _GEN_0 = {{31'd0}, _shiftedSig_T}; // @[RecFNToIN.scala 80:50]
  assign shiftedSig = _GEN_0 << _shiftedSig_T_2; // @[RecFNToIN.scala 80:50]
  assign alignedSig_hi = shiftedSig[83:51]; // @[RecFNToIN.scala 86:23]
  assign alignedSig_lo = |shiftedSig[50:0]; // @[RecFNToIN.scala 86:69]
  assign alignedSig = {alignedSig_hi,alignedSig_lo}; // @[Cat.scala 30:58]
  assign unroundedInt = alignedSig[33:2]; // @[RecFNToIN.scala 87:54]
  assign _common_inexact_T_1 = |alignedSig[1:0]; // @[RecFNToIN.scala 89:57]
  assign common_inexact = magGeOne ? _common_inexact_T_1 : rawIn_out_sig_hi_lo; // @[RecFNToIN.scala 89:29]
  assign _roundIncr_near_even_T_1 = &alignedSig[2:1]; // @[RecFNToIN.scala 91:46]
  assign _roundIncr_near_even_T_3 = &alignedSig[1:0]; // @[RecFNToIN.scala 91:71]
  assign _roundIncr_near_even_T_4 = _roundIncr_near_even_T_1 | _roundIncr_near_even_T_3; // @[RecFNToIN.scala 91:51]
  assign _roundIncr_near_even_T_5 = magGeOne & _roundIncr_near_even_T_4; // @[RecFNToIN.scala 91:25]
  assign _roundIncr_near_even_T_8 = magJustBelowOne & _common_inexact_T_1; // @[RecFNToIN.scala 92:26]
  assign roundIncr_near_even = _roundIncr_near_even_T_5 | _roundIncr_near_even_T_8; // @[RecFNToIN.scala 91:78]
  assign _roundIncr_near_maxMag_T_1 = magGeOne & alignedSig[1]; // @[RecFNToIN.scala 93:43]
  assign roundIncr_near_maxMag = _roundIncr_near_maxMag_T_1 | magJustBelowOne; // @[RecFNToIN.scala 93:61]
  assign _roundIncr_T = roundingMode_near_even & roundIncr_near_even; // @[RecFNToIN.scala 95:35]
  assign _roundIncr_T_1 = roundingMode_near_maxMag & roundIncr_near_maxMag; // @[RecFNToIN.scala 96:35]
  assign _roundIncr_T_2 = _roundIncr_T | _roundIncr_T_1; // @[RecFNToIN.scala 95:61]
  assign _roundIncr_T_3 = roundingMode_min | roundingMode_odd; // @[RecFNToIN.scala 97:28]
  assign _roundIncr_T_4 = rawIn__sign & common_inexact; // @[RecFNToIN.scala 98:26]
  assign _roundIncr_T_5 = _roundIncr_T_3 & _roundIncr_T_4; // @[RecFNToIN.scala 97:49]
  assign _roundIncr_T_6 = _roundIncr_T_2 | _roundIncr_T_5; // @[RecFNToIN.scala 96:61]
  assign _roundIncr_T_8 = ~rawIn__sign & common_inexact; // @[RecFNToIN.scala 99:43]
  assign _roundIncr_T_9 = roundingMode_max & _roundIncr_T_8; // @[RecFNToIN.scala 99:27]
  assign roundIncr = _roundIncr_T_6 | _roundIncr_T_9; // @[RecFNToIN.scala 98:46]
  assign magGeOne_atOverflowEdge = posExp == 11'h1f; // @[RecFNToIN.scala 107:43]
  assign _roundCarryBut2_T_1 = &unroundedInt[29:0]; // @[RecFNToIN.scala 110:56]
  assign roundCarryBut2 = _roundCarryBut2_T_1 & roundIncr; // @[RecFNToIN.scala 110:61]
  assign _common_overflow_T = posExp >= 11'h20; // @[RecFNToIN.scala 113:21]
  assign _common_overflow_T_2 = |unroundedInt[30:0]; // @[RecFNToIN.scala 117:60]
  assign _common_overflow_T_3 = _common_overflow_T_2 | roundIncr; // @[RecFNToIN.scala 117:64]
  assign _common_overflow_T_4 = magGeOne_atOverflowEdge & _common_overflow_T_3; // @[RecFNToIN.scala 116:49]
  assign _common_overflow_T_5 = posExp == 11'h1e; // @[RecFNToIN.scala 119:38]
  assign _common_overflow_T_6 = _common_overflow_T_5 & roundCarryBut2; // @[RecFNToIN.scala 119:62]
  assign _common_overflow_T_7 = magGeOne_atOverflowEdge | _common_overflow_T_6; // @[RecFNToIN.scala 118:49]
  assign _common_overflow_T_8 = rawIn__sign ? _common_overflow_T_4 : _common_overflow_T_7; // @[RecFNToIN.scala 115:24]
  assign _common_overflow_T_10 = magGeOne_atOverflowEdge & unroundedInt[30]; // @[RecFNToIN.scala 122:50]
  assign _common_overflow_T_11 = _common_overflow_T_10 & roundCarryBut2; // @[RecFNToIN.scala 123:57]
  assign _common_overflow_T_12 = rawIn__sign | _common_overflow_T_11; // @[RecFNToIN.scala 121:32]
  assign _common_overflow_T_13 = io_signedOut ? _common_overflow_T_8 : _common_overflow_T_12; // @[RecFNToIN.scala 114:20]
  assign _common_overflow_T_14 = _common_overflow_T | _common_overflow_T_13; // @[RecFNToIN.scala 113:40]
  assign _common_overflow_T_16 = ~io_signedOut & rawIn__sign; // @[RecFNToIN.scala 125:27]
  assign _common_overflow_T_17 = _common_overflow_T_16 & roundIncr; // @[RecFNToIN.scala 125:41]
  assign common_overflow = magGeOne ? _common_overflow_T_14 : _common_overflow_T_17; // @[RecFNToIN.scala 112:12]
  assign invalidExc = rawIn__isNaN | rawIn__isInf; // @[RecFNToIN.scala 130:34]
  assign overflow = ~invalidExc & common_overflow; // @[RecFNToIN.scala 131:32]
  assign _inexact_T_2 = ~invalidExc & ~common_overflow; // @[RecFNToIN.scala 132:32]
  assign inexact = _inexact_T_2 & common_inexact; // @[RecFNToIN.scala 132:52]
  assign io_intExceptionFlags_hi = {invalidExc,overflow}; // @[Cat.scala 30:58]
  assign io_intExceptionFlags = {io_intExceptionFlags_hi,inexact}; // @[RecFNToIN.scala 143:26]
  assign RecFNToIN_1_covSum = 30'h0;
  assign io_covSum = RecFNToIN_1_covSum;
  assign metaAssert = 1'h0;
endmodule
module INToRecFN(
  input         io_signedIn,
  input  [63:0] io_in,
  input  [2:0]  io_roundingMode,
  output [32:0] io_out,
  output [4:0]  io_exceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  roundAnyRawFNToRecFN_io_in_isZero; // @[INToRecFN.scala 59:15]
  wire  roundAnyRawFNToRecFN_io_in_sign; // @[INToRecFN.scala 59:15]
  wire [8:0] roundAnyRawFNToRecFN_io_in_sExp; // @[INToRecFN.scala 59:15]
  wire [64:0] roundAnyRawFNToRecFN_io_in_sig; // @[INToRecFN.scala 59:15]
  wire [2:0] roundAnyRawFNToRecFN_io_roundingMode; // @[INToRecFN.scala 59:15]
  wire [32:0] roundAnyRawFNToRecFN_io_out; // @[INToRecFN.scala 59:15]
  wire [4:0] roundAnyRawFNToRecFN_io_exceptionFlags; // @[INToRecFN.scala 59:15]
  wire [29:0] roundAnyRawFNToRecFN_io_covSum; // @[INToRecFN.scala 59:15]
  wire  roundAnyRawFNToRecFN_metaAssert; // @[INToRecFN.scala 59:15]
  wire  intAsRawFloat_sign; // @[rawFloatFromIN.scala 50:29]
  wire [63:0] _intAsRawFloat_absIn_T_1; // @[rawFloatFromIN.scala 51:31]
  wire [63:0] intAsRawFloat_extAbsIn_lo; // @[rawFloatFromIN.scala 51:24]
  wire [127:0] _intAsRawFloat_extAbsIn_T; // @[Cat.scala 30:58]
  wire [63:0] intAsRawFloat_extAbsIn; // @[rawFloatFromIN.scala 52:56]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_64; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_65; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_66; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_67; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_68; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_69; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_70; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_71; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_72; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_73; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_74; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_75; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_76; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_77; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_78; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_79; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_80; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_81; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_82; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_83; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_84; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_85; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_86; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_87; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_88; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_89; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_90; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_91; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_92; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_93; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_94; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_95; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_96; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_97; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_98; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_99; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_100; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_101; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_102; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_103; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_104; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_105; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_106; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_107; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_108; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_109; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_110; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_111; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_112; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_113; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_114; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_115; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_116; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_117; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_118; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_119; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_120; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_121; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_122; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_123; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_124; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_125; // @[Mux.scala 47:69]
  wire [5:0] intAsRawFloat_adjustedNormDist; // @[Mux.scala 47:69]
  wire [126:0] _GEN_0; // @[rawFloatFromIN.scala 55:22]
  wire [126:0] _intAsRawFloat_sig_T; // @[rawFloatFromIN.scala 55:22]
  wire [63:0] intAsRawFloat_sig; // @[rawFloatFromIN.scala 55:41]
  wire [5:0] intAsRawFloat_out_sExp_lo; // @[rawFloatFromIN.scala 63:39]
  wire [7:0] _intAsRawFloat_out_sExp_T_1; // @[Cat.scala 30:58]
  wire [29:0] INToRecFN_covSum;
  wire [29:0] roundAnyRawFNToRecFN_sum;
  wire  roundAnyRawFNToRecFN_metaAssert_wire;
  RoundAnyRawFNToRecFN_1 roundAnyRawFNToRecFN ( // @[INToRecFN.scala 59:15]
    .io_in_isZero(roundAnyRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundAnyRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundAnyRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundAnyRawFNToRecFN_io_in_sig),
    .io_roundingMode(roundAnyRawFNToRecFN_io_roundingMode),
    .io_out(roundAnyRawFNToRecFN_io_out),
    .io_exceptionFlags(roundAnyRawFNToRecFN_io_exceptionFlags),
    .io_covSum(roundAnyRawFNToRecFN_io_covSum),
    .metaAssert(roundAnyRawFNToRecFN_metaAssert)
  );
  assign intAsRawFloat_sign = io_signedIn & io_in[63]; // @[rawFloatFromIN.scala 50:29]
  assign _intAsRawFloat_absIn_T_1 = 64'h0 - io_in; // @[rawFloatFromIN.scala 51:31]
  assign intAsRawFloat_extAbsIn_lo = intAsRawFloat_sign ? _intAsRawFloat_absIn_T_1 : io_in; // @[rawFloatFromIN.scala 51:24]
  assign _intAsRawFloat_extAbsIn_T = {64'h0,intAsRawFloat_extAbsIn_lo}; // @[Cat.scala 30:58]
  assign intAsRawFloat_extAbsIn = _intAsRawFloat_extAbsIn_T[63:0]; // @[rawFloatFromIN.scala 52:56]
  assign _intAsRawFloat_adjustedNormDist_T_64 = intAsRawFloat_extAbsIn[1] ? 6'h3e : 6'h3f; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_65 = intAsRawFloat_extAbsIn[2] ? 6'h3d : _intAsRawFloat_adjustedNormDist_T_64; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_66 = intAsRawFloat_extAbsIn[3] ? 6'h3c : _intAsRawFloat_adjustedNormDist_T_65; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_67 = intAsRawFloat_extAbsIn[4] ? 6'h3b : _intAsRawFloat_adjustedNormDist_T_66; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_68 = intAsRawFloat_extAbsIn[5] ? 6'h3a : _intAsRawFloat_adjustedNormDist_T_67; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_69 = intAsRawFloat_extAbsIn[6] ? 6'h39 : _intAsRawFloat_adjustedNormDist_T_68; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_70 = intAsRawFloat_extAbsIn[7] ? 6'h38 : _intAsRawFloat_adjustedNormDist_T_69; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_71 = intAsRawFloat_extAbsIn[8] ? 6'h37 : _intAsRawFloat_adjustedNormDist_T_70; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_72 = intAsRawFloat_extAbsIn[9] ? 6'h36 : _intAsRawFloat_adjustedNormDist_T_71; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_73 = intAsRawFloat_extAbsIn[10] ? 6'h35 : _intAsRawFloat_adjustedNormDist_T_72; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_74 = intAsRawFloat_extAbsIn[11] ? 6'h34 : _intAsRawFloat_adjustedNormDist_T_73; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_75 = intAsRawFloat_extAbsIn[12] ? 6'h33 : _intAsRawFloat_adjustedNormDist_T_74; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_76 = intAsRawFloat_extAbsIn[13] ? 6'h32 : _intAsRawFloat_adjustedNormDist_T_75; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_77 = intAsRawFloat_extAbsIn[14] ? 6'h31 : _intAsRawFloat_adjustedNormDist_T_76; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_78 = intAsRawFloat_extAbsIn[15] ? 6'h30 : _intAsRawFloat_adjustedNormDist_T_77; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_79 = intAsRawFloat_extAbsIn[16] ? 6'h2f : _intAsRawFloat_adjustedNormDist_T_78; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_80 = intAsRawFloat_extAbsIn[17] ? 6'h2e : _intAsRawFloat_adjustedNormDist_T_79; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_81 = intAsRawFloat_extAbsIn[18] ? 6'h2d : _intAsRawFloat_adjustedNormDist_T_80; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_82 = intAsRawFloat_extAbsIn[19] ? 6'h2c : _intAsRawFloat_adjustedNormDist_T_81; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_83 = intAsRawFloat_extAbsIn[20] ? 6'h2b : _intAsRawFloat_adjustedNormDist_T_82; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_84 = intAsRawFloat_extAbsIn[21] ? 6'h2a : _intAsRawFloat_adjustedNormDist_T_83; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_85 = intAsRawFloat_extAbsIn[22] ? 6'h29 : _intAsRawFloat_adjustedNormDist_T_84; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_86 = intAsRawFloat_extAbsIn[23] ? 6'h28 : _intAsRawFloat_adjustedNormDist_T_85; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_87 = intAsRawFloat_extAbsIn[24] ? 6'h27 : _intAsRawFloat_adjustedNormDist_T_86; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_88 = intAsRawFloat_extAbsIn[25] ? 6'h26 : _intAsRawFloat_adjustedNormDist_T_87; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_89 = intAsRawFloat_extAbsIn[26] ? 6'h25 : _intAsRawFloat_adjustedNormDist_T_88; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_90 = intAsRawFloat_extAbsIn[27] ? 6'h24 : _intAsRawFloat_adjustedNormDist_T_89; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_91 = intAsRawFloat_extAbsIn[28] ? 6'h23 : _intAsRawFloat_adjustedNormDist_T_90; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_92 = intAsRawFloat_extAbsIn[29] ? 6'h22 : _intAsRawFloat_adjustedNormDist_T_91; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_93 = intAsRawFloat_extAbsIn[30] ? 6'h21 : _intAsRawFloat_adjustedNormDist_T_92; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_94 = intAsRawFloat_extAbsIn[31] ? 6'h20 : _intAsRawFloat_adjustedNormDist_T_93; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_95 = intAsRawFloat_extAbsIn[32] ? 6'h1f : _intAsRawFloat_adjustedNormDist_T_94; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_96 = intAsRawFloat_extAbsIn[33] ? 6'h1e : _intAsRawFloat_adjustedNormDist_T_95; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_97 = intAsRawFloat_extAbsIn[34] ? 6'h1d : _intAsRawFloat_adjustedNormDist_T_96; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_98 = intAsRawFloat_extAbsIn[35] ? 6'h1c : _intAsRawFloat_adjustedNormDist_T_97; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_99 = intAsRawFloat_extAbsIn[36] ? 6'h1b : _intAsRawFloat_adjustedNormDist_T_98; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_100 = intAsRawFloat_extAbsIn[37] ? 6'h1a : _intAsRawFloat_adjustedNormDist_T_99; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_101 = intAsRawFloat_extAbsIn[38] ? 6'h19 : _intAsRawFloat_adjustedNormDist_T_100; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_102 = intAsRawFloat_extAbsIn[39] ? 6'h18 : _intAsRawFloat_adjustedNormDist_T_101; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_103 = intAsRawFloat_extAbsIn[40] ? 6'h17 : _intAsRawFloat_adjustedNormDist_T_102; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_104 = intAsRawFloat_extAbsIn[41] ? 6'h16 : _intAsRawFloat_adjustedNormDist_T_103; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_105 = intAsRawFloat_extAbsIn[42] ? 6'h15 : _intAsRawFloat_adjustedNormDist_T_104; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_106 = intAsRawFloat_extAbsIn[43] ? 6'h14 : _intAsRawFloat_adjustedNormDist_T_105; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_107 = intAsRawFloat_extAbsIn[44] ? 6'h13 : _intAsRawFloat_adjustedNormDist_T_106; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_108 = intAsRawFloat_extAbsIn[45] ? 6'h12 : _intAsRawFloat_adjustedNormDist_T_107; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_109 = intAsRawFloat_extAbsIn[46] ? 6'h11 : _intAsRawFloat_adjustedNormDist_T_108; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_110 = intAsRawFloat_extAbsIn[47] ? 6'h10 : _intAsRawFloat_adjustedNormDist_T_109; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_111 = intAsRawFloat_extAbsIn[48] ? 6'hf : _intAsRawFloat_adjustedNormDist_T_110; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_112 = intAsRawFloat_extAbsIn[49] ? 6'he : _intAsRawFloat_adjustedNormDist_T_111; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_113 = intAsRawFloat_extAbsIn[50] ? 6'hd : _intAsRawFloat_adjustedNormDist_T_112; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_114 = intAsRawFloat_extAbsIn[51] ? 6'hc : _intAsRawFloat_adjustedNormDist_T_113; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_115 = intAsRawFloat_extAbsIn[52] ? 6'hb : _intAsRawFloat_adjustedNormDist_T_114; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_116 = intAsRawFloat_extAbsIn[53] ? 6'ha : _intAsRawFloat_adjustedNormDist_T_115; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_117 = intAsRawFloat_extAbsIn[54] ? 6'h9 : _intAsRawFloat_adjustedNormDist_T_116; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_118 = intAsRawFloat_extAbsIn[55] ? 6'h8 : _intAsRawFloat_adjustedNormDist_T_117; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_119 = intAsRawFloat_extAbsIn[56] ? 6'h7 : _intAsRawFloat_adjustedNormDist_T_118; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_120 = intAsRawFloat_extAbsIn[57] ? 6'h6 : _intAsRawFloat_adjustedNormDist_T_119; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_121 = intAsRawFloat_extAbsIn[58] ? 6'h5 : _intAsRawFloat_adjustedNormDist_T_120; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_122 = intAsRawFloat_extAbsIn[59] ? 6'h4 : _intAsRawFloat_adjustedNormDist_T_121; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_123 = intAsRawFloat_extAbsIn[60] ? 6'h3 : _intAsRawFloat_adjustedNormDist_T_122; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_124 = intAsRawFloat_extAbsIn[61] ? 6'h2 : _intAsRawFloat_adjustedNormDist_T_123; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_125 = intAsRawFloat_extAbsIn[62] ? 6'h1 : _intAsRawFloat_adjustedNormDist_T_124; // @[Mux.scala 47:69]
  assign intAsRawFloat_adjustedNormDist = intAsRawFloat_extAbsIn[63] ? 6'h0 : _intAsRawFloat_adjustedNormDist_T_125; // @[Mux.scala 47:69]
  assign _GEN_0 = {{63'd0}, intAsRawFloat_extAbsIn}; // @[rawFloatFromIN.scala 55:22]
  assign _intAsRawFloat_sig_T = _GEN_0 << intAsRawFloat_adjustedNormDist; // @[rawFloatFromIN.scala 55:22]
  assign intAsRawFloat_sig = _intAsRawFloat_sig_T[63:0]; // @[rawFloatFromIN.scala 55:41]
  assign intAsRawFloat_out_sExp_lo = ~intAsRawFloat_adjustedNormDist; // @[rawFloatFromIN.scala 63:39]
  assign _intAsRawFloat_out_sExp_T_1 = {2'h2,intAsRawFloat_out_sExp_lo}; // @[Cat.scala 30:58]
  assign io_out = roundAnyRawFNToRecFN_io_out; // @[INToRecFN.scala 72:23]
  assign io_exceptionFlags = roundAnyRawFNToRecFN_io_exceptionFlags; // @[INToRecFN.scala 73:23]
  assign roundAnyRawFNToRecFN_io_in_isZero = ~intAsRawFloat_sig[63]; // @[INToRecFN.scala 69:44]
  assign roundAnyRawFNToRecFN_io_in_sign = io_signedIn & io_in[63]; // @[INToRecFN.scala 69:44]
  assign roundAnyRawFNToRecFN_io_in_sExp = {1'b0,$signed(_intAsRawFloat_out_sExp_T_1)}; // @[INToRecFN.scala 69:44]
  assign roundAnyRawFNToRecFN_io_in_sig = {{1'd0}, intAsRawFloat_sig}; // @[INToRecFN.scala 69:44]
  assign roundAnyRawFNToRecFN_io_roundingMode = io_roundingMode; // @[INToRecFN.scala 70:44]
  assign INToRecFN_covSum = 30'h0;
  assign roundAnyRawFNToRecFN_sum = INToRecFN_covSum + roundAnyRawFNToRecFN_io_covSum;
  assign io_covSum = roundAnyRawFNToRecFN_sum;
  assign roundAnyRawFNToRecFN_metaAssert_wire = roundAnyRawFNToRecFN_metaAssert;
  assign metaAssert = roundAnyRawFNToRecFN_metaAssert_wire;
endmodule
module INToRecFN_1(
  input         io_signedIn,
  input  [63:0] io_in,
  input  [2:0]  io_roundingMode,
  output [64:0] io_out,
  output [4:0]  io_exceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  roundAnyRawFNToRecFN_io_in_isZero; // @[INToRecFN.scala 59:15]
  wire  roundAnyRawFNToRecFN_io_in_sign; // @[INToRecFN.scala 59:15]
  wire [8:0] roundAnyRawFNToRecFN_io_in_sExp; // @[INToRecFN.scala 59:15]
  wire [64:0] roundAnyRawFNToRecFN_io_in_sig; // @[INToRecFN.scala 59:15]
  wire [2:0] roundAnyRawFNToRecFN_io_roundingMode; // @[INToRecFN.scala 59:15]
  wire [64:0] roundAnyRawFNToRecFN_io_out; // @[INToRecFN.scala 59:15]
  wire [4:0] roundAnyRawFNToRecFN_io_exceptionFlags; // @[INToRecFN.scala 59:15]
  wire [29:0] roundAnyRawFNToRecFN_io_covSum; // @[INToRecFN.scala 59:15]
  wire  roundAnyRawFNToRecFN_metaAssert; // @[INToRecFN.scala 59:15]
  wire  intAsRawFloat_sign; // @[rawFloatFromIN.scala 50:29]
  wire [63:0] _intAsRawFloat_absIn_T_1; // @[rawFloatFromIN.scala 51:31]
  wire [63:0] intAsRawFloat_extAbsIn_lo; // @[rawFloatFromIN.scala 51:24]
  wire [127:0] _intAsRawFloat_extAbsIn_T; // @[Cat.scala 30:58]
  wire [63:0] intAsRawFloat_extAbsIn; // @[rawFloatFromIN.scala 52:56]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_64; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_65; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_66; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_67; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_68; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_69; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_70; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_71; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_72; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_73; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_74; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_75; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_76; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_77; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_78; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_79; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_80; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_81; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_82; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_83; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_84; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_85; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_86; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_87; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_88; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_89; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_90; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_91; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_92; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_93; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_94; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_95; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_96; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_97; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_98; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_99; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_100; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_101; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_102; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_103; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_104; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_105; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_106; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_107; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_108; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_109; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_110; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_111; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_112; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_113; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_114; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_115; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_116; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_117; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_118; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_119; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_120; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_121; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_122; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_123; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_124; // @[Mux.scala 47:69]
  wire [5:0] _intAsRawFloat_adjustedNormDist_T_125; // @[Mux.scala 47:69]
  wire [5:0] intAsRawFloat_adjustedNormDist; // @[Mux.scala 47:69]
  wire [126:0] _GEN_0; // @[rawFloatFromIN.scala 55:22]
  wire [126:0] _intAsRawFloat_sig_T; // @[rawFloatFromIN.scala 55:22]
  wire [63:0] intAsRawFloat_sig; // @[rawFloatFromIN.scala 55:41]
  wire [5:0] intAsRawFloat_out_sExp_lo; // @[rawFloatFromIN.scala 63:39]
  wire [7:0] _intAsRawFloat_out_sExp_T_1; // @[Cat.scala 30:58]
  wire [29:0] INToRecFN_1_covSum;
  wire [29:0] roundAnyRawFNToRecFN_sum;
  wire  roundAnyRawFNToRecFN_metaAssert_wire;
  RoundAnyRawFNToRecFN_2 roundAnyRawFNToRecFN ( // @[INToRecFN.scala 59:15]
    .io_in_isZero(roundAnyRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundAnyRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundAnyRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundAnyRawFNToRecFN_io_in_sig),
    .io_roundingMode(roundAnyRawFNToRecFN_io_roundingMode),
    .io_out(roundAnyRawFNToRecFN_io_out),
    .io_exceptionFlags(roundAnyRawFNToRecFN_io_exceptionFlags),
    .io_covSum(roundAnyRawFNToRecFN_io_covSum),
    .metaAssert(roundAnyRawFNToRecFN_metaAssert)
  );
  assign intAsRawFloat_sign = io_signedIn & io_in[63]; // @[rawFloatFromIN.scala 50:29]
  assign _intAsRawFloat_absIn_T_1 = 64'h0 - io_in; // @[rawFloatFromIN.scala 51:31]
  assign intAsRawFloat_extAbsIn_lo = intAsRawFloat_sign ? _intAsRawFloat_absIn_T_1 : io_in; // @[rawFloatFromIN.scala 51:24]
  assign _intAsRawFloat_extAbsIn_T = {64'h0,intAsRawFloat_extAbsIn_lo}; // @[Cat.scala 30:58]
  assign intAsRawFloat_extAbsIn = _intAsRawFloat_extAbsIn_T[63:0]; // @[rawFloatFromIN.scala 52:56]
  assign _intAsRawFloat_adjustedNormDist_T_64 = intAsRawFloat_extAbsIn[1] ? 6'h3e : 6'h3f; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_65 = intAsRawFloat_extAbsIn[2] ? 6'h3d : _intAsRawFloat_adjustedNormDist_T_64; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_66 = intAsRawFloat_extAbsIn[3] ? 6'h3c : _intAsRawFloat_adjustedNormDist_T_65; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_67 = intAsRawFloat_extAbsIn[4] ? 6'h3b : _intAsRawFloat_adjustedNormDist_T_66; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_68 = intAsRawFloat_extAbsIn[5] ? 6'h3a : _intAsRawFloat_adjustedNormDist_T_67; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_69 = intAsRawFloat_extAbsIn[6] ? 6'h39 : _intAsRawFloat_adjustedNormDist_T_68; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_70 = intAsRawFloat_extAbsIn[7] ? 6'h38 : _intAsRawFloat_adjustedNormDist_T_69; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_71 = intAsRawFloat_extAbsIn[8] ? 6'h37 : _intAsRawFloat_adjustedNormDist_T_70; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_72 = intAsRawFloat_extAbsIn[9] ? 6'h36 : _intAsRawFloat_adjustedNormDist_T_71; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_73 = intAsRawFloat_extAbsIn[10] ? 6'h35 : _intAsRawFloat_adjustedNormDist_T_72; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_74 = intAsRawFloat_extAbsIn[11] ? 6'h34 : _intAsRawFloat_adjustedNormDist_T_73; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_75 = intAsRawFloat_extAbsIn[12] ? 6'h33 : _intAsRawFloat_adjustedNormDist_T_74; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_76 = intAsRawFloat_extAbsIn[13] ? 6'h32 : _intAsRawFloat_adjustedNormDist_T_75; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_77 = intAsRawFloat_extAbsIn[14] ? 6'h31 : _intAsRawFloat_adjustedNormDist_T_76; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_78 = intAsRawFloat_extAbsIn[15] ? 6'h30 : _intAsRawFloat_adjustedNormDist_T_77; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_79 = intAsRawFloat_extAbsIn[16] ? 6'h2f : _intAsRawFloat_adjustedNormDist_T_78; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_80 = intAsRawFloat_extAbsIn[17] ? 6'h2e : _intAsRawFloat_adjustedNormDist_T_79; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_81 = intAsRawFloat_extAbsIn[18] ? 6'h2d : _intAsRawFloat_adjustedNormDist_T_80; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_82 = intAsRawFloat_extAbsIn[19] ? 6'h2c : _intAsRawFloat_adjustedNormDist_T_81; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_83 = intAsRawFloat_extAbsIn[20] ? 6'h2b : _intAsRawFloat_adjustedNormDist_T_82; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_84 = intAsRawFloat_extAbsIn[21] ? 6'h2a : _intAsRawFloat_adjustedNormDist_T_83; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_85 = intAsRawFloat_extAbsIn[22] ? 6'h29 : _intAsRawFloat_adjustedNormDist_T_84; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_86 = intAsRawFloat_extAbsIn[23] ? 6'h28 : _intAsRawFloat_adjustedNormDist_T_85; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_87 = intAsRawFloat_extAbsIn[24] ? 6'h27 : _intAsRawFloat_adjustedNormDist_T_86; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_88 = intAsRawFloat_extAbsIn[25] ? 6'h26 : _intAsRawFloat_adjustedNormDist_T_87; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_89 = intAsRawFloat_extAbsIn[26] ? 6'h25 : _intAsRawFloat_adjustedNormDist_T_88; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_90 = intAsRawFloat_extAbsIn[27] ? 6'h24 : _intAsRawFloat_adjustedNormDist_T_89; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_91 = intAsRawFloat_extAbsIn[28] ? 6'h23 : _intAsRawFloat_adjustedNormDist_T_90; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_92 = intAsRawFloat_extAbsIn[29] ? 6'h22 : _intAsRawFloat_adjustedNormDist_T_91; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_93 = intAsRawFloat_extAbsIn[30] ? 6'h21 : _intAsRawFloat_adjustedNormDist_T_92; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_94 = intAsRawFloat_extAbsIn[31] ? 6'h20 : _intAsRawFloat_adjustedNormDist_T_93; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_95 = intAsRawFloat_extAbsIn[32] ? 6'h1f : _intAsRawFloat_adjustedNormDist_T_94; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_96 = intAsRawFloat_extAbsIn[33] ? 6'h1e : _intAsRawFloat_adjustedNormDist_T_95; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_97 = intAsRawFloat_extAbsIn[34] ? 6'h1d : _intAsRawFloat_adjustedNormDist_T_96; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_98 = intAsRawFloat_extAbsIn[35] ? 6'h1c : _intAsRawFloat_adjustedNormDist_T_97; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_99 = intAsRawFloat_extAbsIn[36] ? 6'h1b : _intAsRawFloat_adjustedNormDist_T_98; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_100 = intAsRawFloat_extAbsIn[37] ? 6'h1a : _intAsRawFloat_adjustedNormDist_T_99; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_101 = intAsRawFloat_extAbsIn[38] ? 6'h19 : _intAsRawFloat_adjustedNormDist_T_100; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_102 = intAsRawFloat_extAbsIn[39] ? 6'h18 : _intAsRawFloat_adjustedNormDist_T_101; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_103 = intAsRawFloat_extAbsIn[40] ? 6'h17 : _intAsRawFloat_adjustedNormDist_T_102; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_104 = intAsRawFloat_extAbsIn[41] ? 6'h16 : _intAsRawFloat_adjustedNormDist_T_103; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_105 = intAsRawFloat_extAbsIn[42] ? 6'h15 : _intAsRawFloat_adjustedNormDist_T_104; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_106 = intAsRawFloat_extAbsIn[43] ? 6'h14 : _intAsRawFloat_adjustedNormDist_T_105; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_107 = intAsRawFloat_extAbsIn[44] ? 6'h13 : _intAsRawFloat_adjustedNormDist_T_106; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_108 = intAsRawFloat_extAbsIn[45] ? 6'h12 : _intAsRawFloat_adjustedNormDist_T_107; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_109 = intAsRawFloat_extAbsIn[46] ? 6'h11 : _intAsRawFloat_adjustedNormDist_T_108; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_110 = intAsRawFloat_extAbsIn[47] ? 6'h10 : _intAsRawFloat_adjustedNormDist_T_109; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_111 = intAsRawFloat_extAbsIn[48] ? 6'hf : _intAsRawFloat_adjustedNormDist_T_110; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_112 = intAsRawFloat_extAbsIn[49] ? 6'he : _intAsRawFloat_adjustedNormDist_T_111; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_113 = intAsRawFloat_extAbsIn[50] ? 6'hd : _intAsRawFloat_adjustedNormDist_T_112; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_114 = intAsRawFloat_extAbsIn[51] ? 6'hc : _intAsRawFloat_adjustedNormDist_T_113; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_115 = intAsRawFloat_extAbsIn[52] ? 6'hb : _intAsRawFloat_adjustedNormDist_T_114; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_116 = intAsRawFloat_extAbsIn[53] ? 6'ha : _intAsRawFloat_adjustedNormDist_T_115; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_117 = intAsRawFloat_extAbsIn[54] ? 6'h9 : _intAsRawFloat_adjustedNormDist_T_116; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_118 = intAsRawFloat_extAbsIn[55] ? 6'h8 : _intAsRawFloat_adjustedNormDist_T_117; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_119 = intAsRawFloat_extAbsIn[56] ? 6'h7 : _intAsRawFloat_adjustedNormDist_T_118; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_120 = intAsRawFloat_extAbsIn[57] ? 6'h6 : _intAsRawFloat_adjustedNormDist_T_119; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_121 = intAsRawFloat_extAbsIn[58] ? 6'h5 : _intAsRawFloat_adjustedNormDist_T_120; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_122 = intAsRawFloat_extAbsIn[59] ? 6'h4 : _intAsRawFloat_adjustedNormDist_T_121; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_123 = intAsRawFloat_extAbsIn[60] ? 6'h3 : _intAsRawFloat_adjustedNormDist_T_122; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_124 = intAsRawFloat_extAbsIn[61] ? 6'h2 : _intAsRawFloat_adjustedNormDist_T_123; // @[Mux.scala 47:69]
  assign _intAsRawFloat_adjustedNormDist_T_125 = intAsRawFloat_extAbsIn[62] ? 6'h1 : _intAsRawFloat_adjustedNormDist_T_124; // @[Mux.scala 47:69]
  assign intAsRawFloat_adjustedNormDist = intAsRawFloat_extAbsIn[63] ? 6'h0 : _intAsRawFloat_adjustedNormDist_T_125; // @[Mux.scala 47:69]
  assign _GEN_0 = {{63'd0}, intAsRawFloat_extAbsIn}; // @[rawFloatFromIN.scala 55:22]
  assign _intAsRawFloat_sig_T = _GEN_0 << intAsRawFloat_adjustedNormDist; // @[rawFloatFromIN.scala 55:22]
  assign intAsRawFloat_sig = _intAsRawFloat_sig_T[63:0]; // @[rawFloatFromIN.scala 55:41]
  assign intAsRawFloat_out_sExp_lo = ~intAsRawFloat_adjustedNormDist; // @[rawFloatFromIN.scala 63:39]
  assign _intAsRawFloat_out_sExp_T_1 = {2'h2,intAsRawFloat_out_sExp_lo}; // @[Cat.scala 30:58]
  assign io_out = roundAnyRawFNToRecFN_io_out; // @[INToRecFN.scala 72:23]
  assign io_exceptionFlags = roundAnyRawFNToRecFN_io_exceptionFlags; // @[INToRecFN.scala 73:23]
  assign roundAnyRawFNToRecFN_io_in_isZero = ~intAsRawFloat_sig[63]; // @[INToRecFN.scala 69:44]
  assign roundAnyRawFNToRecFN_io_in_sign = io_signedIn & io_in[63]; // @[INToRecFN.scala 69:44]
  assign roundAnyRawFNToRecFN_io_in_sExp = {1'b0,$signed(_intAsRawFloat_out_sExp_T_1)}; // @[INToRecFN.scala 69:44]
  assign roundAnyRawFNToRecFN_io_in_sig = {{1'd0}, intAsRawFloat_sig}; // @[INToRecFN.scala 69:44]
  assign roundAnyRawFNToRecFN_io_roundingMode = io_roundingMode; // @[INToRecFN.scala 70:44]
  assign INToRecFN_1_covSum = 30'h0;
  assign roundAnyRawFNToRecFN_sum = INToRecFN_1_covSum + roundAnyRawFNToRecFN_io_covSum;
  assign io_covSum = roundAnyRawFNToRecFN_sum;
  assign roundAnyRawFNToRecFN_metaAssert_wire = roundAnyRawFNToRecFN_metaAssert;
  assign metaAssert = roundAnyRawFNToRecFN_metaAssert_wire;
endmodule
module RecFNToRecFN(
  input  [64:0] io_in,
  input  [2:0]  io_roundingMode,
  output [32:0] io_out,
  output [4:0]  io_exceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  roundAnyRawFNToRecFN_io_invalidExc; // @[RecFNToRecFN.scala 72:19]
  wire  roundAnyRawFNToRecFN_io_in_isNaN; // @[RecFNToRecFN.scala 72:19]
  wire  roundAnyRawFNToRecFN_io_in_isInf; // @[RecFNToRecFN.scala 72:19]
  wire  roundAnyRawFNToRecFN_io_in_isZero; // @[RecFNToRecFN.scala 72:19]
  wire  roundAnyRawFNToRecFN_io_in_sign; // @[RecFNToRecFN.scala 72:19]
  wire [12:0] roundAnyRawFNToRecFN_io_in_sExp; // @[RecFNToRecFN.scala 72:19]
  wire [53:0] roundAnyRawFNToRecFN_io_in_sig; // @[RecFNToRecFN.scala 72:19]
  wire [2:0] roundAnyRawFNToRecFN_io_roundingMode; // @[RecFNToRecFN.scala 72:19]
  wire [32:0] roundAnyRawFNToRecFN_io_out; // @[RecFNToRecFN.scala 72:19]
  wire [4:0] roundAnyRawFNToRecFN_io_exceptionFlags; // @[RecFNToRecFN.scala 72:19]
  wire [29:0] roundAnyRawFNToRecFN_io_covSum; // @[RecFNToRecFN.scala 72:19]
  wire  roundAnyRawFNToRecFN_metaAssert; // @[RecFNToRecFN.scala 72:19]
  wire [11:0] rawIn_exp; // @[rawFloatFromRecFN.scala 50:21]
  wire  rawIn_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  rawIn_isSpecial; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawIn__isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawIn_out_sig_hi_lo; // @[rawFloatFromRecFN.scala 60:39]
  wire [51:0] rawIn_out_sig_lo; // @[rawFloatFromRecFN.scala 60:51]
  wire [1:0] rawIn_out_sig_hi; // @[Cat.scala 30:58]
  wire [53:0] rawIn__sig; // @[Cat.scala 30:58]
  wire [29:0] RecFNToRecFN_covSum;
  wire [29:0] roundAnyRawFNToRecFN_sum;
  wire  roundAnyRawFNToRecFN_metaAssert_wire;
  RoundAnyRawFNToRecFN_3 roundAnyRawFNToRecFN ( // @[RecFNToRecFN.scala 72:19]
    .io_invalidExc(roundAnyRawFNToRecFN_io_invalidExc),
    .io_in_isNaN(roundAnyRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundAnyRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundAnyRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundAnyRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundAnyRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundAnyRawFNToRecFN_io_in_sig),
    .io_roundingMode(roundAnyRawFNToRecFN_io_roundingMode),
    .io_out(roundAnyRawFNToRecFN_io_out),
    .io_exceptionFlags(roundAnyRawFNToRecFN_io_exceptionFlags),
    .io_covSum(roundAnyRawFNToRecFN_io_covSum),
    .metaAssert(roundAnyRawFNToRecFN_metaAssert)
  );
  assign rawIn_exp = io_in[63:52]; // @[rawFloatFromRecFN.scala 50:21]
  assign rawIn_isZero = rawIn_exp[11:9] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign rawIn_isSpecial = rawIn_exp[11:10] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawIn__isNaN = rawIn_isSpecial & rawIn_exp[9]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawIn_out_sig_hi_lo = ~rawIn_isZero; // @[rawFloatFromRecFN.scala 60:39]
  assign rawIn_out_sig_lo = io_in[51:0]; // @[rawFloatFromRecFN.scala 60:51]
  assign rawIn_out_sig_hi = {1'h0,rawIn_out_sig_hi_lo}; // @[Cat.scala 30:58]
  assign rawIn__sig = {1'h0,rawIn_out_sig_hi_lo,rawIn_out_sig_lo}; // @[Cat.scala 30:58]
  assign io_out = roundAnyRawFNToRecFN_io_out; // @[RecFNToRecFN.scala 85:27]
  assign io_exceptionFlags = roundAnyRawFNToRecFN_io_exceptionFlags; // @[RecFNToRecFN.scala 86:27]
  assign roundAnyRawFNToRecFN_io_invalidExc = rawIn__isNaN & ~rawIn__sig[51]; // @[RecFNToRecFN.scala 80:48]
  assign roundAnyRawFNToRecFN_io_in_isNaN = rawIn_isSpecial & rawIn_exp[9]; // @[RecFNToRecFN.scala 82:48]
  assign roundAnyRawFNToRecFN_io_in_isInf = rawIn_isSpecial & ~rawIn_exp[9]; // @[RecFNToRecFN.scala 82:48]
  assign roundAnyRawFNToRecFN_io_in_isZero = rawIn_exp[11:9] == 3'h0; // @[RecFNToRecFN.scala 82:48]
  assign roundAnyRawFNToRecFN_io_in_sign = io_in[64]; // @[RecFNToRecFN.scala 82:48]
  assign roundAnyRawFNToRecFN_io_in_sExp = {1'b0,$signed(rawIn_exp)}; // @[RecFNToRecFN.scala 82:48]
  assign roundAnyRawFNToRecFN_io_in_sig = {rawIn_out_sig_hi,rawIn_out_sig_lo}; // @[RecFNToRecFN.scala 82:48]
  assign roundAnyRawFNToRecFN_io_roundingMode = io_roundingMode; // @[RecFNToRecFN.scala 83:48]
  assign RecFNToRecFN_covSum = 30'h0;
  assign roundAnyRawFNToRecFN_sum = RecFNToRecFN_covSum + roundAnyRawFNToRecFN_io_covSum;
  assign io_covSum = roundAnyRawFNToRecFN_sum;
  assign roundAnyRawFNToRecFN_metaAssert_wire = roundAnyRawFNToRecFN_metaAssert;
  assign metaAssert = roundAnyRawFNToRecFN_metaAssert_wire;
endmodule
module MulAddRecFNPipe_1(
  input         clock,
  input         reset,
  input         io_validin,
  input  [1:0]  io_op,
  input  [64:0] io_a,
  input  [64:0] io_b,
  input  [64:0] io_c,
  input  [2:0]  io_roundingMode,
  output [64:0] io_out,
  output [4:0]  io_exceptionFlags,
  output        io_validout,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  wire [1:0] mulAddRecFNToRaw_preMul_io_op; // @[FPU.scala 648:41]
  wire [64:0] mulAddRecFNToRaw_preMul_io_a; // @[FPU.scala 648:41]
  wire [64:0] mulAddRecFNToRaw_preMul_io_b; // @[FPU.scala 648:41]
  wire [64:0] mulAddRecFNToRaw_preMul_io_c; // @[FPU.scala 648:41]
  wire [52:0] mulAddRecFNToRaw_preMul_io_mulAddA; // @[FPU.scala 648:41]
  wire [52:0] mulAddRecFNToRaw_preMul_io_mulAddB; // @[FPU.scala 648:41]
  wire [105:0] mulAddRecFNToRaw_preMul_io_mulAddC; // @[FPU.scala 648:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny; // @[FPU.scala 648:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB; // @[FPU.scala 648:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfA; // @[FPU.scala 648:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA; // @[FPU.scala 648:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfB; // @[FPU.scala 648:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB; // @[FPU.scala 648:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_signProd; // @[FPU.scala 648:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC; // @[FPU.scala 648:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfC; // @[FPU.scala 648:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC; // @[FPU.scala 648:41]
  wire [12:0] mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum; // @[FPU.scala 648:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags; // @[FPU.scala 648:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant; // @[FPU.scala 648:41]
  wire [5:0] mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist; // @[FPU.scala 648:41]
  wire [54:0] mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC; // @[FPU.scala 648:41]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC; // @[FPU.scala 648:41]
  wire [29:0] mulAddRecFNToRaw_preMul_io_covSum; // @[FPU.scala 648:41]
  wire  mulAddRecFNToRaw_preMul_metaAssert; // @[FPU.scala 648:41]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny; // @[FPU.scala 649:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB; // @[FPU.scala 649:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA; // @[FPU.scala 649:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA; // @[FPU.scala 649:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB; // @[FPU.scala 649:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB; // @[FPU.scala 649:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_signProd; // @[FPU.scala 649:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC; // @[FPU.scala 649:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC; // @[FPU.scala 649:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC; // @[FPU.scala 649:42]
  wire [12:0] mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum; // @[FPU.scala 649:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags; // @[FPU.scala 649:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant; // @[FPU.scala 649:42]
  wire [5:0] mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist; // @[FPU.scala 649:42]
  wire [54:0] mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC; // @[FPU.scala 649:42]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC; // @[FPU.scala 649:42]
  wire [106:0] mulAddRecFNToRaw_postMul_io_mulAddResult; // @[FPU.scala 649:42]
  wire [2:0] mulAddRecFNToRaw_postMul_io_roundingMode; // @[FPU.scala 649:42]
  wire  mulAddRecFNToRaw_postMul_io_invalidExc; // @[FPU.scala 649:42]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isNaN; // @[FPU.scala 649:42]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isInf; // @[FPU.scala 649:42]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isZero; // @[FPU.scala 649:42]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_sign; // @[FPU.scala 649:42]
  wire [12:0] mulAddRecFNToRaw_postMul_io_rawOut_sExp; // @[FPU.scala 649:42]
  wire [55:0] mulAddRecFNToRaw_postMul_io_rawOut_sig; // @[FPU.scala 649:42]
  wire [29:0] mulAddRecFNToRaw_postMul_io_covSum; // @[FPU.scala 649:42]
  wire  mulAddRecFNToRaw_postMul_metaAssert; // @[FPU.scala 649:42]
  wire  roundRawFNToRecFN_io_invalidExc; // @[FPU.scala 676:35]
  wire  roundRawFNToRecFN_io_infiniteExc; // @[FPU.scala 676:35]
  wire  roundRawFNToRecFN_io_in_isNaN; // @[FPU.scala 676:35]
  wire  roundRawFNToRecFN_io_in_isInf; // @[FPU.scala 676:35]
  wire  roundRawFNToRecFN_io_in_isZero; // @[FPU.scala 676:35]
  wire  roundRawFNToRecFN_io_in_sign; // @[FPU.scala 676:35]
  wire [12:0] roundRawFNToRecFN_io_in_sExp; // @[FPU.scala 676:35]
  wire [55:0] roundRawFNToRecFN_io_in_sig; // @[FPU.scala 676:35]
  wire [2:0] roundRawFNToRecFN_io_roundingMode; // @[FPU.scala 676:35]
  wire  roundRawFNToRecFN_io_detectTininess; // @[FPU.scala 676:35]
  wire [64:0] roundRawFNToRecFN_io_out; // @[FPU.scala 676:35]
  wire [4:0] roundRawFNToRecFN_io_exceptionFlags; // @[FPU.scala 676:35]
  wire [29:0] roundRawFNToRecFN_io_covSum; // @[FPU.scala 676:35]
  wire  roundRawFNToRecFN_metaAssert; // @[FPU.scala 676:35]
  wire [105:0] _mulAddResult_T; // @[FPU.scala 657:45]
  wire [106:0] mulAddResult; // @[FPU.scala 658:50]
  reg  mulAddRecFNToRaw_postMul_io_fromPreMul_b_isSigNaNAny; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  reg  mulAddRecFNToRaw_postMul_io_fromPreMul_b_isNaNAOrB; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  reg  mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfA; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg  mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroA; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg  mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfB; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg  mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroB; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg  mulAddRecFNToRaw_postMul_io_fromPreMul_b_signProd; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg  mulAddRecFNToRaw_postMul_io_fromPreMul_b_isNaNC; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7;
  reg  mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfC; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8;
  reg  mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroC; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  reg [12:0] mulAddRecFNToRaw_postMul_io_fromPreMul_b_sExpSum; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10;
  reg  mulAddRecFNToRaw_postMul_io_fromPreMul_b_doSubMags; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11;
  reg  mulAddRecFNToRaw_postMul_io_fromPreMul_b_CIsDominant; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12;
  reg [5:0] mulAddRecFNToRaw_postMul_io_fromPreMul_b_CDom_CAlignDist; // @[Reg.scala 15:16]
  reg [31:0] _RAND_13;
  reg [54:0] mulAddRecFNToRaw_postMul_io_fromPreMul_b_highAlignedSigC; // @[Reg.scala 15:16]
  reg [63:0] _RAND_14;
  reg  mulAddRecFNToRaw_postMul_io_fromPreMul_b_bit0AlignedSigC; // @[Reg.scala 15:16]
  reg [31:0] _RAND_15;
  reg [106:0] mulAddRecFNToRaw_postMul_io_mulAddResult_b; // @[Reg.scala 15:16]
  reg [127:0] _RAND_16;
  reg [2:0] mulAddRecFNToRaw_postMul_io_roundingMode_b; // @[Reg.scala 15:16]
  reg [31:0] _RAND_17;
  reg [2:0] roundingMode_stage0_b; // @[Reg.scala 15:16]
  reg [31:0] _RAND_18;
  reg  detectTininess_stage0_b; // @[Reg.scala 15:16]
  reg [31:0] _RAND_19;
  reg  valid_stage0_v; // @[Valid.scala 117:22]
  reg [31:0] _RAND_20;
  reg  roundRawFNToRecFN_io_invalidExc_b; // @[Reg.scala 15:16]
  reg [31:0] _RAND_21;
  reg  roundRawFNToRecFN_io_in_b_isNaN; // @[Reg.scala 15:16]
  reg [31:0] _RAND_22;
  reg  roundRawFNToRecFN_io_in_b_isInf; // @[Reg.scala 15:16]
  reg [31:0] _RAND_23;
  reg  roundRawFNToRecFN_io_in_b_isZero; // @[Reg.scala 15:16]
  reg [31:0] _RAND_24;
  reg  roundRawFNToRecFN_io_in_b_sign; // @[Reg.scala 15:16]
  reg [31:0] _RAND_25;
  reg [12:0] roundRawFNToRecFN_io_in_b_sExp; // @[Reg.scala 15:16]
  reg [31:0] _RAND_26;
  reg [55:0] roundRawFNToRecFN_io_in_b_sig; // @[Reg.scala 15:16]
  reg [63:0] _RAND_27;
  reg [2:0] roundRawFNToRecFN_io_roundingMode_b; // @[Reg.scala 15:16]
  reg [31:0] _RAND_28;
  reg  roundRawFNToRecFN_io_detectTininess_b; // @[Reg.scala 15:16]
  reg [31:0] _RAND_29;
  reg  io_validout_v; // @[Valid.scala 117:22]
  reg [31:0] _RAND_30;
  reg  MulAddRecFNPipe_1_state; // @[Register tracking MulAddRecFNPipe_1 state]
  reg [31:0] _RAND_31;
  reg  MulAddRecFNPipe_1_cov [0:1]; // @[Coverage map for MulAddRecFNPipe_1]
  reg [31:0] _RAND_32;
  wire  MulAddRecFNPipe_1_cov_read_data; // @[Coverage map for MulAddRecFNPipe_1]
  wire  MulAddRecFNPipe_1_cov_read_addr; // @[Coverage map for MulAddRecFNPipe_1]
  wire  MulAddRecFNPipe_1_cov_write_data; // @[Coverage map for MulAddRecFNPipe_1]
  wire  MulAddRecFNPipe_1_cov_write_addr; // @[Coverage map for MulAddRecFNPipe_1]
  wire  MulAddRecFNPipe_1_cov_write_mask; // @[Coverage map for MulAddRecFNPipe_1]
  wire  MulAddRecFNPipe_1_cov_write_en; // @[Coverage map for MulAddRecFNPipe_1]
  reg [29:0] MulAddRecFNPipe_1_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_33;
  wire  valid_stage0_v_shl;
  wire  valid_stage0_v_pad;
  wire [29:0] mulAddRecFNToRaw_preMul_sum;
  wire [29:0] mulAddRecFNToRaw_postMul_sum;
  wire [29:0] roundRawFNToRecFN_sum;
  wire  mulAddRecFNToRaw_preMul_metaAssert_wire;
  wire  mulAddRecFNToRaw_postMul_metaAssert_wire;
  wire  roundRawFNToRecFN_metaAssert_wire;
  wire  MulAddRecFNPipe_1_or2;
  wire  MulAddRecFNPipe_1_or0;
  reg  MulAddRecFNPipe_1_metaAssert;
  reg [31:0] _RAND_34;
  MulAddRecFNToRaw_preMul_1 mulAddRecFNToRaw_preMul ( // @[FPU.scala 648:41]
    .io_op(mulAddRecFNToRaw_preMul_io_op),
    .io_a(mulAddRecFNToRaw_preMul_io_a),
    .io_b(mulAddRecFNToRaw_preMul_io_b),
    .io_c(mulAddRecFNToRaw_preMul_io_c),
    .io_mulAddA(mulAddRecFNToRaw_preMul_io_mulAddA),
    .io_mulAddB(mulAddRecFNToRaw_preMul_io_mulAddB),
    .io_mulAddC(mulAddRecFNToRaw_preMul_io_mulAddC),
    .io_toPostMul_isSigNaNAny(mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny),
    .io_toPostMul_isNaNAOrB(mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB),
    .io_toPostMul_isInfA(mulAddRecFNToRaw_preMul_io_toPostMul_isInfA),
    .io_toPostMul_isZeroA(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA),
    .io_toPostMul_isInfB(mulAddRecFNToRaw_preMul_io_toPostMul_isInfB),
    .io_toPostMul_isZeroB(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB),
    .io_toPostMul_signProd(mulAddRecFNToRaw_preMul_io_toPostMul_signProd),
    .io_toPostMul_isNaNC(mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC),
    .io_toPostMul_isInfC(mulAddRecFNToRaw_preMul_io_toPostMul_isInfC),
    .io_toPostMul_isZeroC(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC),
    .io_toPostMul_sExpSum(mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum),
    .io_toPostMul_doSubMags(mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags),
    .io_toPostMul_CIsDominant(mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant),
    .io_toPostMul_CDom_CAlignDist(mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist),
    .io_toPostMul_highAlignedSigC(mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC),
    .io_toPostMul_bit0AlignedSigC(mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC),
    .io_covSum(mulAddRecFNToRaw_preMul_io_covSum),
    .metaAssert(mulAddRecFNToRaw_preMul_metaAssert)
  );
  MulAddRecFNToRaw_postMul_1 mulAddRecFNToRaw_postMul ( // @[FPU.scala 649:42]
    .io_fromPreMul_isSigNaNAny(mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny),
    .io_fromPreMul_isNaNAOrB(mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB),
    .io_fromPreMul_isInfA(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA),
    .io_fromPreMul_isZeroA(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA),
    .io_fromPreMul_isInfB(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB),
    .io_fromPreMul_isZeroB(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB),
    .io_fromPreMul_signProd(mulAddRecFNToRaw_postMul_io_fromPreMul_signProd),
    .io_fromPreMul_isNaNC(mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC),
    .io_fromPreMul_isInfC(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC),
    .io_fromPreMul_isZeroC(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC),
    .io_fromPreMul_sExpSum(mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum),
    .io_fromPreMul_doSubMags(mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags),
    .io_fromPreMul_CIsDominant(mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant),
    .io_fromPreMul_CDom_CAlignDist(mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist),
    .io_fromPreMul_highAlignedSigC(mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC),
    .io_fromPreMul_bit0AlignedSigC(mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC),
    .io_mulAddResult(mulAddRecFNToRaw_postMul_io_mulAddResult),
    .io_roundingMode(mulAddRecFNToRaw_postMul_io_roundingMode),
    .io_invalidExc(mulAddRecFNToRaw_postMul_io_invalidExc),
    .io_rawOut_isNaN(mulAddRecFNToRaw_postMul_io_rawOut_isNaN),
    .io_rawOut_isInf(mulAddRecFNToRaw_postMul_io_rawOut_isInf),
    .io_rawOut_isZero(mulAddRecFNToRaw_postMul_io_rawOut_isZero),
    .io_rawOut_sign(mulAddRecFNToRaw_postMul_io_rawOut_sign),
    .io_rawOut_sExp(mulAddRecFNToRaw_postMul_io_rawOut_sExp),
    .io_rawOut_sig(mulAddRecFNToRaw_postMul_io_rawOut_sig),
    .io_covSum(mulAddRecFNToRaw_postMul_io_covSum),
    .metaAssert(mulAddRecFNToRaw_postMul_metaAssert)
  );
  RoundRawFNToRecFN_3 roundRawFNToRecFN ( // @[FPU.scala 676:35]
    .io_invalidExc(roundRawFNToRecFN_io_invalidExc),
    .io_infiniteExc(roundRawFNToRecFN_io_infiniteExc),
    .io_in_isNaN(roundRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundRawFNToRecFN_io_in_sig),
    .io_roundingMode(roundRawFNToRecFN_io_roundingMode),
    .io_detectTininess(roundRawFNToRecFN_io_detectTininess),
    .io_out(roundRawFNToRecFN_io_out),
    .io_exceptionFlags(roundRawFNToRecFN_io_exceptionFlags),
    .io_covSum(roundRawFNToRecFN_io_covSum),
    .metaAssert(roundRawFNToRecFN_metaAssert)
  );
  assign _mulAddResult_T = mulAddRecFNToRaw_preMul_io_mulAddA * mulAddRecFNToRaw_preMul_io_mulAddB; // @[FPU.scala 657:45]
  assign mulAddResult = _mulAddResult_T + mulAddRecFNToRaw_preMul_io_mulAddC; // @[FPU.scala 658:50]
  assign io_out = roundRawFNToRecFN_io_out; // @[FPU.scala 687:23]
  assign io_exceptionFlags = roundRawFNToRecFN_io_exceptionFlags; // @[FPU.scala 688:23]
  assign io_validout = io_validout_v; // @[FPU.scala 683:45]
  assign mulAddRecFNToRaw_preMul_io_op = io_op; // @[FPU.scala 651:35]
  assign mulAddRecFNToRaw_preMul_io_a = io_a; // @[FPU.scala 652:35]
  assign mulAddRecFNToRaw_preMul_io_b = io_b; // @[FPU.scala 653:35]
  assign mulAddRecFNToRaw_preMul_io_c = io_c; // @[FPU.scala 654:35]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny = mulAddRecFNToRaw_postMul_io_fromPreMul_b_isSigNaNAny; // @[FPU.scala 666:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB = mulAddRecFNToRaw_postMul_io_fromPreMul_b_isNaNAOrB; // @[FPU.scala 666:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA = mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfA; // @[FPU.scala 666:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA = mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroA; // @[FPU.scala 666:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB = mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfB; // @[FPU.scala 666:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB = mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroB; // @[FPU.scala 666:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_signProd = mulAddRecFNToRaw_postMul_io_fromPreMul_b_signProd; // @[FPU.scala 666:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC = mulAddRecFNToRaw_postMul_io_fromPreMul_b_isNaNC; // @[FPU.scala 666:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC = mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfC; // @[FPU.scala 666:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC = mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroC; // @[FPU.scala 666:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum = mulAddRecFNToRaw_postMul_io_fromPreMul_b_sExpSum; // @[FPU.scala 666:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags = mulAddRecFNToRaw_postMul_io_fromPreMul_b_doSubMags; // @[FPU.scala 666:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant = mulAddRecFNToRaw_postMul_io_fromPreMul_b_CIsDominant; // @[FPU.scala 666:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist = mulAddRecFNToRaw_postMul_io_fromPreMul_b_CDom_CAlignDist; // @[FPU.scala 666:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC = mulAddRecFNToRaw_postMul_io_fromPreMul_b_highAlignedSigC; // @[FPU.scala 666:46]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC = mulAddRecFNToRaw_postMul_io_fromPreMul_b_bit0AlignedSigC; // @[FPU.scala 666:46]
  assign mulAddRecFNToRaw_postMul_io_mulAddResult = mulAddRecFNToRaw_postMul_io_mulAddResult_b; // @[FPU.scala 667:46]
  assign mulAddRecFNToRaw_postMul_io_roundingMode = mulAddRecFNToRaw_postMul_io_roundingMode_b; // @[FPU.scala 668:46]
  assign roundRawFNToRecFN_io_invalidExc = roundRawFNToRecFN_io_invalidExc_b; // @[FPU.scala 679:45]
  assign roundRawFNToRecFN_io_infiniteExc = 1'h0; // @[FPU.scala 685:38]
  assign roundRawFNToRecFN_io_in_isNaN = roundRawFNToRecFN_io_in_b_isNaN; // @[FPU.scala 680:45]
  assign roundRawFNToRecFN_io_in_isInf = roundRawFNToRecFN_io_in_b_isInf; // @[FPU.scala 680:45]
  assign roundRawFNToRecFN_io_in_isZero = roundRawFNToRecFN_io_in_b_isZero; // @[FPU.scala 680:45]
  assign roundRawFNToRecFN_io_in_sign = roundRawFNToRecFN_io_in_b_sign; // @[FPU.scala 680:45]
  assign roundRawFNToRecFN_io_in_sExp = roundRawFNToRecFN_io_in_b_sExp; // @[FPU.scala 680:45]
  assign roundRawFNToRecFN_io_in_sig = roundRawFNToRecFN_io_in_b_sig; // @[FPU.scala 680:45]
  assign roundRawFNToRecFN_io_roundingMode = roundRawFNToRecFN_io_roundingMode_b; // @[FPU.scala 681:45]
  assign roundRawFNToRecFN_io_detectTininess = roundRawFNToRecFN_io_detectTininess_b; // @[FPU.scala 682:45]
  assign MulAddRecFNPipe_1_cov_read_addr = MulAddRecFNPipe_1_state;
  assign MulAddRecFNPipe_1_cov_read_data = MulAddRecFNPipe_1_cov[MulAddRecFNPipe_1_cov_read_addr]; // @[Coverage map for MulAddRecFNPipe_1]
  assign MulAddRecFNPipe_1_cov_write_data = 1'h1;
  assign MulAddRecFNPipe_1_cov_write_addr = MulAddRecFNPipe_1_state;
  assign MulAddRecFNPipe_1_cov_write_mask = 1'h1;
  assign MulAddRecFNPipe_1_cov_write_en = 1'h1;
  assign valid_stage0_v_shl = valid_stage0_v;
  assign valid_stage0_v_pad = valid_stage0_v_shl;
  assign mulAddRecFNToRaw_preMul_sum = MulAddRecFNPipe_1_covSum + mulAddRecFNToRaw_preMul_io_covSum;
  assign mulAddRecFNToRaw_postMul_sum = mulAddRecFNToRaw_preMul_sum + mulAddRecFNToRaw_postMul_io_covSum;
  assign roundRawFNToRecFN_sum = mulAddRecFNToRaw_postMul_sum + roundRawFNToRecFN_io_covSum;
  assign io_covSum = roundRawFNToRecFN_sum;
  assign mulAddRecFNToRaw_preMul_metaAssert_wire = mulAddRecFNToRaw_preMul_metaAssert;
  assign mulAddRecFNToRaw_postMul_metaAssert_wire = mulAddRecFNToRaw_postMul_metaAssert;
  assign roundRawFNToRecFN_metaAssert_wire = roundRawFNToRecFN_metaAssert;
  assign MulAddRecFNPipe_1_or2 = mulAddRecFNToRaw_postMul_metaAssert_wire | roundRawFNToRecFN_metaAssert_wire;
  assign MulAddRecFNPipe_1_or0 = mulAddRecFNToRaw_preMul_metaAssert_wire | MulAddRecFNPipe_1_or2;
  assign metaAssert = MulAddRecFNPipe_1_metaAssert;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mulAddRecFNToRaw_postMul_io_fromPreMul_b_isSigNaNAny = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mulAddRecFNToRaw_postMul_io_fromPreMul_b_isNaNAOrB = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfA = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroA = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfB = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroB = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  mulAddRecFNToRaw_postMul_io_fromPreMul_b_signProd = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  mulAddRecFNToRaw_postMul_io_fromPreMul_b_isNaNC = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfC = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroC = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  mulAddRecFNToRaw_postMul_io_fromPreMul_b_sExpSum = _RAND_10[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  mulAddRecFNToRaw_postMul_io_fromPreMul_b_doSubMags = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  mulAddRecFNToRaw_postMul_io_fromPreMul_b_CIsDominant = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  mulAddRecFNToRaw_postMul_io_fromPreMul_b_CDom_CAlignDist = _RAND_13[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {2{`RANDOM}};
  mulAddRecFNToRaw_postMul_io_fromPreMul_b_highAlignedSigC = _RAND_14[54:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  mulAddRecFNToRaw_postMul_io_fromPreMul_b_bit0AlignedSigC = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {4{`RANDOM}};
  mulAddRecFNToRaw_postMul_io_mulAddResult_b = _RAND_16[106:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  mulAddRecFNToRaw_postMul_io_roundingMode_b = _RAND_17[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  roundingMode_stage0_b = _RAND_18[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  detectTininess_stage0_b = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  valid_stage0_v = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  roundRawFNToRecFN_io_invalidExc_b = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  roundRawFNToRecFN_io_in_b_isNaN = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  roundRawFNToRecFN_io_in_b_isInf = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  roundRawFNToRecFN_io_in_b_isZero = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  roundRawFNToRecFN_io_in_b_sign = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  roundRawFNToRecFN_io_in_b_sExp = _RAND_26[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {2{`RANDOM}};
  roundRawFNToRecFN_io_in_b_sig = _RAND_27[55:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  roundRawFNToRecFN_io_roundingMode_b = _RAND_28[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  roundRawFNToRecFN_io_detectTininess_b = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  io_validout_v = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  MulAddRecFNPipe_1_state = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    MulAddRecFNPipe_1_cov[initvar] = _RAND_32[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  MulAddRecFNPipe_1_covSum = _RAND_33[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  MulAddRecFNPipe_1_metaAssert = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_isSigNaNAny <= 1'h0;
    end else if (io_validin) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_isSigNaNAny <= mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny;
    end
    if (metaReset) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_isNaNAOrB <= 1'h0;
    end else if (io_validin) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_isNaNAOrB <= mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB;
    end
    if (metaReset) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfA <= 1'h0;
    end else if (io_validin) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfA <= mulAddRecFNToRaw_preMul_io_toPostMul_isInfA;
    end
    if (metaReset) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroA <= 1'h0;
    end else if (io_validin) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroA <= mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA;
    end
    if (metaReset) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfB <= 1'h0;
    end else if (io_validin) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfB <= mulAddRecFNToRaw_preMul_io_toPostMul_isInfB;
    end
    if (metaReset) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroB <= 1'h0;
    end else if (io_validin) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroB <= mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB;
    end
    if (metaReset) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_signProd <= 1'h0;
    end else if (io_validin) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_signProd <= mulAddRecFNToRaw_preMul_io_toPostMul_signProd;
    end
    if (metaReset) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_isNaNC <= 1'h0;
    end else if (io_validin) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_isNaNC <= mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC;
    end
    if (metaReset) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfC <= 1'h0;
    end else if (io_validin) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfC <= mulAddRecFNToRaw_preMul_io_toPostMul_isInfC;
    end
    if (metaReset) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroC <= 1'h0;
    end else if (io_validin) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroC <= mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC;
    end
    if (metaReset) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_sExpSum <= 13'h0;
    end else if (io_validin) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_sExpSum <= mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum;
    end
    if (metaReset) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_doSubMags <= 1'h0;
    end else if (io_validin) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_doSubMags <= mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags;
    end
    if (metaReset) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_CIsDominant <= 1'h0;
    end else if (io_validin) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_CIsDominant <= mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant;
    end
    if (metaReset) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_CDom_CAlignDist <= 6'h0;
    end else if (io_validin) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_CDom_CAlignDist <= mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist;
    end
    if (metaReset) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_highAlignedSigC <= 55'h0;
    end else if (io_validin) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_highAlignedSigC <= mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC;
    end
    if (metaReset) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_bit0AlignedSigC <= 1'h0;
    end else if (io_validin) begin
      mulAddRecFNToRaw_postMul_io_fromPreMul_b_bit0AlignedSigC <= mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC;
    end
    if (metaReset) begin
      mulAddRecFNToRaw_postMul_io_mulAddResult_b <= 107'h0;
    end else if (io_validin) begin
      mulAddRecFNToRaw_postMul_io_mulAddResult_b <= mulAddResult;
    end
    if (metaReset) begin
      mulAddRecFNToRaw_postMul_io_roundingMode_b <= 3'h0;
    end else if (io_validin) begin
      mulAddRecFNToRaw_postMul_io_roundingMode_b <= io_roundingMode;
    end
    if (metaReset) begin
      roundingMode_stage0_b <= 3'h0;
    end else if (io_validin) begin
      roundingMode_stage0_b <= io_roundingMode;
    end
    if (metaReset) begin
      detectTininess_stage0_b <= 1'h0;
    end else begin
      detectTininess_stage0_b <= io_validin | detectTininess_stage0_b;
    end
    if (metaReset) begin
      valid_stage0_v <= 1'h0;
    end else if (reset) begin
      valid_stage0_v <= 1'h0;
    end else begin
      valid_stage0_v <= io_validin;
    end
    if (metaReset) begin
      roundRawFNToRecFN_io_invalidExc_b <= 1'h0;
    end else if (valid_stage0_v) begin
      roundRawFNToRecFN_io_invalidExc_b <= mulAddRecFNToRaw_postMul_io_invalidExc;
    end
    if (metaReset) begin
      roundRawFNToRecFN_io_in_b_isNaN <= 1'h0;
    end else if (valid_stage0_v) begin
      roundRawFNToRecFN_io_in_b_isNaN <= mulAddRecFNToRaw_postMul_io_rawOut_isNaN;
    end
    if (metaReset) begin
      roundRawFNToRecFN_io_in_b_isInf <= 1'h0;
    end else if (valid_stage0_v) begin
      roundRawFNToRecFN_io_in_b_isInf <= mulAddRecFNToRaw_postMul_io_rawOut_isInf;
    end
    if (metaReset) begin
      roundRawFNToRecFN_io_in_b_isZero <= 1'h0;
    end else if (valid_stage0_v) begin
      roundRawFNToRecFN_io_in_b_isZero <= mulAddRecFNToRaw_postMul_io_rawOut_isZero;
    end
    if (metaReset) begin
      roundRawFNToRecFN_io_in_b_sign <= 1'h0;
    end else if (valid_stage0_v) begin
      roundRawFNToRecFN_io_in_b_sign <= mulAddRecFNToRaw_postMul_io_rawOut_sign;
    end
    if (metaReset) begin
      roundRawFNToRecFN_io_in_b_sExp <= 13'h0;
    end else if (valid_stage0_v) begin
      roundRawFNToRecFN_io_in_b_sExp <= mulAddRecFNToRaw_postMul_io_rawOut_sExp;
    end
    if (metaReset) begin
      roundRawFNToRecFN_io_in_b_sig <= 56'h0;
    end else if (valid_stage0_v) begin
      roundRawFNToRecFN_io_in_b_sig <= mulAddRecFNToRaw_postMul_io_rawOut_sig;
    end
    if (metaReset) begin
      roundRawFNToRecFN_io_roundingMode_b <= 3'h0;
    end else if (valid_stage0_v) begin
      roundRawFNToRecFN_io_roundingMode_b <= roundingMode_stage0_b;
    end
    if (metaReset) begin
      roundRawFNToRecFN_io_detectTininess_b <= 1'h0;
    end else if (valid_stage0_v) begin
      roundRawFNToRecFN_io_detectTininess_b <= detectTininess_stage0_b;
    end
    if (metaReset) begin
      io_validout_v <= 1'h0;
    end else if (reset) begin
      io_validout_v <= 1'h0;
    end else begin
      io_validout_v <= valid_stage0_v;
    end
    MulAddRecFNPipe_1_state <= valid_stage0_v_pad;
    if (!(MulAddRecFNPipe_1_cov_read_data)) begin
      MulAddRecFNPipe_1_covSum <= MulAddRecFNPipe_1_covSum + 1'h1;
    end
    if (metaReset) begin
      MulAddRecFNPipe_1_metaAssert <= 1'h0;
    end else begin
      MulAddRecFNPipe_1_metaAssert <= MulAddRecFNPipe_1_metaAssert | MulAddRecFNPipe_1_or0;
    end
  end
  always @(posedge clock) begin
    if(MulAddRecFNPipe_1_cov_write_en & MulAddRecFNPipe_1_cov_write_mask) begin
      MulAddRecFNPipe_1_cov[MulAddRecFNPipe_1_cov_write_addr] <= MulAddRecFNPipe_1_cov_write_data; // @[Coverage map for MulAddRecFNPipe_1]
    end
  end
endmodule
module DivSqrtRecFNToRaw_small(
  input         clock,
  input         reset,
  output        io_inReady,
  input         io_inValid,
  input         io_sqrtOp,
  input  [32:0] io_a,
  input  [32:0] io_b,
  input  [2:0]  io_roundingMode,
  output        io_rawOutValid_div,
  output        io_rawOutValid_sqrt,
  output [2:0]  io_roundingModeOut,
  output        io_invalidExc,
  output        io_infiniteExc,
  output        io_rawOut_isNaN,
  output        io_rawOut_isInf,
  output        io_rawOut_isZero,
  output        io_rawOut_sign,
  output [9:0]  io_rawOut_sExp,
  output [26:0] io_rawOut_sig,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset,
  input         divSqrtRawFN__halt
);
  wire  divSqrtRawFN__clock; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN__reset; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN__io_inReady; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN__io_inValid; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN__io_sqrtOp; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN__io_a_isNaN; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN__io_a_isInf; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN__io_a_isZero; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN__io_a_sign; // @[DivSqrtRecFN_small.scala 416:15]
  wire [9:0] divSqrtRawFN__io_a_sExp; // @[DivSqrtRecFN_small.scala 416:15]
  wire [24:0] divSqrtRawFN__io_a_sig; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN__io_b_isNaN; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN__io_b_isInf; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN__io_b_isZero; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN__io_b_sign; // @[DivSqrtRecFN_small.scala 416:15]
  wire [9:0] divSqrtRawFN__io_b_sExp; // @[DivSqrtRecFN_small.scala 416:15]
  wire [24:0] divSqrtRawFN__io_b_sig; // @[DivSqrtRecFN_small.scala 416:15]
  wire [2:0] divSqrtRawFN__io_roundingMode; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN__io_rawOutValid_div; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN__io_rawOutValid_sqrt; // @[DivSqrtRecFN_small.scala 416:15]
  wire [2:0] divSqrtRawFN__io_roundingModeOut; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN__io_invalidExc; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN__io_infiniteExc; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN__io_rawOut_isNaN; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN__io_rawOut_isInf; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN__io_rawOut_isZero; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN__io_rawOut_sign; // @[DivSqrtRecFN_small.scala 416:15]
  wire [9:0] divSqrtRawFN__io_rawOut_sExp; // @[DivSqrtRecFN_small.scala 416:15]
  wire [26:0] divSqrtRawFN__io_rawOut_sig; // @[DivSqrtRecFN_small.scala 416:15]
  wire [29:0] divSqrtRawFN__io_covSum; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN__metaAssert; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN__metaReset; // @[DivSqrtRecFN_small.scala 416:15]
  wire [8:0] divSqrtRawFN_io_a_exp; // @[rawFloatFromRecFN.scala 50:21]
  wire  divSqrtRawFN_io_a_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  divSqrtRawFN_io_a_isSpecial; // @[rawFloatFromRecFN.scala 52:54]
  wire  divSqrtRawFN_io_a_out_sig_hi_lo; // @[rawFloatFromRecFN.scala 60:39]
  wire [22:0] divSqrtRawFN_io_a_out_sig_lo; // @[rawFloatFromRecFN.scala 60:51]
  wire [1:0] divSqrtRawFN_io_a_out_sig_hi; // @[Cat.scala 30:58]
  wire [8:0] divSqrtRawFN_io_b_exp; // @[rawFloatFromRecFN.scala 50:21]
  wire  divSqrtRawFN_io_b_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  divSqrtRawFN_io_b_isSpecial; // @[rawFloatFromRecFN.scala 52:54]
  wire  divSqrtRawFN_io_b_out_sig_hi_lo; // @[rawFloatFromRecFN.scala 60:39]
  wire [22:0] divSqrtRawFN_io_b_out_sig_lo; // @[rawFloatFromRecFN.scala 60:51]
  wire [1:0] divSqrtRawFN_io_b_out_sig_hi; // @[Cat.scala 30:58]
  wire [29:0] DivSqrtRecFNToRaw_small_covSum;
  wire [29:0] divSqrtRawFN__sum;
  wire  divSqrtRawFN__metaAssert_wire;
  reg  DivSqrtRecFNToRaw_small_metaAssert;
  reg [31:0] _RAND_0;
  DivSqrtRawFN_small divSqrtRawFN_ ( // @[DivSqrtRecFN_small.scala 416:15]
    .clock(divSqrtRawFN__clock),
    .reset(divSqrtRawFN__reset),
    .io_inReady(divSqrtRawFN__io_inReady),
    .io_inValid(divSqrtRawFN__io_inValid),
    .io_sqrtOp(divSqrtRawFN__io_sqrtOp),
    .io_a_isNaN(divSqrtRawFN__io_a_isNaN),
    .io_a_isInf(divSqrtRawFN__io_a_isInf),
    .io_a_isZero(divSqrtRawFN__io_a_isZero),
    .io_a_sign(divSqrtRawFN__io_a_sign),
    .io_a_sExp(divSqrtRawFN__io_a_sExp),
    .io_a_sig(divSqrtRawFN__io_a_sig),
    .io_b_isNaN(divSqrtRawFN__io_b_isNaN),
    .io_b_isInf(divSqrtRawFN__io_b_isInf),
    .io_b_isZero(divSqrtRawFN__io_b_isZero),
    .io_b_sign(divSqrtRawFN__io_b_sign),
    .io_b_sExp(divSqrtRawFN__io_b_sExp),
    .io_b_sig(divSqrtRawFN__io_b_sig),
    .io_roundingMode(divSqrtRawFN__io_roundingMode),
    .io_rawOutValid_div(divSqrtRawFN__io_rawOutValid_div),
    .io_rawOutValid_sqrt(divSqrtRawFN__io_rawOutValid_sqrt),
    .io_roundingModeOut(divSqrtRawFN__io_roundingModeOut),
    .io_invalidExc(divSqrtRawFN__io_invalidExc),
    .io_infiniteExc(divSqrtRawFN__io_infiniteExc),
    .io_rawOut_isNaN(divSqrtRawFN__io_rawOut_isNaN),
    .io_rawOut_isInf(divSqrtRawFN__io_rawOut_isInf),
    .io_rawOut_isZero(divSqrtRawFN__io_rawOut_isZero),
    .io_rawOut_sign(divSqrtRawFN__io_rawOut_sign),
    .io_rawOut_sExp(divSqrtRawFN__io_rawOut_sExp),
    .io_rawOut_sig(divSqrtRawFN__io_rawOut_sig),
    .io_covSum(divSqrtRawFN__io_covSum),
    .metaAssert(divSqrtRawFN__metaAssert),
    .metaReset(divSqrtRawFN__metaReset)
  );
  assign divSqrtRawFN_io_a_exp = io_a[31:23]; // @[rawFloatFromRecFN.scala 50:21]
  assign divSqrtRawFN_io_a_isZero = divSqrtRawFN_io_a_exp[8:6] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign divSqrtRawFN_io_a_isSpecial = divSqrtRawFN_io_a_exp[8:7] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign divSqrtRawFN_io_a_out_sig_hi_lo = ~divSqrtRawFN_io_a_isZero; // @[rawFloatFromRecFN.scala 60:39]
  assign divSqrtRawFN_io_a_out_sig_lo = io_a[22:0]; // @[rawFloatFromRecFN.scala 60:51]
  assign divSqrtRawFN_io_a_out_sig_hi = {1'h0,divSqrtRawFN_io_a_out_sig_hi_lo}; // @[Cat.scala 30:58]
  assign divSqrtRawFN_io_b_exp = io_b[31:23]; // @[rawFloatFromRecFN.scala 50:21]
  assign divSqrtRawFN_io_b_isZero = divSqrtRawFN_io_b_exp[8:6] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign divSqrtRawFN_io_b_isSpecial = divSqrtRawFN_io_b_exp[8:7] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign divSqrtRawFN_io_b_out_sig_hi_lo = ~divSqrtRawFN_io_b_isZero; // @[rawFloatFromRecFN.scala 60:39]
  assign divSqrtRawFN_io_b_out_sig_lo = io_b[22:0]; // @[rawFloatFromRecFN.scala 60:51]
  assign divSqrtRawFN_io_b_out_sig_hi = {1'h0,divSqrtRawFN_io_b_out_sig_hi_lo}; // @[Cat.scala 30:58]
  assign io_inReady = divSqrtRawFN__io_inReady; // @[DivSqrtRecFN_small.scala 418:16]
  assign io_rawOutValid_div = divSqrtRawFN__io_rawOutValid_div; // @[DivSqrtRecFN_small.scala 425:25]
  assign io_rawOutValid_sqrt = divSqrtRawFN__io_rawOutValid_sqrt; // @[DivSqrtRecFN_small.scala 426:25]
  assign io_roundingModeOut = divSqrtRawFN__io_roundingModeOut; // @[DivSqrtRecFN_small.scala 427:25]
  assign io_invalidExc = divSqrtRawFN__io_invalidExc; // @[DivSqrtRecFN_small.scala 428:25]
  assign io_infiniteExc = divSqrtRawFN__io_infiniteExc; // @[DivSqrtRecFN_small.scala 429:25]
  assign io_rawOut_isNaN = divSqrtRawFN__io_rawOut_isNaN; // @[DivSqrtRecFN_small.scala 430:25]
  assign io_rawOut_isInf = divSqrtRawFN__io_rawOut_isInf; // @[DivSqrtRecFN_small.scala 430:25]
  assign io_rawOut_isZero = divSqrtRawFN__io_rawOut_isZero; // @[DivSqrtRecFN_small.scala 430:25]
  assign io_rawOut_sign = divSqrtRawFN__io_rawOut_sign; // @[DivSqrtRecFN_small.scala 430:25]
  assign io_rawOut_sExp = divSqrtRawFN__io_rawOut_sExp; // @[DivSqrtRecFN_small.scala 430:25]
  assign io_rawOut_sig = divSqrtRawFN__io_rawOut_sig; // @[DivSqrtRecFN_small.scala 430:25]
  assign divSqrtRawFN__clock = clock;
  assign divSqrtRawFN__reset = reset;
  assign divSqrtRawFN__io_inValid = io_inValid; // @[DivSqrtRecFN_small.scala 419:34]
  assign divSqrtRawFN__io_sqrtOp = io_sqrtOp; // @[DivSqrtRecFN_small.scala 420:34]
  assign divSqrtRawFN__io_a_isNaN = divSqrtRawFN_io_a_isSpecial & divSqrtRawFN_io_a_exp[6]; // @[DivSqrtRecFN_small.scala 421:34]
  assign divSqrtRawFN__io_a_isInf = divSqrtRawFN_io_a_isSpecial & ~divSqrtRawFN_io_a_exp[6]; // @[DivSqrtRecFN_small.scala 421:34]
  assign divSqrtRawFN__io_a_isZero = divSqrtRawFN_io_a_exp[8:6] == 3'h0; // @[DivSqrtRecFN_small.scala 421:34]
  assign divSqrtRawFN__io_a_sign = io_a[32]; // @[DivSqrtRecFN_small.scala 421:34]
  assign divSqrtRawFN__io_a_sExp = {1'b0,$signed(divSqrtRawFN_io_a_exp)}; // @[DivSqrtRecFN_small.scala 421:34]
  assign divSqrtRawFN__io_a_sig = {divSqrtRawFN_io_a_out_sig_hi,divSqrtRawFN_io_a_out_sig_lo}; // @[DivSqrtRecFN_small.scala 421:34]
  assign divSqrtRawFN__io_b_isNaN = divSqrtRawFN_io_b_isSpecial & divSqrtRawFN_io_b_exp[6]; // @[DivSqrtRecFN_small.scala 422:34]
  assign divSqrtRawFN__io_b_isInf = divSqrtRawFN_io_b_isSpecial & ~divSqrtRawFN_io_b_exp[6]; // @[DivSqrtRecFN_small.scala 422:34]
  assign divSqrtRawFN__io_b_isZero = divSqrtRawFN_io_b_exp[8:6] == 3'h0; // @[DivSqrtRecFN_small.scala 422:34]
  assign divSqrtRawFN__io_b_sign = io_b[32]; // @[DivSqrtRecFN_small.scala 422:34]
  assign divSqrtRawFN__io_b_sExp = {1'b0,$signed(divSqrtRawFN_io_b_exp)}; // @[DivSqrtRecFN_small.scala 422:34]
  assign divSqrtRawFN__io_b_sig = {divSqrtRawFN_io_b_out_sig_hi,divSqrtRawFN_io_b_out_sig_lo}; // @[DivSqrtRecFN_small.scala 422:34]
  assign divSqrtRawFN__io_roundingMode = io_roundingMode; // @[DivSqrtRecFN_small.scala 423:34]
  assign DivSqrtRecFNToRaw_small_covSum = 30'h0;
  assign divSqrtRawFN__sum = DivSqrtRecFNToRaw_small_covSum + divSqrtRawFN__io_covSum;
  assign io_covSum = divSqrtRawFN__sum;
  assign divSqrtRawFN__metaAssert_wire = divSqrtRawFN__metaAssert;
  assign metaAssert = DivSqrtRecFNToRaw_small_metaAssert;
  assign divSqrtRawFN__metaReset = metaReset | divSqrtRawFN__halt;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  DivSqrtRecFNToRaw_small_metaAssert = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      DivSqrtRecFNToRaw_small_metaAssert <= 1'h0;
    end else begin
      DivSqrtRecFNToRaw_small_metaAssert <= DivSqrtRecFNToRaw_small_metaAssert | divSqrtRawFN__metaAssert_wire;
    end
  end
endmodule
module RoundRawFNToRecFN_2(
  input         io_invalidExc,
  input         io_infiniteExc,
  input         io_in_isNaN,
  input         io_in_isInf,
  input         io_in_isZero,
  input         io_in_sign,
  input  [9:0]  io_in_sExp,
  input  [26:0] io_in_sig,
  input  [2:0]  io_roundingMode,
  input         io_detectTininess,
  output [32:0] io_out,
  output [4:0]  io_exceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  roundAnyRawFNToRecFN_io_invalidExc; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_infiniteExc; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_sign; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [9:0] roundAnyRawFNToRecFN_io_in_sExp; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [26:0] roundAnyRawFNToRecFN_io_in_sig; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [2:0] roundAnyRawFNToRecFN_io_roundingMode; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_detectTininess; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [32:0] roundAnyRawFNToRecFN_io_out; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [4:0] roundAnyRawFNToRecFN_io_exceptionFlags; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [29:0] roundAnyRawFNToRecFN_io_covSum; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_metaAssert; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [29:0] RoundRawFNToRecFN_2_covSum;
  wire [29:0] roundAnyRawFNToRecFN_sum;
  wire  roundAnyRawFNToRecFN_metaAssert_wire;
  RoundAnyRawFNToRecFN_5 roundAnyRawFNToRecFN ( // @[RoundAnyRawFNToRecFN.scala 307:15]
    .io_invalidExc(roundAnyRawFNToRecFN_io_invalidExc),
    .io_infiniteExc(roundAnyRawFNToRecFN_io_infiniteExc),
    .io_in_isNaN(roundAnyRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundAnyRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundAnyRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundAnyRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundAnyRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundAnyRawFNToRecFN_io_in_sig),
    .io_roundingMode(roundAnyRawFNToRecFN_io_roundingMode),
    .io_detectTininess(roundAnyRawFNToRecFN_io_detectTininess),
    .io_out(roundAnyRawFNToRecFN_io_out),
    .io_exceptionFlags(roundAnyRawFNToRecFN_io_exceptionFlags),
    .io_covSum(roundAnyRawFNToRecFN_io_covSum),
    .metaAssert(roundAnyRawFNToRecFN_metaAssert)
  );
  assign io_out = roundAnyRawFNToRecFN_io_out; // @[RoundAnyRawFNToRecFN.scala 315:23]
  assign io_exceptionFlags = roundAnyRawFNToRecFN_io_exceptionFlags; // @[RoundAnyRawFNToRecFN.scala 316:23]
  assign roundAnyRawFNToRecFN_io_invalidExc = io_invalidExc; // @[RoundAnyRawFNToRecFN.scala 310:44]
  assign roundAnyRawFNToRecFN_io_infiniteExc = io_infiniteExc; // @[RoundAnyRawFNToRecFN.scala 311:44]
  assign roundAnyRawFNToRecFN_io_in_isNaN = io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_isInf = io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_isZero = io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_sign = io_in_sign; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_sExp = io_in_sExp; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_sig = io_in_sig; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_roundingMode = io_roundingMode; // @[RoundAnyRawFNToRecFN.scala 313:44]
  assign roundAnyRawFNToRecFN_io_detectTininess = io_detectTininess; // @[RoundAnyRawFNToRecFN.scala 314:44]
  assign RoundRawFNToRecFN_2_covSum = 30'h0;
  assign roundAnyRawFNToRecFN_sum = RoundRawFNToRecFN_2_covSum + roundAnyRawFNToRecFN_io_covSum;
  assign io_covSum = roundAnyRawFNToRecFN_sum;
  assign roundAnyRawFNToRecFN_metaAssert_wire = roundAnyRawFNToRecFN_metaAssert;
  assign metaAssert = roundAnyRawFNToRecFN_metaAssert_wire;
endmodule
module DivSqrtRecFNToRaw_small_1(
  input         clock,
  input         reset,
  output        io_inReady,
  input         io_inValid,
  input         io_sqrtOp,
  input  [64:0] io_a,
  input  [64:0] io_b,
  input  [2:0]  io_roundingMode,
  output        io_rawOutValid_div,
  output        io_rawOutValid_sqrt,
  output [2:0]  io_roundingModeOut,
  output        io_invalidExc,
  output        io_infiniteExc,
  output        io_rawOut_isNaN,
  output        io_rawOut_isInf,
  output        io_rawOut_isZero,
  output        io_rawOut_sign,
  output [12:0] io_rawOut_sExp,
  output [55:0] io_rawOut_sig,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset,
  input         divSqrtRawFN__halt
);
  wire  divSqrtRawFN__clock; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN__reset; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN__io_inReady; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN__io_inValid; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN__io_sqrtOp; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN__io_a_isNaN; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN__io_a_isInf; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN__io_a_isZero; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN__io_a_sign; // @[DivSqrtRecFN_small.scala 416:15]
  wire [12:0] divSqrtRawFN__io_a_sExp; // @[DivSqrtRecFN_small.scala 416:15]
  wire [53:0] divSqrtRawFN__io_a_sig; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN__io_b_isNaN; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN__io_b_isInf; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN__io_b_isZero; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN__io_b_sign; // @[DivSqrtRecFN_small.scala 416:15]
  wire [12:0] divSqrtRawFN__io_b_sExp; // @[DivSqrtRecFN_small.scala 416:15]
  wire [53:0] divSqrtRawFN__io_b_sig; // @[DivSqrtRecFN_small.scala 416:15]
  wire [2:0] divSqrtRawFN__io_roundingMode; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN__io_rawOutValid_div; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN__io_rawOutValid_sqrt; // @[DivSqrtRecFN_small.scala 416:15]
  wire [2:0] divSqrtRawFN__io_roundingModeOut; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN__io_invalidExc; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN__io_infiniteExc; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN__io_rawOut_isNaN; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN__io_rawOut_isInf; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN__io_rawOut_isZero; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN__io_rawOut_sign; // @[DivSqrtRecFN_small.scala 416:15]
  wire [12:0] divSqrtRawFN__io_rawOut_sExp; // @[DivSqrtRecFN_small.scala 416:15]
  wire [55:0] divSqrtRawFN__io_rawOut_sig; // @[DivSqrtRecFN_small.scala 416:15]
  wire [29:0] divSqrtRawFN__io_covSum; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN__metaAssert; // @[DivSqrtRecFN_small.scala 416:15]
  wire  divSqrtRawFN__metaReset; // @[DivSqrtRecFN_small.scala 416:15]
  wire [11:0] divSqrtRawFN_io_a_exp; // @[rawFloatFromRecFN.scala 50:21]
  wire  divSqrtRawFN_io_a_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  divSqrtRawFN_io_a_isSpecial; // @[rawFloatFromRecFN.scala 52:54]
  wire  divSqrtRawFN_io_a_out_sig_hi_lo; // @[rawFloatFromRecFN.scala 60:39]
  wire [51:0] divSqrtRawFN_io_a_out_sig_lo; // @[rawFloatFromRecFN.scala 60:51]
  wire [1:0] divSqrtRawFN_io_a_out_sig_hi; // @[Cat.scala 30:58]
  wire [11:0] divSqrtRawFN_io_b_exp; // @[rawFloatFromRecFN.scala 50:21]
  wire  divSqrtRawFN_io_b_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  divSqrtRawFN_io_b_isSpecial; // @[rawFloatFromRecFN.scala 52:54]
  wire  divSqrtRawFN_io_b_out_sig_hi_lo; // @[rawFloatFromRecFN.scala 60:39]
  wire [51:0] divSqrtRawFN_io_b_out_sig_lo; // @[rawFloatFromRecFN.scala 60:51]
  wire [1:0] divSqrtRawFN_io_b_out_sig_hi; // @[Cat.scala 30:58]
  wire [29:0] DivSqrtRecFNToRaw_small_1_covSum;
  wire [29:0] divSqrtRawFN__sum;
  wire  divSqrtRawFN__metaAssert_wire;
  reg  DivSqrtRecFNToRaw_small_1_metaAssert;
  reg [31:0] _RAND_0;
  DivSqrtRawFN_small_1 divSqrtRawFN_ ( // @[DivSqrtRecFN_small.scala 416:15]
    .clock(divSqrtRawFN__clock),
    .reset(divSqrtRawFN__reset),
    .io_inReady(divSqrtRawFN__io_inReady),
    .io_inValid(divSqrtRawFN__io_inValid),
    .io_sqrtOp(divSqrtRawFN__io_sqrtOp),
    .io_a_isNaN(divSqrtRawFN__io_a_isNaN),
    .io_a_isInf(divSqrtRawFN__io_a_isInf),
    .io_a_isZero(divSqrtRawFN__io_a_isZero),
    .io_a_sign(divSqrtRawFN__io_a_sign),
    .io_a_sExp(divSqrtRawFN__io_a_sExp),
    .io_a_sig(divSqrtRawFN__io_a_sig),
    .io_b_isNaN(divSqrtRawFN__io_b_isNaN),
    .io_b_isInf(divSqrtRawFN__io_b_isInf),
    .io_b_isZero(divSqrtRawFN__io_b_isZero),
    .io_b_sign(divSqrtRawFN__io_b_sign),
    .io_b_sExp(divSqrtRawFN__io_b_sExp),
    .io_b_sig(divSqrtRawFN__io_b_sig),
    .io_roundingMode(divSqrtRawFN__io_roundingMode),
    .io_rawOutValid_div(divSqrtRawFN__io_rawOutValid_div),
    .io_rawOutValid_sqrt(divSqrtRawFN__io_rawOutValid_sqrt),
    .io_roundingModeOut(divSqrtRawFN__io_roundingModeOut),
    .io_invalidExc(divSqrtRawFN__io_invalidExc),
    .io_infiniteExc(divSqrtRawFN__io_infiniteExc),
    .io_rawOut_isNaN(divSqrtRawFN__io_rawOut_isNaN),
    .io_rawOut_isInf(divSqrtRawFN__io_rawOut_isInf),
    .io_rawOut_isZero(divSqrtRawFN__io_rawOut_isZero),
    .io_rawOut_sign(divSqrtRawFN__io_rawOut_sign),
    .io_rawOut_sExp(divSqrtRawFN__io_rawOut_sExp),
    .io_rawOut_sig(divSqrtRawFN__io_rawOut_sig),
    .io_covSum(divSqrtRawFN__io_covSum),
    .metaAssert(divSqrtRawFN__metaAssert),
    .metaReset(divSqrtRawFN__metaReset)
  );
  assign divSqrtRawFN_io_a_exp = io_a[63:52]; // @[rawFloatFromRecFN.scala 50:21]
  assign divSqrtRawFN_io_a_isZero = divSqrtRawFN_io_a_exp[11:9] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign divSqrtRawFN_io_a_isSpecial = divSqrtRawFN_io_a_exp[11:10] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign divSqrtRawFN_io_a_out_sig_hi_lo = ~divSqrtRawFN_io_a_isZero; // @[rawFloatFromRecFN.scala 60:39]
  assign divSqrtRawFN_io_a_out_sig_lo = io_a[51:0]; // @[rawFloatFromRecFN.scala 60:51]
  assign divSqrtRawFN_io_a_out_sig_hi = {1'h0,divSqrtRawFN_io_a_out_sig_hi_lo}; // @[Cat.scala 30:58]
  assign divSqrtRawFN_io_b_exp = io_b[63:52]; // @[rawFloatFromRecFN.scala 50:21]
  assign divSqrtRawFN_io_b_isZero = divSqrtRawFN_io_b_exp[11:9] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign divSqrtRawFN_io_b_isSpecial = divSqrtRawFN_io_b_exp[11:10] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign divSqrtRawFN_io_b_out_sig_hi_lo = ~divSqrtRawFN_io_b_isZero; // @[rawFloatFromRecFN.scala 60:39]
  assign divSqrtRawFN_io_b_out_sig_lo = io_b[51:0]; // @[rawFloatFromRecFN.scala 60:51]
  assign divSqrtRawFN_io_b_out_sig_hi = {1'h0,divSqrtRawFN_io_b_out_sig_hi_lo}; // @[Cat.scala 30:58]
  assign io_inReady = divSqrtRawFN__io_inReady; // @[DivSqrtRecFN_small.scala 418:16]
  assign io_rawOutValid_div = divSqrtRawFN__io_rawOutValid_div; // @[DivSqrtRecFN_small.scala 425:25]
  assign io_rawOutValid_sqrt = divSqrtRawFN__io_rawOutValid_sqrt; // @[DivSqrtRecFN_small.scala 426:25]
  assign io_roundingModeOut = divSqrtRawFN__io_roundingModeOut; // @[DivSqrtRecFN_small.scala 427:25]
  assign io_invalidExc = divSqrtRawFN__io_invalidExc; // @[DivSqrtRecFN_small.scala 428:25]
  assign io_infiniteExc = divSqrtRawFN__io_infiniteExc; // @[DivSqrtRecFN_small.scala 429:25]
  assign io_rawOut_isNaN = divSqrtRawFN__io_rawOut_isNaN; // @[DivSqrtRecFN_small.scala 430:25]
  assign io_rawOut_isInf = divSqrtRawFN__io_rawOut_isInf; // @[DivSqrtRecFN_small.scala 430:25]
  assign io_rawOut_isZero = divSqrtRawFN__io_rawOut_isZero; // @[DivSqrtRecFN_small.scala 430:25]
  assign io_rawOut_sign = divSqrtRawFN__io_rawOut_sign; // @[DivSqrtRecFN_small.scala 430:25]
  assign io_rawOut_sExp = divSqrtRawFN__io_rawOut_sExp; // @[DivSqrtRecFN_small.scala 430:25]
  assign io_rawOut_sig = divSqrtRawFN__io_rawOut_sig; // @[DivSqrtRecFN_small.scala 430:25]
  assign divSqrtRawFN__clock = clock;
  assign divSqrtRawFN__reset = reset;
  assign divSqrtRawFN__io_inValid = io_inValid; // @[DivSqrtRecFN_small.scala 419:34]
  assign divSqrtRawFN__io_sqrtOp = io_sqrtOp; // @[DivSqrtRecFN_small.scala 420:34]
  assign divSqrtRawFN__io_a_isNaN = divSqrtRawFN_io_a_isSpecial & divSqrtRawFN_io_a_exp[9]; // @[DivSqrtRecFN_small.scala 421:34]
  assign divSqrtRawFN__io_a_isInf = divSqrtRawFN_io_a_isSpecial & ~divSqrtRawFN_io_a_exp[9]; // @[DivSqrtRecFN_small.scala 421:34]
  assign divSqrtRawFN__io_a_isZero = divSqrtRawFN_io_a_exp[11:9] == 3'h0; // @[DivSqrtRecFN_small.scala 421:34]
  assign divSqrtRawFN__io_a_sign = io_a[64]; // @[DivSqrtRecFN_small.scala 421:34]
  assign divSqrtRawFN__io_a_sExp = {1'b0,$signed(divSqrtRawFN_io_a_exp)}; // @[DivSqrtRecFN_small.scala 421:34]
  assign divSqrtRawFN__io_a_sig = {divSqrtRawFN_io_a_out_sig_hi,divSqrtRawFN_io_a_out_sig_lo}; // @[DivSqrtRecFN_small.scala 421:34]
  assign divSqrtRawFN__io_b_isNaN = divSqrtRawFN_io_b_isSpecial & divSqrtRawFN_io_b_exp[9]; // @[DivSqrtRecFN_small.scala 422:34]
  assign divSqrtRawFN__io_b_isInf = divSqrtRawFN_io_b_isSpecial & ~divSqrtRawFN_io_b_exp[9]; // @[DivSqrtRecFN_small.scala 422:34]
  assign divSqrtRawFN__io_b_isZero = divSqrtRawFN_io_b_exp[11:9] == 3'h0; // @[DivSqrtRecFN_small.scala 422:34]
  assign divSqrtRawFN__io_b_sign = io_b[64]; // @[DivSqrtRecFN_small.scala 422:34]
  assign divSqrtRawFN__io_b_sExp = {1'b0,$signed(divSqrtRawFN_io_b_exp)}; // @[DivSqrtRecFN_small.scala 422:34]
  assign divSqrtRawFN__io_b_sig = {divSqrtRawFN_io_b_out_sig_hi,divSqrtRawFN_io_b_out_sig_lo}; // @[DivSqrtRecFN_small.scala 422:34]
  assign divSqrtRawFN__io_roundingMode = io_roundingMode; // @[DivSqrtRecFN_small.scala 423:34]
  assign DivSqrtRecFNToRaw_small_1_covSum = 30'h0;
  assign divSqrtRawFN__sum = DivSqrtRecFNToRaw_small_1_covSum + divSqrtRawFN__io_covSum;
  assign io_covSum = divSqrtRawFN__sum;
  assign divSqrtRawFN__metaAssert_wire = divSqrtRawFN__metaAssert;
  assign metaAssert = DivSqrtRecFNToRaw_small_1_metaAssert;
  assign divSqrtRawFN__metaReset = metaReset | divSqrtRawFN__halt;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  DivSqrtRecFNToRaw_small_1_metaAssert = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      DivSqrtRecFNToRaw_small_1_metaAssert <= 1'h0;
    end else begin
      DivSqrtRecFNToRaw_small_1_metaAssert <= DivSqrtRecFNToRaw_small_1_metaAssert | divSqrtRawFN__metaAssert_wire;
    end
  end
endmodule
module RoundRawFNToRecFN_3(
  input         io_invalidExc,
  input         io_infiniteExc,
  input         io_in_isNaN,
  input         io_in_isInf,
  input         io_in_isZero,
  input         io_in_sign,
  input  [12:0] io_in_sExp,
  input  [55:0] io_in_sig,
  input  [2:0]  io_roundingMode,
  input         io_detectTininess,
  output [64:0] io_out,
  output [4:0]  io_exceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  roundAnyRawFNToRecFN_io_invalidExc; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_infiniteExc; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_sign; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [12:0] roundAnyRawFNToRecFN_io_in_sExp; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [55:0] roundAnyRawFNToRecFN_io_in_sig; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [2:0] roundAnyRawFNToRecFN_io_roundingMode; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_detectTininess; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [64:0] roundAnyRawFNToRecFN_io_out; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [4:0] roundAnyRawFNToRecFN_io_exceptionFlags; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [29:0] roundAnyRawFNToRecFN_io_covSum; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_metaAssert; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [29:0] RoundRawFNToRecFN_3_covSum;
  wire [29:0] roundAnyRawFNToRecFN_sum;
  wire  roundAnyRawFNToRecFN_metaAssert_wire;
  RoundAnyRawFNToRecFN_6 roundAnyRawFNToRecFN ( // @[RoundAnyRawFNToRecFN.scala 307:15]
    .io_invalidExc(roundAnyRawFNToRecFN_io_invalidExc),
    .io_infiniteExc(roundAnyRawFNToRecFN_io_infiniteExc),
    .io_in_isNaN(roundAnyRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundAnyRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundAnyRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundAnyRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundAnyRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundAnyRawFNToRecFN_io_in_sig),
    .io_roundingMode(roundAnyRawFNToRecFN_io_roundingMode),
    .io_detectTininess(roundAnyRawFNToRecFN_io_detectTininess),
    .io_out(roundAnyRawFNToRecFN_io_out),
    .io_exceptionFlags(roundAnyRawFNToRecFN_io_exceptionFlags),
    .io_covSum(roundAnyRawFNToRecFN_io_covSum),
    .metaAssert(roundAnyRawFNToRecFN_metaAssert)
  );
  assign io_out = roundAnyRawFNToRecFN_io_out; // @[RoundAnyRawFNToRecFN.scala 315:23]
  assign io_exceptionFlags = roundAnyRawFNToRecFN_io_exceptionFlags; // @[RoundAnyRawFNToRecFN.scala 316:23]
  assign roundAnyRawFNToRecFN_io_invalidExc = io_invalidExc; // @[RoundAnyRawFNToRecFN.scala 310:44]
  assign roundAnyRawFNToRecFN_io_infiniteExc = io_infiniteExc; // @[RoundAnyRawFNToRecFN.scala 311:44]
  assign roundAnyRawFNToRecFN_io_in_isNaN = io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_isInf = io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_isZero = io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_sign = io_in_sign; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_sExp = io_in_sExp; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_sig = io_in_sig; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_roundingMode = io_roundingMode; // @[RoundAnyRawFNToRecFN.scala 313:44]
  assign roundAnyRawFNToRecFN_io_detectTininess = io_detectTininess; // @[RoundAnyRawFNToRecFN.scala 314:44]
  assign RoundRawFNToRecFN_3_covSum = 30'h0;
  assign roundAnyRawFNToRecFN_sum = RoundRawFNToRecFN_3_covSum + roundAnyRawFNToRecFN_io_covSum;
  assign io_covSum = roundAnyRawFNToRecFN_sum;
  assign roundAnyRawFNToRecFN_metaAssert_wire = roundAnyRawFNToRecFN_metaAssert;
  assign metaAssert = roundAnyRawFNToRecFN_metaAssert_wire;
endmodule
module RVCExpander(
  input  [31:0] io_in,
  output [31:0] io_out_bits,
  output [4:0]  io_out_rd,
  output [4:0]  io_out_rs1,
  output [4:0]  io_out_rs2,
  output [4:0]  io_out_rs3,
  output        io_rvc,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  _io_out_s_opc_T_1; // @[RVC.scala 53:29]
  wire [6:0] io_out_s_lo_lo; // @[RVC.scala 53:20]
  wire [3:0] io_out_s_hi_hi_hi; // @[RVC.scala 34:26]
  wire [1:0] io_out_s_hi_hi_lo; // @[RVC.scala 34:35]
  wire  io_out_s_hi_lo; // @[RVC.scala 34:45]
  wire  io_out_s_lo_hi; // @[RVC.scala 34:51]
  wire [2:0] io_out_s_lo_1; // @[RVC.scala 31:29]
  wire [4:0] io_out_s_lo_hi_1; // @[Cat.scala 30:58]
  wire [29:0] _io_out_s_T; // @[Cat.scala 30:58]
  wire [4:0] io_out_s_0_rs3; // @[RVC.scala 20:101]
  wire [1:0] io_out_s_hi_hi_2; // @[RVC.scala 36:20]
  wire [2:0] io_out_s_hi_lo_1; // @[RVC.scala 36:28]
  wire [7:0] io_out_s_hi_hi_hi_2; // @[Cat.scala 30:58]
  wire [2:0] io_out_s_lo_5; // @[RVC.scala 30:29]
  wire [4:0] io_out_s_hi_hi_lo_1; // @[Cat.scala 30:58]
  wire [27:0] _io_out_s_T_4; // @[Cat.scala 30:58]
  wire [6:0] io_out_s_hi_hi_hi_3; // @[Cat.scala 30:58]
  wire [26:0] _io_out_s_T_9; // @[Cat.scala 30:58]
  wire [27:0] _io_out_s_T_14; // @[Cat.scala 30:58]
  wire [1:0] io_out_s_hi_hi_hi_5; // @[RVC.scala 63:32]
  wire [4:0] io_out_s_lo_hi_lo; // @[RVC.scala 63:65]
  wire [26:0] _io_out_s_T_21; // @[Cat.scala 30:58]
  wire [2:0] io_out_s_hi_hi_hi_6; // @[RVC.scala 66:30]
  wire [4:0] io_out_s_lo_hi_lo_1; // @[RVC.scala 66:63]
  wire [27:0] _io_out_s_T_28; // @[Cat.scala 30:58]
  wire [26:0] _io_out_s_T_35; // @[Cat.scala 30:58]
  wire [27:0] _io_out_s_T_42; // @[Cat.scala 30:58]
  wire [6:0] io_out_s_hi_20; // @[Bitwise.scala 72:12]
  wire [4:0] io_out_s_lo_52; // @[RVC.scala 43:38]
  wire [11:0] io_out_s_hi_hi_hi_9; // @[Cat.scala 30:58]
  wire [4:0] io_out_s_hi_hi_lo_8; // @[RVC.scala 33:13]
  wire [31:0] io_out_s_8_bits; // @[Cat.scala 30:58]
  wire  _io_out_s_opc_T_3; // @[RVC.scala 77:24]
  wire [6:0] io_out_s_lo_lo_1; // @[RVC.scala 77:20]
  wire [31:0] io_out_s_9_bits; // @[Cat.scala 30:58]
  wire [31:0] io_out_s_10_bits; // @[Cat.scala 30:58]
  wire  _io_out_s_opc_T_7; // @[RVC.scala 90:29]
  wire [6:0] io_out_s_me_lo; // @[RVC.scala 90:20]
  wire [14:0] io_out_s_me_hi_hi; // @[Bitwise.scala 72:12]
  wire [31:0] _io_out_s_me_T_2; // @[Cat.scala 30:58]
  wire [19:0] io_out_s_me_hi_hi_1; // @[RVC.scala 91:31]
  wire [31:0] io_out_s_me_bits; // @[Cat.scala 30:58]
  wire  _io_out_s_T_68; // @[RVC.scala 92:14]
  wire  _io_out_s_T_70; // @[RVC.scala 92:27]
  wire  _io_out_s_T_71; // @[RVC.scala 92:21]
  wire [6:0] io_out_s_lo_lo_2; // @[RVC.scala 86:20]
  wire [2:0] io_out_s_hi_hi_hi_12; // @[Bitwise.scala 72:12]
  wire [1:0] io_out_s_hi_hi_lo_10; // @[RVC.scala 42:42]
  wire  io_out_s_lo_hi_hi; // @[RVC.scala 42:56]
  wire [31:0] io_out_s_res_bits; // @[Cat.scala 30:58]
  wire [31:0] io_out_s_11_bits; // @[RVC.scala 92:10]
  wire [4:0] io_out_s_11_rd; // @[RVC.scala 92:10]
  wire [4:0] io_out_s_11_rs2; // @[RVC.scala 92:10]
  wire [4:0] io_out_s_11_rs3; // @[RVC.scala 92:10]
  wire [25:0] _io_out_s_T_79; // @[Cat.scala 30:58]
  wire [30:0] _GEN_0; // @[RVC.scala 99:23]
  wire [30:0] _io_out_s_T_81; // @[RVC.scala 99:23]
  wire [31:0] _io_out_s_T_84; // @[Cat.scala 30:58]
  wire [2:0] _io_out_s_funct_T; // @[Cat.scala 30:58]
  wire  _io_out_s_funct_T_1; // @[package.scala 32:86]
  wire [2:0] _io_out_s_funct_T_2; // @[package.scala 32:76]
  wire  _io_out_s_funct_T_3; // @[package.scala 32:86]
  wire [2:0] _io_out_s_funct_T_4; // @[package.scala 32:76]
  wire  _io_out_s_funct_T_5; // @[package.scala 32:86]
  wire [2:0] _io_out_s_funct_T_6; // @[package.scala 32:76]
  wire  _io_out_s_funct_T_7; // @[package.scala 32:86]
  wire [2:0] _io_out_s_funct_T_8; // @[package.scala 32:76]
  wire  _io_out_s_funct_T_9; // @[package.scala 32:86]
  wire [2:0] _io_out_s_funct_T_10; // @[package.scala 32:76]
  wire  _io_out_s_funct_T_11; // @[package.scala 32:86]
  wire [2:0] _io_out_s_funct_T_12; // @[package.scala 32:76]
  wire  _io_out_s_funct_T_13; // @[package.scala 32:86]
  wire [2:0] io_out_s_hi_lo_17; // @[package.scala 32:76]
  wire  _io_out_s_sub_T_1; // @[RVC.scala 103:30]
  wire [30:0] io_out_s_sub; // @[RVC.scala 103:22]
  wire [6:0] io_out_s_lo_lo_3; // @[RVC.scala 104:22]
  wire [24:0] _io_out_s_T_85; // @[Cat.scala 30:58]
  wire [30:0] _GEN_1; // @[RVC.scala 105:43]
  wire [30:0] _io_out_s_T_86; // @[RVC.scala 105:43]
  wire  _io_out_s_T_88; // @[package.scala 32:86]
  wire [30:0] _io_out_s_T_89; // @[package.scala 32:76]
  wire  _io_out_s_T_90; // @[package.scala 32:86]
  wire [31:0] _io_out_s_T_91; // @[package.scala 32:76]
  wire  _io_out_s_T_92; // @[package.scala 32:86]
  wire [31:0] io_out_s_12_bits; // @[package.scala 32:76]
  wire [9:0] io_out_s_hi_hi_hi_hi; // @[Bitwise.scala 72:12]
  wire  io_out_s_hi_hi_hi_lo; // @[RVC.scala 44:36]
  wire [1:0] io_out_s_hi_hi_lo_16; // @[RVC.scala 44:42]
  wire  io_out_s_hi_lo_lo; // @[RVC.scala 44:57]
  wire  io_out_s_lo_hi_lo_5; // @[RVC.scala 44:69]
  wire [2:0] io_out_s_lo_lo_hi; // @[RVC.scala 44:76]
  wire [20:0] _io_out_s_T_100; // @[Cat.scala 30:58]
  wire  io_out_s_hi_hi_hi_19; // @[RVC.scala 94:26]
  wire [9:0] io_out_s_hi_hi_lo_18; // @[RVC.scala 94:36]
  wire  io_out_s_hi_lo_21; // @[RVC.scala 94:48]
  wire [7:0] io_out_s_lo_hi_hi_5; // @[RVC.scala 94:58]
  wire [31:0] io_out_s_13_bits; // @[Cat.scala 30:58]
  wire [4:0] io_out_s_hi_hi_hi_23; // @[Bitwise.scala 72:12]
  wire [12:0] _io_out_s_T_116; // @[Cat.scala 30:58]
  wire  io_out_s_hi_hi_hi_24; // @[RVC.scala 95:29]
  wire [5:0] io_out_s_hi_hi_lo_23; // @[RVC.scala 95:39]
  wire [3:0] io_out_s_lo_hi_lo_12; // @[RVC.scala 95:71]
  wire  io_out_s_lo_lo_hi_4; // @[RVC.scala 95:82]
  wire [31:0] io_out_s_14_bits; // @[Cat.scala 30:58]
  wire [31:0] io_out_s_15_bits; // @[Cat.scala 30:58]
  wire [6:0] io_out_s_lo_lo_10; // @[RVC.scala 113:23]
  wire [25:0] _io_out_s_T_145; // @[Cat.scala 30:58]
  wire [28:0] _io_out_s_T_150; // @[Cat.scala 30:58]
  wire [1:0] io_out_s_hi_hi_47; // @[RVC.scala 37:22]
  wire [2:0] io_out_s_lo_hi_41; // @[RVC.scala 37:37]
  wire [27:0] _io_out_s_T_154; // @[Cat.scala 30:58]
  wire [28:0] _io_out_s_T_158; // @[Cat.scala 30:58]
  wire [24:0] _io_out_s_mv_T; // @[Cat.scala 30:58]
  wire [24:0] _io_out_s_add_T; // @[Cat.scala 30:58]
  wire [24:0] io_out_s_jr; // @[Cat.scala 30:58]
  wire [17:0] io_out_s_reserved_hi; // @[RVC.scala 133:29]
  wire [24:0] io_out_s_reserved; // @[Cat.scala 30:58]
  wire [24:0] _io_out_s_jr_reserved_T_2; // @[RVC.scala 134:33]
  wire  _io_out_s_jr_mv_T_1; // @[RVC.scala 135:27]
  wire [31:0] io_out_s_mv_bits; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] io_out_s_jr_reserved_bits; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] io_out_s_jr_mv_bits; // @[RVC.scala 135:22]
  wire [4:0] io_out_s_jr_mv_rd; // @[RVC.scala 135:22]
  wire [4:0] io_out_s_jr_mv_rs1; // @[RVC.scala 135:22]
  wire [4:0] io_out_s_jr_mv_rs2; // @[RVC.scala 135:22]
  wire [4:0] io_out_s_jr_mv_rs3; // @[RVC.scala 135:22]
  wire [24:0] io_out_s_jalr; // @[Cat.scala 30:58]
  wire [24:0] _io_out_s_ebreak_T; // @[Cat.scala 30:58]
  wire [24:0] io_out_s_ebreak; // @[RVC.scala 137:46]
  wire [24:0] _io_out_s_jalr_ebreak_T_2; // @[RVC.scala 138:33]
  wire [31:0] io_out_s_add_bits; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] io_out_s_jalr_ebreak_bits; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] io_out_s_jalr_add_bits; // @[RVC.scala 139:25]
  wire [4:0] io_out_s_jalr_add_rd; // @[RVC.scala 139:25]
  wire [4:0] io_out_s_jalr_add_rs1; // @[RVC.scala 139:25]
  wire [31:0] io_out_s_20_bits; // @[RVC.scala 140:10]
  wire [4:0] io_out_s_20_rd; // @[RVC.scala 140:10]
  wire [4:0] io_out_s_20_rs1; // @[RVC.scala 140:10]
  wire [4:0] io_out_s_20_rs2; // @[RVC.scala 140:10]
  wire [4:0] io_out_s_20_rs3; // @[RVC.scala 140:10]
  wire [8:0] _io_out_s_T_163; // @[Cat.scala 30:58]
  wire [3:0] io_out_s_hi_hi_hi_37; // @[RVC.scala 124:34]
  wire [4:0] io_out_s_lo_hi_lo_19; // @[RVC.scala 124:66]
  wire [28:0] _io_out_s_T_165; // @[Cat.scala 30:58]
  wire [1:0] io_out_s_hi_hi_54; // @[RVC.scala 39:22]
  wire [3:0] io_out_s_hi_lo_38; // @[RVC.scala 39:30]
  wire [7:0] _io_out_s_T_169; // @[Cat.scala 30:58]
  wire [2:0] io_out_s_hi_hi_hi_38; // @[RVC.scala 123:33]
  wire [4:0] io_out_s_lo_hi_lo_20; // @[RVC.scala 123:65]
  wire [27:0] _io_out_s_T_171; // @[Cat.scala 30:58]
  wire [28:0] _io_out_s_T_177; // @[Cat.scala 30:58]
  wire [4:0] io_out_s_24_rs1; // @[RVC.scala 20:57]
  wire [4:0] io_out_s_24_rs2; // @[RVC.scala 20:79]
  wire [2:0] io_out_lo; // @[RVC.scala 151:20]
  wire [4:0] _io_out_T; // @[Cat.scala 30:58]
  wire  _io_out_T_1; // @[package.scala 32:86]
  wire [31:0] io_out_s_1_bits; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] io_out_s_0_bits; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _io_out_T_2_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_2_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_2_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_2_rs3; // @[package.scala 32:76]
  wire  _io_out_T_3; // @[package.scala 32:86]
  wire [31:0] io_out_s_2_bits; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _io_out_T_4_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_4_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_4_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_4_rs3; // @[package.scala 32:76]
  wire  _io_out_T_5; // @[package.scala 32:86]
  wire [31:0] io_out_s_3_bits; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _io_out_T_6_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_6_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_6_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_6_rs3; // @[package.scala 32:76]
  wire  _io_out_T_7; // @[package.scala 32:86]
  wire [31:0] io_out_s_4_bits; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _io_out_T_8_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_8_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_8_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_8_rs3; // @[package.scala 32:76]
  wire  _io_out_T_9; // @[package.scala 32:86]
  wire [31:0] io_out_s_5_bits; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _io_out_T_10_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_10_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_10_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_10_rs3; // @[package.scala 32:76]
  wire  _io_out_T_11; // @[package.scala 32:86]
  wire [31:0] io_out_s_6_bits; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _io_out_T_12_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_12_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_12_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_12_rs3; // @[package.scala 32:76]
  wire  _io_out_T_13; // @[package.scala 32:86]
  wire [31:0] io_out_s_7_bits; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _io_out_T_14_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_14_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_14_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_14_rs3; // @[package.scala 32:76]
  wire  _io_out_T_15; // @[package.scala 32:86]
  wire [31:0] _io_out_T_16_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_16_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_16_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_16_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_16_rs3; // @[package.scala 32:76]
  wire  _io_out_T_17; // @[package.scala 32:86]
  wire [31:0] _io_out_T_18_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_18_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_18_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_18_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_18_rs3; // @[package.scala 32:76]
  wire  _io_out_T_19; // @[package.scala 32:86]
  wire [31:0] _io_out_T_20_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_20_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_20_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_20_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_20_rs3; // @[package.scala 32:76]
  wire  _io_out_T_21; // @[package.scala 32:86]
  wire [31:0] _io_out_T_22_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_22_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_22_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_22_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_22_rs3; // @[package.scala 32:76]
  wire  _io_out_T_23; // @[package.scala 32:86]
  wire [31:0] _io_out_T_24_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_24_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_24_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_24_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_24_rs3; // @[package.scala 32:76]
  wire  _io_out_T_25; // @[package.scala 32:86]
  wire [31:0] _io_out_T_26_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_26_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_26_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_26_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_26_rs3; // @[package.scala 32:76]
  wire  _io_out_T_27; // @[package.scala 32:86]
  wire [31:0] _io_out_T_28_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_28_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_28_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_28_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_28_rs3; // @[package.scala 32:76]
  wire  _io_out_T_29; // @[package.scala 32:86]
  wire [31:0] _io_out_T_30_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_30_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_30_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_30_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_30_rs3; // @[package.scala 32:76]
  wire  _io_out_T_31; // @[package.scala 32:86]
  wire [31:0] io_out_s_16_bits; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _io_out_T_32_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_32_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_32_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_32_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_32_rs3; // @[package.scala 32:76]
  wire  _io_out_T_33; // @[package.scala 32:86]
  wire [31:0] io_out_s_17_bits; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _io_out_T_34_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_34_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_34_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_34_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_34_rs3; // @[package.scala 32:76]
  wire  _io_out_T_35; // @[package.scala 32:86]
  wire [31:0] io_out_s_18_bits; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _io_out_T_36_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_36_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_36_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_36_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_36_rs3; // @[package.scala 32:76]
  wire  _io_out_T_37; // @[package.scala 32:86]
  wire [31:0] io_out_s_19_bits; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _io_out_T_38_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_38_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_38_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_38_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_38_rs3; // @[package.scala 32:76]
  wire  _io_out_T_39; // @[package.scala 32:86]
  wire [31:0] _io_out_T_40_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_40_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_40_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_40_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_40_rs3; // @[package.scala 32:76]
  wire  _io_out_T_41; // @[package.scala 32:86]
  wire [31:0] io_out_s_21_bits; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _io_out_T_42_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_42_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_42_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_42_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_42_rs3; // @[package.scala 32:76]
  wire  _io_out_T_43; // @[package.scala 32:86]
  wire [31:0] io_out_s_22_bits; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _io_out_T_44_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_44_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_44_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_44_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_44_rs3; // @[package.scala 32:76]
  wire  _io_out_T_45; // @[package.scala 32:86]
  wire [31:0] io_out_s_23_bits; // @[RVC.scala 21:19 RVC.scala 22:14]
  wire [31:0] _io_out_T_46_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_46_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_46_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_46_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_46_rs3; // @[package.scala 32:76]
  wire  _io_out_T_47; // @[package.scala 32:86]
  wire [31:0] _io_out_T_48_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_48_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_48_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_48_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_48_rs3; // @[package.scala 32:76]
  wire  _io_out_T_49; // @[package.scala 32:86]
  wire [31:0] _io_out_T_50_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_50_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_50_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_50_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_50_rs3; // @[package.scala 32:76]
  wire  _io_out_T_51; // @[package.scala 32:86]
  wire [31:0] _io_out_T_52_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_52_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_52_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_52_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_52_rs3; // @[package.scala 32:76]
  wire  _io_out_T_53; // @[package.scala 32:86]
  wire [31:0] _io_out_T_54_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_54_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_54_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_54_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_54_rs3; // @[package.scala 32:76]
  wire  _io_out_T_55; // @[package.scala 32:86]
  wire [31:0] _io_out_T_56_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_56_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_56_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_56_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_56_rs3; // @[package.scala 32:76]
  wire  _io_out_T_57; // @[package.scala 32:86]
  wire [31:0] _io_out_T_58_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_58_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_58_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_58_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_58_rs3; // @[package.scala 32:76]
  wire  _io_out_T_59; // @[package.scala 32:86]
  wire [31:0] _io_out_T_60_bits; // @[package.scala 32:76]
  wire [4:0] _io_out_T_60_rd; // @[package.scala 32:76]
  wire [4:0] _io_out_T_60_rs1; // @[package.scala 32:76]
  wire [4:0] _io_out_T_60_rs2; // @[package.scala 32:76]
  wire [4:0] _io_out_T_60_rs3; // @[package.scala 32:76]
  wire  _io_out_T_61; // @[package.scala 32:86]
  wire [29:0] RVCExpander_covSum;
  assign _io_out_s_opc_T_1 = |io_in[12:5]; // @[RVC.scala 53:29]
  assign io_out_s_lo_lo = _io_out_s_opc_T_1 ? 7'h13 : 7'h1f; // @[RVC.scala 53:20]
  assign io_out_s_hi_hi_hi = io_in[10:7]; // @[RVC.scala 34:26]
  assign io_out_s_hi_hi_lo = io_in[12:11]; // @[RVC.scala 34:35]
  assign io_out_s_hi_lo = io_in[5]; // @[RVC.scala 34:45]
  assign io_out_s_lo_hi = io_in[6]; // @[RVC.scala 34:51]
  assign io_out_s_lo_1 = io_in[4:2]; // @[RVC.scala 31:29]
  assign io_out_s_lo_hi_1 = {2'h1,io_out_s_lo_1}; // @[Cat.scala 30:58]
  assign _io_out_s_T = {io_out_s_hi_hi_hi,io_out_s_hi_hi_lo,io_out_s_hi_lo,io_out_s_lo_hi,2'h0,5'h2,3'h0,2'h1,io_out_s_lo_1,io_out_s_lo_lo}; // @[Cat.scala 30:58]
  assign io_out_s_0_rs3 = io_in[31:27]; // @[RVC.scala 20:101]
  assign io_out_s_hi_hi_2 = io_in[6:5]; // @[RVC.scala 36:20]
  assign io_out_s_hi_lo_1 = io_in[12:10]; // @[RVC.scala 36:28]
  assign io_out_s_hi_hi_hi_2 = {io_out_s_hi_hi_2,io_out_s_hi_lo_1,3'h0}; // @[Cat.scala 30:58]
  assign io_out_s_lo_5 = io_in[9:7]; // @[RVC.scala 30:29]
  assign io_out_s_hi_hi_lo_1 = {2'h1,io_out_s_lo_5}; // @[Cat.scala 30:58]
  assign _io_out_s_T_4 = {io_out_s_hi_hi_2,io_out_s_hi_lo_1,3'h0,2'h1,io_out_s_lo_5,3'h3,2'h1,io_out_s_lo_1,7'h7}; // @[Cat.scala 30:58]
  assign io_out_s_hi_hi_hi_3 = {io_out_s_hi_lo,io_out_s_hi_lo_1,io_out_s_lo_hi,2'h0}; // @[Cat.scala 30:58]
  assign _io_out_s_T_9 = {io_out_s_hi_lo,io_out_s_hi_lo_1,io_out_s_lo_hi,2'h0,2'h1,io_out_s_lo_5,3'h2,2'h1,io_out_s_lo_1,7'h3}; // @[Cat.scala 30:58]
  assign _io_out_s_T_14 = {io_out_s_hi_hi_2,io_out_s_hi_lo_1,3'h0,2'h1,io_out_s_lo_5,3'h3,2'h1,io_out_s_lo_1,7'h3}; // @[Cat.scala 30:58]
  assign io_out_s_hi_hi_hi_5 = io_out_s_hi_hi_hi_3[6:5]; // @[RVC.scala 63:32]
  assign io_out_s_lo_hi_lo = io_out_s_hi_hi_hi_3[4:0]; // @[RVC.scala 63:65]
  assign _io_out_s_T_21 = {io_out_s_hi_hi_hi_5,2'h1,io_out_s_lo_1,2'h1,io_out_s_lo_5,3'h2,io_out_s_lo_hi_lo,7'h3f}; // @[Cat.scala 30:58]
  assign io_out_s_hi_hi_hi_6 = io_out_s_hi_hi_hi_2[7:5]; // @[RVC.scala 66:30]
  assign io_out_s_lo_hi_lo_1 = io_out_s_hi_hi_hi_2[4:0]; // @[RVC.scala 66:63]
  assign _io_out_s_T_28 = {io_out_s_hi_hi_hi_6,2'h1,io_out_s_lo_1,2'h1,io_out_s_lo_5,3'h3,io_out_s_lo_hi_lo_1,7'h27}; // @[Cat.scala 30:58]
  assign _io_out_s_T_35 = {io_out_s_hi_hi_hi_5,2'h1,io_out_s_lo_1,2'h1,io_out_s_lo_5,3'h2,io_out_s_lo_hi_lo,7'h23}; // @[Cat.scala 30:58]
  assign _io_out_s_T_42 = {io_out_s_hi_hi_hi_6,2'h1,io_out_s_lo_1,2'h1,io_out_s_lo_5,3'h3,io_out_s_lo_hi_lo_1,7'h23}; // @[Cat.scala 30:58]
  assign io_out_s_hi_20 = io_in[12] ? 7'h7f : 7'h0; // @[Bitwise.scala 72:12]
  assign io_out_s_lo_52 = io_in[6:2]; // @[RVC.scala 43:38]
  assign io_out_s_hi_hi_hi_9 = {io_out_s_hi_20,io_out_s_lo_52}; // @[Cat.scala 30:58]
  assign io_out_s_hi_hi_lo_8 = io_in[11:7]; // @[RVC.scala 33:13]
  assign io_out_s_8_bits = {io_out_s_hi_20,io_out_s_lo_52,io_out_s_hi_hi_lo_8,3'h0,io_out_s_hi_hi_lo_8,7'h13}; // @[Cat.scala 30:58]
  assign _io_out_s_opc_T_3 = |io_out_s_hi_hi_lo_8; // @[RVC.scala 77:24]
  assign io_out_s_lo_lo_1 = _io_out_s_opc_T_3 ? 7'h1b : 7'h1f; // @[RVC.scala 77:20]
  assign io_out_s_9_bits = {io_out_s_hi_20,io_out_s_lo_52,io_out_s_hi_hi_lo_8,3'h0,io_out_s_hi_hi_lo_8,io_out_s_lo_lo_1}; // @[Cat.scala 30:58]
  assign io_out_s_10_bits = {io_out_s_hi_20,io_out_s_lo_52,5'h0,3'h0,io_out_s_hi_hi_lo_8,7'h13}; // @[Cat.scala 30:58]
  assign _io_out_s_opc_T_7 = |io_out_s_hi_hi_hi_9; // @[RVC.scala 90:29]
  assign io_out_s_me_lo = _io_out_s_opc_T_7 ? 7'h37 : 7'h3f; // @[RVC.scala 90:20]
  assign io_out_s_me_hi_hi = io_in[12] ? 15'h7fff : 15'h0; // @[Bitwise.scala 72:12]
  assign _io_out_s_me_T_2 = {io_out_s_me_hi_hi,io_out_s_lo_52,12'h0}; // @[Cat.scala 30:58]
  assign io_out_s_me_hi_hi_1 = _io_out_s_me_T_2[31:12]; // @[RVC.scala 91:31]
  assign io_out_s_me_bits = {io_out_s_me_hi_hi_1,io_out_s_hi_hi_lo_8,io_out_s_me_lo}; // @[Cat.scala 30:58]
  assign _io_out_s_T_68 = io_out_s_hi_hi_lo_8 == 5'h0; // @[RVC.scala 92:14]
  assign _io_out_s_T_70 = io_out_s_hi_hi_lo_8 == 5'h2; // @[RVC.scala 92:27]
  assign _io_out_s_T_71 = _io_out_s_T_68 | _io_out_s_T_70; // @[RVC.scala 92:21]
  assign io_out_s_lo_lo_2 = _io_out_s_opc_T_7 ? 7'h13 : 7'h1f; // @[RVC.scala 86:20]
  assign io_out_s_hi_hi_hi_12 = io_in[12] ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  assign io_out_s_hi_hi_lo_10 = io_in[4:3]; // @[RVC.scala 42:42]
  assign io_out_s_lo_hi_hi = io_in[2]; // @[RVC.scala 42:56]
  assign io_out_s_res_bits = {io_out_s_hi_hi_hi_12,io_out_s_hi_hi_lo_10,io_out_s_hi_lo,io_out_s_lo_hi_hi,io_out_s_lo_hi,4'h0,io_out_s_hi_hi_lo_8,3'h0,io_out_s_hi_hi_lo_8,io_out_s_lo_lo_2}; // @[Cat.scala 30:58]
  assign io_out_s_11_bits = _io_out_s_T_71 ? io_out_s_res_bits : io_out_s_me_bits; // @[RVC.scala 92:10]
  assign io_out_s_11_rd = _io_out_s_T_71 ? io_out_s_hi_hi_lo_8 : io_out_s_hi_hi_lo_8; // @[RVC.scala 92:10]
  assign io_out_s_11_rs2 = _io_out_s_T_71 ? io_out_s_lo_hi_1 : io_out_s_lo_hi_1; // @[RVC.scala 92:10]
  assign io_out_s_11_rs3 = _io_out_s_T_71 ? io_out_s_0_rs3 : io_out_s_0_rs3; // @[RVC.scala 92:10]
  assign _io_out_s_T_79 = {io_in[12],io_out_s_lo_52,2'h1,io_out_s_lo_5,3'h5,2'h1,io_out_s_lo_5,7'h13}; // @[Cat.scala 30:58]
  assign _GEN_0 = {{5'd0}, _io_out_s_T_79}; // @[RVC.scala 99:23]
  assign _io_out_s_T_81 = _GEN_0 | 31'h40000000; // @[RVC.scala 99:23]
  assign _io_out_s_T_84 = {io_out_s_hi_20,io_out_s_lo_52,2'h1,io_out_s_lo_5,3'h7,2'h1,io_out_s_lo_5,7'h13}; // @[Cat.scala 30:58]
  assign _io_out_s_funct_T = {io_in[12],io_out_s_hi_hi_2}; // @[Cat.scala 30:58]
  assign _io_out_s_funct_T_1 = _io_out_s_funct_T == 3'h1; // @[package.scala 32:86]
  assign _io_out_s_funct_T_2 = _io_out_s_funct_T_1 ? 3'h4 : 3'h0; // @[package.scala 32:76]
  assign _io_out_s_funct_T_3 = _io_out_s_funct_T == 3'h2; // @[package.scala 32:86]
  assign _io_out_s_funct_T_4 = _io_out_s_funct_T_3 ? 3'h6 : _io_out_s_funct_T_2; // @[package.scala 32:76]
  assign _io_out_s_funct_T_5 = _io_out_s_funct_T == 3'h3; // @[package.scala 32:86]
  assign _io_out_s_funct_T_6 = _io_out_s_funct_T_5 ? 3'h7 : _io_out_s_funct_T_4; // @[package.scala 32:76]
  assign _io_out_s_funct_T_7 = _io_out_s_funct_T == 3'h4; // @[package.scala 32:86]
  assign _io_out_s_funct_T_8 = _io_out_s_funct_T_7 ? 3'h0 : _io_out_s_funct_T_6; // @[package.scala 32:76]
  assign _io_out_s_funct_T_9 = _io_out_s_funct_T == 3'h5; // @[package.scala 32:86]
  assign _io_out_s_funct_T_10 = _io_out_s_funct_T_9 ? 3'h0 : _io_out_s_funct_T_8; // @[package.scala 32:76]
  assign _io_out_s_funct_T_11 = _io_out_s_funct_T == 3'h6; // @[package.scala 32:86]
  assign _io_out_s_funct_T_12 = _io_out_s_funct_T_11 ? 3'h2 : _io_out_s_funct_T_10; // @[package.scala 32:76]
  assign _io_out_s_funct_T_13 = _io_out_s_funct_T == 3'h7; // @[package.scala 32:86]
  assign io_out_s_hi_lo_17 = _io_out_s_funct_T_13 ? 3'h3 : _io_out_s_funct_T_12; // @[package.scala 32:76]
  assign _io_out_s_sub_T_1 = io_out_s_hi_hi_2 == 2'h0; // @[RVC.scala 103:30]
  assign io_out_s_sub = _io_out_s_sub_T_1 ? 31'h40000000 : 31'h0; // @[RVC.scala 103:22]
  assign io_out_s_lo_lo_3 = io_in[12] ? 7'h3b : 7'h33; // @[RVC.scala 104:22]
  assign _io_out_s_T_85 = {2'h1,io_out_s_lo_1,2'h1,io_out_s_lo_5,io_out_s_hi_lo_17,2'h1,io_out_s_lo_5,io_out_s_lo_lo_3}; // @[Cat.scala 30:58]
  assign _GEN_1 = {{6'd0}, _io_out_s_T_85}; // @[RVC.scala 105:43]
  assign _io_out_s_T_86 = _GEN_1 | io_out_s_sub; // @[RVC.scala 105:43]
  assign _io_out_s_T_88 = io_in[11:10] == 2'h1; // @[package.scala 32:86]
  assign _io_out_s_T_89 = _io_out_s_T_88 ? _io_out_s_T_81 : {{5'd0}, _io_out_s_T_79}; // @[package.scala 32:76]
  assign _io_out_s_T_90 = io_in[11:10] == 2'h2; // @[package.scala 32:86]
  assign _io_out_s_T_91 = _io_out_s_T_90 ? _io_out_s_T_84 : {{1'd0}, _io_out_s_T_89}; // @[package.scala 32:76]
  assign _io_out_s_T_92 = io_in[11:10] == 2'h3; // @[package.scala 32:86]
  assign io_out_s_12_bits = _io_out_s_T_92 ? {{1'd0}, _io_out_s_T_86} : _io_out_s_T_91; // @[package.scala 32:76]
  assign io_out_s_hi_hi_hi_hi = io_in[12] ? 10'h3ff : 10'h0; // @[Bitwise.scala 72:12]
  assign io_out_s_hi_hi_hi_lo = io_in[8]; // @[RVC.scala 44:36]
  assign io_out_s_hi_hi_lo_16 = io_in[10:9]; // @[RVC.scala 44:42]
  assign io_out_s_hi_lo_lo = io_in[7]; // @[RVC.scala 44:57]
  assign io_out_s_lo_hi_lo_5 = io_in[11]; // @[RVC.scala 44:69]
  assign io_out_s_lo_lo_hi = io_in[5:3]; // @[RVC.scala 44:76]
  assign _io_out_s_T_100 = {io_out_s_hi_hi_hi_hi,io_out_s_hi_hi_hi_lo,io_out_s_hi_hi_lo_16,io_out_s_lo_hi,io_out_s_hi_lo_lo,io_out_s_lo_hi_hi,io_out_s_lo_hi_lo_5,io_out_s_lo_lo_hi,1'h0}; // @[Cat.scala 30:58]
  assign io_out_s_hi_hi_hi_19 = _io_out_s_T_100[20]; // @[RVC.scala 94:26]
  assign io_out_s_hi_hi_lo_18 = _io_out_s_T_100[10:1]; // @[RVC.scala 94:36]
  assign io_out_s_hi_lo_21 = _io_out_s_T_100[11]; // @[RVC.scala 94:48]
  assign io_out_s_lo_hi_hi_5 = _io_out_s_T_100[19:12]; // @[RVC.scala 94:58]
  assign io_out_s_13_bits = {io_out_s_hi_hi_hi_19,io_out_s_hi_hi_lo_18,io_out_s_hi_lo_21,io_out_s_lo_hi_hi_5,5'h0,7'h6f}; // @[Cat.scala 30:58]
  assign io_out_s_hi_hi_hi_23 = io_in[12] ? 5'h1f : 5'h0; // @[Bitwise.scala 72:12]
  assign _io_out_s_T_116 = {io_out_s_hi_hi_hi_23,io_out_s_hi_hi_2,io_out_s_lo_hi_hi,io_in[11:10],io_out_s_hi_hi_lo_10,1'h0}; // @[Cat.scala 30:58]
  assign io_out_s_hi_hi_hi_24 = _io_out_s_T_116[12]; // @[RVC.scala 95:29]
  assign io_out_s_hi_hi_lo_23 = _io_out_s_T_116[10:5]; // @[RVC.scala 95:39]
  assign io_out_s_lo_hi_lo_12 = _io_out_s_T_116[4:1]; // @[RVC.scala 95:71]
  assign io_out_s_lo_lo_hi_4 = _io_out_s_T_116[11]; // @[RVC.scala 95:82]
  assign io_out_s_14_bits = {io_out_s_hi_hi_hi_24,io_out_s_hi_hi_lo_23,5'h0,2'h1,io_out_s_lo_5,3'h0,io_out_s_lo_hi_lo_12,io_out_s_lo_lo_hi_4,7'h63}; // @[Cat.scala 30:58]
  assign io_out_s_15_bits = {io_out_s_hi_hi_hi_24,io_out_s_hi_hi_lo_23,5'h0,2'h1,io_out_s_lo_5,3'h1,io_out_s_lo_hi_lo_12,io_out_s_lo_lo_hi_4,7'h63}; // @[Cat.scala 30:58]
  assign io_out_s_lo_lo_10 = _io_out_s_opc_T_3 ? 7'h3 : 7'h1f; // @[RVC.scala 113:23]
  assign _io_out_s_T_145 = {io_in[12],io_out_s_lo_52,io_out_s_hi_hi_lo_8,3'h1,io_out_s_hi_hi_lo_8,7'h13}; // @[Cat.scala 30:58]
  assign _io_out_s_T_150 = {io_out_s_lo_1,io_in[12],io_out_s_hi_hi_2,3'h0,5'h2,3'h3,io_out_s_hi_hi_lo_8,7'h7}; // @[Cat.scala 30:58]
  assign io_out_s_hi_hi_47 = io_in[3:2]; // @[RVC.scala 37:22]
  assign io_out_s_lo_hi_41 = io_in[6:4]; // @[RVC.scala 37:37]
  assign _io_out_s_T_154 = {io_out_s_hi_hi_47,io_in[12],io_out_s_lo_hi_41,2'h0,5'h2,3'h2,io_out_s_hi_hi_lo_8,io_out_s_lo_lo_10}; // @[Cat.scala 30:58]
  assign _io_out_s_T_158 = {io_out_s_lo_1,io_in[12],io_out_s_hi_hi_2,3'h0,5'h2,3'h3,io_out_s_hi_hi_lo_8,io_out_s_lo_lo_10}; // @[Cat.scala 30:58]
  assign _io_out_s_mv_T = {io_out_s_lo_52,5'h0,3'h0,io_out_s_hi_hi_lo_8,7'h33}; // @[Cat.scala 30:58]
  assign _io_out_s_add_T = {io_out_s_lo_52,io_out_s_hi_hi_lo_8,3'h0,io_out_s_hi_hi_lo_8,7'h33}; // @[Cat.scala 30:58]
  assign io_out_s_jr = {io_out_s_lo_52,io_out_s_hi_hi_lo_8,3'h0,12'h67}; // @[Cat.scala 30:58]
  assign io_out_s_reserved_hi = io_out_s_jr[24:7]; // @[RVC.scala 133:29]
  assign io_out_s_reserved = {io_out_s_reserved_hi,7'h1f}; // @[Cat.scala 30:58]
  assign _io_out_s_jr_reserved_T_2 = _io_out_s_opc_T_3 ? io_out_s_jr : io_out_s_reserved; // @[RVC.scala 134:33]
  assign _io_out_s_jr_mv_T_1 = |io_out_s_lo_52; // @[RVC.scala 135:27]
  assign io_out_s_mv_bits = {{7'd0}, _io_out_s_mv_T}; // @[RVC.scala 21:19 RVC.scala 22:14]
  assign io_out_s_jr_reserved_bits = {{7'd0}, _io_out_s_jr_reserved_T_2}; // @[RVC.scala 21:19 RVC.scala 22:14]
  assign io_out_s_jr_mv_bits = _io_out_s_jr_mv_T_1 ? io_out_s_mv_bits : io_out_s_jr_reserved_bits; // @[RVC.scala 135:22]
  assign io_out_s_jr_mv_rd = _io_out_s_jr_mv_T_1 ? io_out_s_hi_hi_lo_8 : 5'h0; // @[RVC.scala 135:22]
  assign io_out_s_jr_mv_rs1 = _io_out_s_jr_mv_T_1 ? 5'h0 : io_out_s_hi_hi_lo_8; // @[RVC.scala 135:22]
  assign io_out_s_jr_mv_rs2 = _io_out_s_jr_mv_T_1 ? io_out_s_lo_52 : io_out_s_lo_52; // @[RVC.scala 135:22]
  assign io_out_s_jr_mv_rs3 = _io_out_s_jr_mv_T_1 ? io_out_s_0_rs3 : io_out_s_0_rs3; // @[RVC.scala 135:22]
  assign io_out_s_jalr = {io_out_s_lo_52,io_out_s_hi_hi_lo_8,3'h0,12'he7}; // @[Cat.scala 30:58]
  assign _io_out_s_ebreak_T = {io_out_s_reserved_hi,7'h73}; // @[Cat.scala 30:58]
  assign io_out_s_ebreak = _io_out_s_ebreak_T | 25'h100000; // @[RVC.scala 137:46]
  assign _io_out_s_jalr_ebreak_T_2 = _io_out_s_opc_T_3 ? io_out_s_jalr : io_out_s_ebreak; // @[RVC.scala 138:33]
  assign io_out_s_add_bits = {{7'd0}, _io_out_s_add_T}; // @[RVC.scala 21:19 RVC.scala 22:14]
  assign io_out_s_jalr_ebreak_bits = {{7'd0}, _io_out_s_jalr_ebreak_T_2}; // @[RVC.scala 21:19 RVC.scala 22:14]
  assign io_out_s_jalr_add_bits = _io_out_s_jr_mv_T_1 ? io_out_s_add_bits : io_out_s_jalr_ebreak_bits; // @[RVC.scala 139:25]
  assign io_out_s_jalr_add_rd = _io_out_s_jr_mv_T_1 ? io_out_s_hi_hi_lo_8 : 5'h1; // @[RVC.scala 139:25]
  assign io_out_s_jalr_add_rs1 = _io_out_s_jr_mv_T_1 ? io_out_s_hi_hi_lo_8 : io_out_s_hi_hi_lo_8; // @[RVC.scala 139:25]
  assign io_out_s_20_bits = io_in[12] ? io_out_s_jalr_add_bits : io_out_s_jr_mv_bits; // @[RVC.scala 140:10]
  assign io_out_s_20_rd = io_in[12] ? io_out_s_jalr_add_rd : io_out_s_jr_mv_rd; // @[RVC.scala 140:10]
  assign io_out_s_20_rs1 = io_in[12] ? io_out_s_jalr_add_rs1 : io_out_s_jr_mv_rs1; // @[RVC.scala 140:10]
  assign io_out_s_20_rs2 = io_in[12] ? io_out_s_jr_mv_rs2 : io_out_s_jr_mv_rs2; // @[RVC.scala 140:10]
  assign io_out_s_20_rs3 = io_in[12] ? io_out_s_jr_mv_rs3 : io_out_s_jr_mv_rs3; // @[RVC.scala 140:10]
  assign _io_out_s_T_163 = {io_out_s_lo_5,io_out_s_hi_lo_1,3'h0}; // @[Cat.scala 30:58]
  assign io_out_s_hi_hi_hi_37 = _io_out_s_T_163[8:5]; // @[RVC.scala 124:34]
  assign io_out_s_lo_hi_lo_19 = _io_out_s_T_163[4:0]; // @[RVC.scala 124:66]
  assign _io_out_s_T_165 = {io_out_s_hi_hi_hi_37,io_out_s_lo_52,5'h2,3'h3,io_out_s_lo_hi_lo_19,7'h27}; // @[Cat.scala 30:58]
  assign io_out_s_hi_hi_54 = io_in[8:7]; // @[RVC.scala 39:22]
  assign io_out_s_hi_lo_38 = io_in[12:9]; // @[RVC.scala 39:30]
  assign _io_out_s_T_169 = {io_out_s_hi_hi_54,io_out_s_hi_lo_38,2'h0}; // @[Cat.scala 30:58]
  assign io_out_s_hi_hi_hi_38 = _io_out_s_T_169[7:5]; // @[RVC.scala 123:33]
  assign io_out_s_lo_hi_lo_20 = _io_out_s_T_169[4:0]; // @[RVC.scala 123:65]
  assign _io_out_s_T_171 = {io_out_s_hi_hi_hi_38,io_out_s_lo_52,5'h2,3'h2,io_out_s_lo_hi_lo_20,7'h23}; // @[Cat.scala 30:58]
  assign _io_out_s_T_177 = {io_out_s_hi_hi_hi_37,io_out_s_lo_52,5'h2,3'h3,io_out_s_lo_hi_lo_19,7'h23}; // @[Cat.scala 30:58]
  assign io_out_s_24_rs1 = io_in[19:15]; // @[RVC.scala 20:57]
  assign io_out_s_24_rs2 = io_in[24:20]; // @[RVC.scala 20:79]
  assign io_out_lo = io_in[15:13]; // @[RVC.scala 151:20]
  assign _io_out_T = {io_in[1:0],io_out_lo}; // @[Cat.scala 30:58]
  assign _io_out_T_1 = _io_out_T == 5'h1; // @[package.scala 32:86]
  assign io_out_s_1_bits = {{4'd0}, _io_out_s_T_4}; // @[RVC.scala 21:19 RVC.scala 22:14]
  assign io_out_s_0_bits = {{2'd0}, _io_out_s_T}; // @[RVC.scala 21:19 RVC.scala 22:14]
  assign _io_out_T_2_bits = _io_out_T_1 ? io_out_s_1_bits : io_out_s_0_bits; // @[package.scala 32:76]
  assign _io_out_T_2_rd = _io_out_T_1 ? io_out_s_lo_hi_1 : io_out_s_lo_hi_1; // @[package.scala 32:76]
  assign _io_out_T_2_rs1 = _io_out_T_1 ? io_out_s_hi_hi_lo_1 : 5'h2; // @[package.scala 32:76]
  assign _io_out_T_2_rs3 = _io_out_T_1 ? io_out_s_0_rs3 : io_out_s_0_rs3; // @[package.scala 32:76]
  assign _io_out_T_3 = _io_out_T == 5'h2; // @[package.scala 32:86]
  assign io_out_s_2_bits = {{5'd0}, _io_out_s_T_9}; // @[RVC.scala 21:19 RVC.scala 22:14]
  assign _io_out_T_4_bits = _io_out_T_3 ? io_out_s_2_bits : _io_out_T_2_bits; // @[package.scala 32:76]
  assign _io_out_T_4_rd = _io_out_T_3 ? io_out_s_lo_hi_1 : _io_out_T_2_rd; // @[package.scala 32:76]
  assign _io_out_T_4_rs1 = _io_out_T_3 ? io_out_s_hi_hi_lo_1 : _io_out_T_2_rs1; // @[package.scala 32:76]
  assign _io_out_T_4_rs3 = _io_out_T_3 ? io_out_s_0_rs3 : _io_out_T_2_rs3; // @[package.scala 32:76]
  assign _io_out_T_5 = _io_out_T == 5'h3; // @[package.scala 32:86]
  assign io_out_s_3_bits = {{4'd0}, _io_out_s_T_14}; // @[RVC.scala 21:19 RVC.scala 22:14]
  assign _io_out_T_6_bits = _io_out_T_5 ? io_out_s_3_bits : _io_out_T_4_bits; // @[package.scala 32:76]
  assign _io_out_T_6_rd = _io_out_T_5 ? io_out_s_lo_hi_1 : _io_out_T_4_rd; // @[package.scala 32:76]
  assign _io_out_T_6_rs1 = _io_out_T_5 ? io_out_s_hi_hi_lo_1 : _io_out_T_4_rs1; // @[package.scala 32:76]
  assign _io_out_T_6_rs3 = _io_out_T_5 ? io_out_s_0_rs3 : _io_out_T_4_rs3; // @[package.scala 32:76]
  assign _io_out_T_7 = _io_out_T == 5'h4; // @[package.scala 32:86]
  assign io_out_s_4_bits = {{5'd0}, _io_out_s_T_21}; // @[RVC.scala 21:19 RVC.scala 22:14]
  assign _io_out_T_8_bits = _io_out_T_7 ? io_out_s_4_bits : _io_out_T_6_bits; // @[package.scala 32:76]
  assign _io_out_T_8_rd = _io_out_T_7 ? io_out_s_lo_hi_1 : _io_out_T_6_rd; // @[package.scala 32:76]
  assign _io_out_T_8_rs1 = _io_out_T_7 ? io_out_s_hi_hi_lo_1 : _io_out_T_6_rs1; // @[package.scala 32:76]
  assign _io_out_T_8_rs3 = _io_out_T_7 ? io_out_s_0_rs3 : _io_out_T_6_rs3; // @[package.scala 32:76]
  assign _io_out_T_9 = _io_out_T == 5'h5; // @[package.scala 32:86]
  assign io_out_s_5_bits = {{4'd0}, _io_out_s_T_28}; // @[RVC.scala 21:19 RVC.scala 22:14]
  assign _io_out_T_10_bits = _io_out_T_9 ? io_out_s_5_bits : _io_out_T_8_bits; // @[package.scala 32:76]
  assign _io_out_T_10_rd = _io_out_T_9 ? io_out_s_lo_hi_1 : _io_out_T_8_rd; // @[package.scala 32:76]
  assign _io_out_T_10_rs1 = _io_out_T_9 ? io_out_s_hi_hi_lo_1 : _io_out_T_8_rs1; // @[package.scala 32:76]
  assign _io_out_T_10_rs3 = _io_out_T_9 ? io_out_s_0_rs3 : _io_out_T_8_rs3; // @[package.scala 32:76]
  assign _io_out_T_11 = _io_out_T == 5'h6; // @[package.scala 32:86]
  assign io_out_s_6_bits = {{5'd0}, _io_out_s_T_35}; // @[RVC.scala 21:19 RVC.scala 22:14]
  assign _io_out_T_12_bits = _io_out_T_11 ? io_out_s_6_bits : _io_out_T_10_bits; // @[package.scala 32:76]
  assign _io_out_T_12_rd = _io_out_T_11 ? io_out_s_lo_hi_1 : _io_out_T_10_rd; // @[package.scala 32:76]
  assign _io_out_T_12_rs1 = _io_out_T_11 ? io_out_s_hi_hi_lo_1 : _io_out_T_10_rs1; // @[package.scala 32:76]
  assign _io_out_T_12_rs3 = _io_out_T_11 ? io_out_s_0_rs3 : _io_out_T_10_rs3; // @[package.scala 32:76]
  assign _io_out_T_13 = _io_out_T == 5'h7; // @[package.scala 32:86]
  assign io_out_s_7_bits = {{4'd0}, _io_out_s_T_42}; // @[RVC.scala 21:19 RVC.scala 22:14]
  assign _io_out_T_14_bits = _io_out_T_13 ? io_out_s_7_bits : _io_out_T_12_bits; // @[package.scala 32:76]
  assign _io_out_T_14_rd = _io_out_T_13 ? io_out_s_lo_hi_1 : _io_out_T_12_rd; // @[package.scala 32:76]
  assign _io_out_T_14_rs1 = _io_out_T_13 ? io_out_s_hi_hi_lo_1 : _io_out_T_12_rs1; // @[package.scala 32:76]
  assign _io_out_T_14_rs3 = _io_out_T_13 ? io_out_s_0_rs3 : _io_out_T_12_rs3; // @[package.scala 32:76]
  assign _io_out_T_15 = _io_out_T == 5'h8; // @[package.scala 32:86]
  assign _io_out_T_16_bits = _io_out_T_15 ? io_out_s_8_bits : _io_out_T_14_bits; // @[package.scala 32:76]
  assign _io_out_T_16_rd = _io_out_T_15 ? io_out_s_hi_hi_lo_8 : _io_out_T_14_rd; // @[package.scala 32:76]
  assign _io_out_T_16_rs1 = _io_out_T_15 ? io_out_s_hi_hi_lo_8 : _io_out_T_14_rs1; // @[package.scala 32:76]
  assign _io_out_T_16_rs2 = _io_out_T_15 ? io_out_s_lo_hi_1 : _io_out_T_14_rd; // @[package.scala 32:76]
  assign _io_out_T_16_rs3 = _io_out_T_15 ? io_out_s_0_rs3 : _io_out_T_14_rs3; // @[package.scala 32:76]
  assign _io_out_T_17 = _io_out_T == 5'h9; // @[package.scala 32:86]
  assign _io_out_T_18_bits = _io_out_T_17 ? io_out_s_9_bits : _io_out_T_16_bits; // @[package.scala 32:76]
  assign _io_out_T_18_rd = _io_out_T_17 ? io_out_s_hi_hi_lo_8 : _io_out_T_16_rd; // @[package.scala 32:76]
  assign _io_out_T_18_rs1 = _io_out_T_17 ? io_out_s_hi_hi_lo_8 : _io_out_T_16_rs1; // @[package.scala 32:76]
  assign _io_out_T_18_rs2 = _io_out_T_17 ? io_out_s_lo_hi_1 : _io_out_T_16_rs2; // @[package.scala 32:76]
  assign _io_out_T_18_rs3 = _io_out_T_17 ? io_out_s_0_rs3 : _io_out_T_16_rs3; // @[package.scala 32:76]
  assign _io_out_T_19 = _io_out_T == 5'ha; // @[package.scala 32:86]
  assign _io_out_T_20_bits = _io_out_T_19 ? io_out_s_10_bits : _io_out_T_18_bits; // @[package.scala 32:76]
  assign _io_out_T_20_rd = _io_out_T_19 ? io_out_s_hi_hi_lo_8 : _io_out_T_18_rd; // @[package.scala 32:76]
  assign _io_out_T_20_rs1 = _io_out_T_19 ? 5'h0 : _io_out_T_18_rs1; // @[package.scala 32:76]
  assign _io_out_T_20_rs2 = _io_out_T_19 ? io_out_s_lo_hi_1 : _io_out_T_18_rs2; // @[package.scala 32:76]
  assign _io_out_T_20_rs3 = _io_out_T_19 ? io_out_s_0_rs3 : _io_out_T_18_rs3; // @[package.scala 32:76]
  assign _io_out_T_21 = _io_out_T == 5'hb; // @[package.scala 32:86]
  assign _io_out_T_22_bits = _io_out_T_21 ? io_out_s_11_bits : _io_out_T_20_bits; // @[package.scala 32:76]
  assign _io_out_T_22_rd = _io_out_T_21 ? io_out_s_11_rd : _io_out_T_20_rd; // @[package.scala 32:76]
  assign _io_out_T_22_rs1 = _io_out_T_21 ? io_out_s_11_rd : _io_out_T_20_rs1; // @[package.scala 32:76]
  assign _io_out_T_22_rs2 = _io_out_T_21 ? io_out_s_11_rs2 : _io_out_T_20_rs2; // @[package.scala 32:76]
  assign _io_out_T_22_rs3 = _io_out_T_21 ? io_out_s_11_rs3 : _io_out_T_20_rs3; // @[package.scala 32:76]
  assign _io_out_T_23 = _io_out_T == 5'hc; // @[package.scala 32:86]
  assign _io_out_T_24_bits = _io_out_T_23 ? io_out_s_12_bits : _io_out_T_22_bits; // @[package.scala 32:76]
  assign _io_out_T_24_rd = _io_out_T_23 ? io_out_s_hi_hi_lo_1 : _io_out_T_22_rd; // @[package.scala 32:76]
  assign _io_out_T_24_rs1 = _io_out_T_23 ? io_out_s_hi_hi_lo_1 : _io_out_T_22_rs1; // @[package.scala 32:76]
  assign _io_out_T_24_rs2 = _io_out_T_23 ? io_out_s_lo_hi_1 : _io_out_T_22_rs2; // @[package.scala 32:76]
  assign _io_out_T_24_rs3 = _io_out_T_23 ? io_out_s_0_rs3 : _io_out_T_22_rs3; // @[package.scala 32:76]
  assign _io_out_T_25 = _io_out_T == 5'hd; // @[package.scala 32:86]
  assign _io_out_T_26_bits = _io_out_T_25 ? io_out_s_13_bits : _io_out_T_24_bits; // @[package.scala 32:76]
  assign _io_out_T_26_rd = _io_out_T_25 ? 5'h0 : _io_out_T_24_rd; // @[package.scala 32:76]
  assign _io_out_T_26_rs1 = _io_out_T_25 ? io_out_s_hi_hi_lo_1 : _io_out_T_24_rs1; // @[package.scala 32:76]
  assign _io_out_T_26_rs2 = _io_out_T_25 ? io_out_s_lo_hi_1 : _io_out_T_24_rs2; // @[package.scala 32:76]
  assign _io_out_T_26_rs3 = _io_out_T_25 ? io_out_s_0_rs3 : _io_out_T_24_rs3; // @[package.scala 32:76]
  assign _io_out_T_27 = _io_out_T == 5'he; // @[package.scala 32:86]
  assign _io_out_T_28_bits = _io_out_T_27 ? io_out_s_14_bits : _io_out_T_26_bits; // @[package.scala 32:76]
  assign _io_out_T_28_rd = _io_out_T_27 ? io_out_s_hi_hi_lo_1 : _io_out_T_26_rd; // @[package.scala 32:76]
  assign _io_out_T_28_rs1 = _io_out_T_27 ? io_out_s_hi_hi_lo_1 : _io_out_T_26_rs1; // @[package.scala 32:76]
  assign _io_out_T_28_rs2 = _io_out_T_27 ? 5'h0 : _io_out_T_26_rs2; // @[package.scala 32:76]
  assign _io_out_T_28_rs3 = _io_out_T_27 ? io_out_s_0_rs3 : _io_out_T_26_rs3; // @[package.scala 32:76]
  assign _io_out_T_29 = _io_out_T == 5'hf; // @[package.scala 32:86]
  assign _io_out_T_30_bits = _io_out_T_29 ? io_out_s_15_bits : _io_out_T_28_bits; // @[package.scala 32:76]
  assign _io_out_T_30_rd = _io_out_T_29 ? 5'h0 : _io_out_T_28_rd; // @[package.scala 32:76]
  assign _io_out_T_30_rs1 = _io_out_T_29 ? io_out_s_hi_hi_lo_1 : _io_out_T_28_rs1; // @[package.scala 32:76]
  assign _io_out_T_30_rs2 = _io_out_T_29 ? 5'h0 : _io_out_T_28_rs2; // @[package.scala 32:76]
  assign _io_out_T_30_rs3 = _io_out_T_29 ? io_out_s_0_rs3 : _io_out_T_28_rs3; // @[package.scala 32:76]
  assign _io_out_T_31 = _io_out_T == 5'h10; // @[package.scala 32:86]
  assign io_out_s_16_bits = {{6'd0}, _io_out_s_T_145}; // @[RVC.scala 21:19 RVC.scala 22:14]
  assign _io_out_T_32_bits = _io_out_T_31 ? io_out_s_16_bits : _io_out_T_30_bits; // @[package.scala 32:76]
  assign _io_out_T_32_rd = _io_out_T_31 ? io_out_s_hi_hi_lo_8 : _io_out_T_30_rd; // @[package.scala 32:76]
  assign _io_out_T_32_rs1 = _io_out_T_31 ? io_out_s_hi_hi_lo_8 : _io_out_T_30_rs1; // @[package.scala 32:76]
  assign _io_out_T_32_rs2 = _io_out_T_31 ? io_out_s_lo_52 : _io_out_T_30_rs2; // @[package.scala 32:76]
  assign _io_out_T_32_rs3 = _io_out_T_31 ? io_out_s_0_rs3 : _io_out_T_30_rs3; // @[package.scala 32:76]
  assign _io_out_T_33 = _io_out_T == 5'h11; // @[package.scala 32:86]
  assign io_out_s_17_bits = {{3'd0}, _io_out_s_T_150}; // @[RVC.scala 21:19 RVC.scala 22:14]
  assign _io_out_T_34_bits = _io_out_T_33 ? io_out_s_17_bits : _io_out_T_32_bits; // @[package.scala 32:76]
  assign _io_out_T_34_rd = _io_out_T_33 ? io_out_s_hi_hi_lo_8 : _io_out_T_32_rd; // @[package.scala 32:76]
  assign _io_out_T_34_rs1 = _io_out_T_33 ? 5'h2 : _io_out_T_32_rs1; // @[package.scala 32:76]
  assign _io_out_T_34_rs2 = _io_out_T_33 ? io_out_s_lo_52 : _io_out_T_32_rs2; // @[package.scala 32:76]
  assign _io_out_T_34_rs3 = _io_out_T_33 ? io_out_s_0_rs3 : _io_out_T_32_rs3; // @[package.scala 32:76]
  assign _io_out_T_35 = _io_out_T == 5'h12; // @[package.scala 32:86]
  assign io_out_s_18_bits = {{4'd0}, _io_out_s_T_154}; // @[RVC.scala 21:19 RVC.scala 22:14]
  assign _io_out_T_36_bits = _io_out_T_35 ? io_out_s_18_bits : _io_out_T_34_bits; // @[package.scala 32:76]
  assign _io_out_T_36_rd = _io_out_T_35 ? io_out_s_hi_hi_lo_8 : _io_out_T_34_rd; // @[package.scala 32:76]
  assign _io_out_T_36_rs1 = _io_out_T_35 ? 5'h2 : _io_out_T_34_rs1; // @[package.scala 32:76]
  assign _io_out_T_36_rs2 = _io_out_T_35 ? io_out_s_lo_52 : _io_out_T_34_rs2; // @[package.scala 32:76]
  assign _io_out_T_36_rs3 = _io_out_T_35 ? io_out_s_0_rs3 : _io_out_T_34_rs3; // @[package.scala 32:76]
  assign _io_out_T_37 = _io_out_T == 5'h13; // @[package.scala 32:86]
  assign io_out_s_19_bits = {{3'd0}, _io_out_s_T_158}; // @[RVC.scala 21:19 RVC.scala 22:14]
  assign _io_out_T_38_bits = _io_out_T_37 ? io_out_s_19_bits : _io_out_T_36_bits; // @[package.scala 32:76]
  assign _io_out_T_38_rd = _io_out_T_37 ? io_out_s_hi_hi_lo_8 : _io_out_T_36_rd; // @[package.scala 32:76]
  assign _io_out_T_38_rs1 = _io_out_T_37 ? 5'h2 : _io_out_T_36_rs1; // @[package.scala 32:76]
  assign _io_out_T_38_rs2 = _io_out_T_37 ? io_out_s_lo_52 : _io_out_T_36_rs2; // @[package.scala 32:76]
  assign _io_out_T_38_rs3 = _io_out_T_37 ? io_out_s_0_rs3 : _io_out_T_36_rs3; // @[package.scala 32:76]
  assign _io_out_T_39 = _io_out_T == 5'h14; // @[package.scala 32:86]
  assign _io_out_T_40_bits = _io_out_T_39 ? io_out_s_20_bits : _io_out_T_38_bits; // @[package.scala 32:76]
  assign _io_out_T_40_rd = _io_out_T_39 ? io_out_s_20_rd : _io_out_T_38_rd; // @[package.scala 32:76]
  assign _io_out_T_40_rs1 = _io_out_T_39 ? io_out_s_20_rs1 : _io_out_T_38_rs1; // @[package.scala 32:76]
  assign _io_out_T_40_rs2 = _io_out_T_39 ? io_out_s_20_rs2 : _io_out_T_38_rs2; // @[package.scala 32:76]
  assign _io_out_T_40_rs3 = _io_out_T_39 ? io_out_s_20_rs3 : _io_out_T_38_rs3; // @[package.scala 32:76]
  assign _io_out_T_41 = _io_out_T == 5'h15; // @[package.scala 32:86]
  assign io_out_s_21_bits = {{3'd0}, _io_out_s_T_165}; // @[RVC.scala 21:19 RVC.scala 22:14]
  assign _io_out_T_42_bits = _io_out_T_41 ? io_out_s_21_bits : _io_out_T_40_bits; // @[package.scala 32:76]
  assign _io_out_T_42_rd = _io_out_T_41 ? io_out_s_hi_hi_lo_8 : _io_out_T_40_rd; // @[package.scala 32:76]
  assign _io_out_T_42_rs1 = _io_out_T_41 ? 5'h2 : _io_out_T_40_rs1; // @[package.scala 32:76]
  assign _io_out_T_42_rs2 = _io_out_T_41 ? io_out_s_lo_52 : _io_out_T_40_rs2; // @[package.scala 32:76]
  assign _io_out_T_42_rs3 = _io_out_T_41 ? io_out_s_0_rs3 : _io_out_T_40_rs3; // @[package.scala 32:76]
  assign _io_out_T_43 = _io_out_T == 5'h16; // @[package.scala 32:86]
  assign io_out_s_22_bits = {{4'd0}, _io_out_s_T_171}; // @[RVC.scala 21:19 RVC.scala 22:14]
  assign _io_out_T_44_bits = _io_out_T_43 ? io_out_s_22_bits : _io_out_T_42_bits; // @[package.scala 32:76]
  assign _io_out_T_44_rd = _io_out_T_43 ? io_out_s_hi_hi_lo_8 : _io_out_T_42_rd; // @[package.scala 32:76]
  assign _io_out_T_44_rs1 = _io_out_T_43 ? 5'h2 : _io_out_T_42_rs1; // @[package.scala 32:76]
  assign _io_out_T_44_rs2 = _io_out_T_43 ? io_out_s_lo_52 : _io_out_T_42_rs2; // @[package.scala 32:76]
  assign _io_out_T_44_rs3 = _io_out_T_43 ? io_out_s_0_rs3 : _io_out_T_42_rs3; // @[package.scala 32:76]
  assign _io_out_T_45 = _io_out_T == 5'h17; // @[package.scala 32:86]
  assign io_out_s_23_bits = {{3'd0}, _io_out_s_T_177}; // @[RVC.scala 21:19 RVC.scala 22:14]
  assign _io_out_T_46_bits = _io_out_T_45 ? io_out_s_23_bits : _io_out_T_44_bits; // @[package.scala 32:76]
  assign _io_out_T_46_rd = _io_out_T_45 ? io_out_s_hi_hi_lo_8 : _io_out_T_44_rd; // @[package.scala 32:76]
  assign _io_out_T_46_rs1 = _io_out_T_45 ? 5'h2 : _io_out_T_44_rs1; // @[package.scala 32:76]
  assign _io_out_T_46_rs2 = _io_out_T_45 ? io_out_s_lo_52 : _io_out_T_44_rs2; // @[package.scala 32:76]
  assign _io_out_T_46_rs3 = _io_out_T_45 ? io_out_s_0_rs3 : _io_out_T_44_rs3; // @[package.scala 32:76]
  assign _io_out_T_47 = _io_out_T == 5'h18; // @[package.scala 32:86]
  assign _io_out_T_48_bits = _io_out_T_47 ? io_in : _io_out_T_46_bits; // @[package.scala 32:76]
  assign _io_out_T_48_rd = _io_out_T_47 ? io_out_s_hi_hi_lo_8 : _io_out_T_46_rd; // @[package.scala 32:76]
  assign _io_out_T_48_rs1 = _io_out_T_47 ? io_out_s_24_rs1 : _io_out_T_46_rs1; // @[package.scala 32:76]
  assign _io_out_T_48_rs2 = _io_out_T_47 ? io_out_s_24_rs2 : _io_out_T_46_rs2; // @[package.scala 32:76]
  assign _io_out_T_48_rs3 = _io_out_T_47 ? io_out_s_0_rs3 : _io_out_T_46_rs3; // @[package.scala 32:76]
  assign _io_out_T_49 = _io_out_T == 5'h19; // @[package.scala 32:86]
  assign _io_out_T_50_bits = _io_out_T_49 ? io_in : _io_out_T_48_bits; // @[package.scala 32:76]
  assign _io_out_T_50_rd = _io_out_T_49 ? io_out_s_hi_hi_lo_8 : _io_out_T_48_rd; // @[package.scala 32:76]
  assign _io_out_T_50_rs1 = _io_out_T_49 ? io_out_s_24_rs1 : _io_out_T_48_rs1; // @[package.scala 32:76]
  assign _io_out_T_50_rs2 = _io_out_T_49 ? io_out_s_24_rs2 : _io_out_T_48_rs2; // @[package.scala 32:76]
  assign _io_out_T_50_rs3 = _io_out_T_49 ? io_out_s_0_rs3 : _io_out_T_48_rs3; // @[package.scala 32:76]
  assign _io_out_T_51 = _io_out_T == 5'h1a; // @[package.scala 32:86]
  assign _io_out_T_52_bits = _io_out_T_51 ? io_in : _io_out_T_50_bits; // @[package.scala 32:76]
  assign _io_out_T_52_rd = _io_out_T_51 ? io_out_s_hi_hi_lo_8 : _io_out_T_50_rd; // @[package.scala 32:76]
  assign _io_out_T_52_rs1 = _io_out_T_51 ? io_out_s_24_rs1 : _io_out_T_50_rs1; // @[package.scala 32:76]
  assign _io_out_T_52_rs2 = _io_out_T_51 ? io_out_s_24_rs2 : _io_out_T_50_rs2; // @[package.scala 32:76]
  assign _io_out_T_52_rs3 = _io_out_T_51 ? io_out_s_0_rs3 : _io_out_T_50_rs3; // @[package.scala 32:76]
  assign _io_out_T_53 = _io_out_T == 5'h1b; // @[package.scala 32:86]
  assign _io_out_T_54_bits = _io_out_T_53 ? io_in : _io_out_T_52_bits; // @[package.scala 32:76]
  assign _io_out_T_54_rd = _io_out_T_53 ? io_out_s_hi_hi_lo_8 : _io_out_T_52_rd; // @[package.scala 32:76]
  assign _io_out_T_54_rs1 = _io_out_T_53 ? io_out_s_24_rs1 : _io_out_T_52_rs1; // @[package.scala 32:76]
  assign _io_out_T_54_rs2 = _io_out_T_53 ? io_out_s_24_rs2 : _io_out_T_52_rs2; // @[package.scala 32:76]
  assign _io_out_T_54_rs3 = _io_out_T_53 ? io_out_s_0_rs3 : _io_out_T_52_rs3; // @[package.scala 32:76]
  assign _io_out_T_55 = _io_out_T == 5'h1c; // @[package.scala 32:86]
  assign _io_out_T_56_bits = _io_out_T_55 ? io_in : _io_out_T_54_bits; // @[package.scala 32:76]
  assign _io_out_T_56_rd = _io_out_T_55 ? io_out_s_hi_hi_lo_8 : _io_out_T_54_rd; // @[package.scala 32:76]
  assign _io_out_T_56_rs1 = _io_out_T_55 ? io_out_s_24_rs1 : _io_out_T_54_rs1; // @[package.scala 32:76]
  assign _io_out_T_56_rs2 = _io_out_T_55 ? io_out_s_24_rs2 : _io_out_T_54_rs2; // @[package.scala 32:76]
  assign _io_out_T_56_rs3 = _io_out_T_55 ? io_out_s_0_rs3 : _io_out_T_54_rs3; // @[package.scala 32:76]
  assign _io_out_T_57 = _io_out_T == 5'h1d; // @[package.scala 32:86]
  assign _io_out_T_58_bits = _io_out_T_57 ? io_in : _io_out_T_56_bits; // @[package.scala 32:76]
  assign _io_out_T_58_rd = _io_out_T_57 ? io_out_s_hi_hi_lo_8 : _io_out_T_56_rd; // @[package.scala 32:76]
  assign _io_out_T_58_rs1 = _io_out_T_57 ? io_out_s_24_rs1 : _io_out_T_56_rs1; // @[package.scala 32:76]
  assign _io_out_T_58_rs2 = _io_out_T_57 ? io_out_s_24_rs2 : _io_out_T_56_rs2; // @[package.scala 32:76]
  assign _io_out_T_58_rs3 = _io_out_T_57 ? io_out_s_0_rs3 : _io_out_T_56_rs3; // @[package.scala 32:76]
  assign _io_out_T_59 = _io_out_T == 5'h1e; // @[package.scala 32:86]
  assign _io_out_T_60_bits = _io_out_T_59 ? io_in : _io_out_T_58_bits; // @[package.scala 32:76]
  assign _io_out_T_60_rd = _io_out_T_59 ? io_out_s_hi_hi_lo_8 : _io_out_T_58_rd; // @[package.scala 32:76]
  assign _io_out_T_60_rs1 = _io_out_T_59 ? io_out_s_24_rs1 : _io_out_T_58_rs1; // @[package.scala 32:76]
  assign _io_out_T_60_rs2 = _io_out_T_59 ? io_out_s_24_rs2 : _io_out_T_58_rs2; // @[package.scala 32:76]
  assign _io_out_T_60_rs3 = _io_out_T_59 ? io_out_s_0_rs3 : _io_out_T_58_rs3; // @[package.scala 32:76]
  assign _io_out_T_61 = _io_out_T == 5'h1f; // @[package.scala 32:86]
  assign io_out_bits = _io_out_T_61 ? io_in : _io_out_T_60_bits; // @[RVC.scala 164:12]
  assign io_out_rd = _io_out_T_61 ? io_out_s_hi_hi_lo_8 : _io_out_T_60_rd; // @[RVC.scala 164:12]
  assign io_out_rs1 = _io_out_T_61 ? io_out_s_24_rs1 : _io_out_T_60_rs1; // @[RVC.scala 164:12]
  assign io_out_rs2 = _io_out_T_61 ? io_out_s_24_rs2 : _io_out_T_60_rs2; // @[RVC.scala 164:12]
  assign io_out_rs3 = _io_out_T_61 ? io_out_s_0_rs3 : _io_out_T_60_rs3; // @[RVC.scala 164:12]
  assign io_rvc = io_in[1:0] != 2'h3; // @[RVC.scala 163:12]
  assign RVCExpander_covSum = 30'h0;
  assign io_covSum = RVCExpander_covSum;
  assign metaAssert = 1'h0;
endmodule
module MulAddRecFNToRaw_preMul(
  input  [1:0]  io_op,
  input  [32:0] io_a,
  input  [32:0] io_b,
  input  [32:0] io_c,
  output [23:0] io_mulAddA,
  output [23:0] io_mulAddB,
  output [47:0] io_mulAddC,
  output        io_toPostMul_isSigNaNAny,
  output        io_toPostMul_isNaNAOrB,
  output        io_toPostMul_isInfA,
  output        io_toPostMul_isZeroA,
  output        io_toPostMul_isInfB,
  output        io_toPostMul_isZeroB,
  output        io_toPostMul_signProd,
  output        io_toPostMul_isNaNC,
  output        io_toPostMul_isInfC,
  output        io_toPostMul_isZeroC,
  output [9:0]  io_toPostMul_sExpSum,
  output        io_toPostMul_doSubMags,
  output        io_toPostMul_CIsDominant,
  output [4:0]  io_toPostMul_CDom_CAlignDist,
  output [25:0] io_toPostMul_highAlignedSigC,
  output        io_toPostMul_bit0AlignedSigC,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire [8:0] rawA_exp; // @[rawFloatFromRecFN.scala 50:21]
  wire  rawA_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  rawA_isSpecial; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawA__isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawA__sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [9:0] rawA__sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire  rawA_out_sig_hi_lo; // @[rawFloatFromRecFN.scala 60:39]
  wire [22:0] rawA_out_sig_lo; // @[rawFloatFromRecFN.scala 60:51]
  wire [24:0] rawA__sig; // @[Cat.scala 30:58]
  wire [8:0] rawB_exp; // @[rawFloatFromRecFN.scala 50:21]
  wire  rawB_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  rawB_isSpecial; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawB__isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawB__sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [9:0] rawB__sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire  rawB_out_sig_hi_lo; // @[rawFloatFromRecFN.scala 60:39]
  wire [22:0] rawB_out_sig_lo; // @[rawFloatFromRecFN.scala 60:51]
  wire [24:0] rawB__sig; // @[Cat.scala 30:58]
  wire [8:0] rawC_exp; // @[rawFloatFromRecFN.scala 50:21]
  wire  rawC_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  rawC_isSpecial; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawC__isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawC__sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [9:0] rawC__sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire  rawC_out_sig_hi_lo; // @[rawFloatFromRecFN.scala 60:39]
  wire [22:0] rawC_out_sig_lo; // @[rawFloatFromRecFN.scala 60:51]
  wire [24:0] rawC__sig; // @[Cat.scala 30:58]
  wire  _signProd_T; // @[MulAddRecFN.scala 98:30]
  wire  signProd; // @[MulAddRecFN.scala 98:42]
  wire [10:0] _sExpAlignedProd_T; // @[MulAddRecFN.scala 101:19]
  wire [10:0] sExpAlignedProd; // @[MulAddRecFN.scala 101:32]
  wire  _doSubMags_T; // @[MulAddRecFN.scala 103:30]
  wire  doSubMags; // @[MulAddRecFN.scala 103:42]
  wire [10:0] _GEN_0; // @[MulAddRecFN.scala 107:42]
  wire [10:0] sNatCAlignDist; // @[MulAddRecFN.scala 107:42]
  wire [9:0] posNatCAlignDist; // @[MulAddRecFN.scala 108:42]
  wire  _isMinCAlign_T; // @[MulAddRecFN.scala 109:35]
  wire  _isMinCAlign_T_1; // @[MulAddRecFN.scala 109:69]
  wire  isMinCAlign; // @[MulAddRecFN.scala 109:50]
  wire  _CIsDominant_T_1; // @[MulAddRecFN.scala 111:60]
  wire  _CIsDominant_T_2; // @[MulAddRecFN.scala 111:39]
  wire  CIsDominant; // @[MulAddRecFN.scala 111:23]
  wire  _CAlignDist_T; // @[MulAddRecFN.scala 115:34]
  wire [6:0] _CAlignDist_T_2; // @[MulAddRecFN.scala 115:16]
  wire [6:0] CAlignDist; // @[MulAddRecFN.scala 113:12]
  wire [24:0] mainAlignedSigC_hi; // @[MulAddRecFN.scala 121:16]
  wire [52:0] mainAlignedSigC_lo; // @[Bitwise.scala 72:12]
  wire [77:0] _mainAlignedSigC_T_3; // @[MulAddRecFN.scala 123:11]
  wire [77:0] mainAlignedSigC; // @[MulAddRecFN.scala 123:17]
  wire [26:0] _reduced4CExtra_T; // @[MulAddRecFN.scala 125:30]
  wire  reduced4CExtra_reducedVec_0; // @[primitives.scala 121:54]
  wire  reduced4CExtra_reducedVec_1; // @[primitives.scala 121:54]
  wire  reduced4CExtra_reducedVec_2; // @[primitives.scala 121:54]
  wire  reduced4CExtra_reducedVec_3; // @[primitives.scala 121:54]
  wire  reduced4CExtra_reducedVec_4; // @[primitives.scala 121:54]
  wire  reduced4CExtra_reducedVec_5; // @[primitives.scala 121:54]
  wire  reduced4CExtra_reducedVec_6; // @[primitives.scala 124:57]
  wire [6:0] _reduced4CExtra_T_1; // @[primitives.scala 125:20]
  wire [32:0] reduced4CExtra_shift; // @[primitives.scala 77:58]
  wire  reduced4CExtra_hi_1; // @[Bitwise.scala 109:18]
  wire  reduced4CExtra_lo_1; // @[Bitwise.scala 109:44]
  wire  reduced4CExtra_hi_3; // @[Bitwise.scala 109:18]
  wire  reduced4CExtra_lo_2; // @[Bitwise.scala 109:44]
  wire  reduced4CExtra_hi_5; // @[Bitwise.scala 109:18]
  wire  reduced4CExtra_lo_4; // @[Bitwise.scala 109:44]
  wire [5:0] _reduced4CExtra_T_8; // @[Cat.scala 30:58]
  wire [6:0] _GEN_1; // @[MulAddRecFN.scala 125:68]
  wire [6:0] _reduced4CExtra_T_9; // @[MulAddRecFN.scala 125:68]
  wire  reduced4CExtra; // @[MulAddRecFN.scala 133:11]
  wire  _alignedSigC_T_2; // @[MulAddRecFN.scala 137:39]
  wire  _alignedSigC_T_4; // @[MulAddRecFN.scala 137:44]
  wire  _alignedSigC_T_6; // @[MulAddRecFN.scala 138:39]
  wire  _alignedSigC_T_7; // @[MulAddRecFN.scala 138:44]
  wire  alignedSigC_lo; // @[MulAddRecFN.scala 136:16]
  wire [74:0] alignedSigC_hi; // @[Cat.scala 30:58]
  wire [75:0] alignedSigC; // @[Cat.scala 30:58]
  wire  _io_toPostMul_isSigNaNAny_T_2; // @[common.scala 81:46]
  wire  _io_toPostMul_isSigNaNAny_T_5; // @[common.scala 81:46]
  wire  _io_toPostMul_isSigNaNAny_T_6; // @[MulAddRecFN.scala 149:32]
  wire  _io_toPostMul_isSigNaNAny_T_9; // @[common.scala 81:46]
  wire [10:0] _io_toPostMul_sExpSum_T_2; // @[MulAddRecFN.scala 161:53]
  wire [10:0] _io_toPostMul_sExpSum_T_3; // @[MulAddRecFN.scala 161:12]
  wire [29:0] MulAddRecFNToRaw_preMul_covSum;
  assign rawA_exp = io_a[31:23]; // @[rawFloatFromRecFN.scala 50:21]
  assign rawA_isZero = rawA_exp[8:6] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign rawA_isSpecial = rawA_exp[8:7] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawA__isNaN = rawA_isSpecial & rawA_exp[6]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawA__sign = io_a[32]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawA__sExp = {1'b0,$signed(rawA_exp)}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawA_out_sig_hi_lo = ~rawA_isZero; // @[rawFloatFromRecFN.scala 60:39]
  assign rawA_out_sig_lo = io_a[22:0]; // @[rawFloatFromRecFN.scala 60:51]
  assign rawA__sig = {1'h0,rawA_out_sig_hi_lo,rawA_out_sig_lo}; // @[Cat.scala 30:58]
  assign rawB_exp = io_b[31:23]; // @[rawFloatFromRecFN.scala 50:21]
  assign rawB_isZero = rawB_exp[8:6] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign rawB_isSpecial = rawB_exp[8:7] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawB__isNaN = rawB_isSpecial & rawB_exp[6]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawB__sign = io_b[32]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawB__sExp = {1'b0,$signed(rawB_exp)}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawB_out_sig_hi_lo = ~rawB_isZero; // @[rawFloatFromRecFN.scala 60:39]
  assign rawB_out_sig_lo = io_b[22:0]; // @[rawFloatFromRecFN.scala 60:51]
  assign rawB__sig = {1'h0,rawB_out_sig_hi_lo,rawB_out_sig_lo}; // @[Cat.scala 30:58]
  assign rawC_exp = io_c[31:23]; // @[rawFloatFromRecFN.scala 50:21]
  assign rawC_isZero = rawC_exp[8:6] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign rawC_isSpecial = rawC_exp[8:7] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawC__isNaN = rawC_isSpecial & rawC_exp[6]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawC__sign = io_c[32]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawC__sExp = {1'b0,$signed(rawC_exp)}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawC_out_sig_hi_lo = ~rawC_isZero; // @[rawFloatFromRecFN.scala 60:39]
  assign rawC_out_sig_lo = io_c[22:0]; // @[rawFloatFromRecFN.scala 60:51]
  assign rawC__sig = {1'h0,rawC_out_sig_hi_lo,rawC_out_sig_lo}; // @[Cat.scala 30:58]
  assign _signProd_T = rawA__sign ^ rawB__sign; // @[MulAddRecFN.scala 98:30]
  assign signProd = _signProd_T ^ io_op[1]; // @[MulAddRecFN.scala 98:42]
  assign _sExpAlignedProd_T = $signed(rawA__sExp) + $signed(rawB__sExp); // @[MulAddRecFN.scala 101:19]
  assign sExpAlignedProd = $signed(_sExpAlignedProd_T) + -11'she5; // @[MulAddRecFN.scala 101:32]
  assign _doSubMags_T = signProd ^ rawC__sign; // @[MulAddRecFN.scala 103:30]
  assign doSubMags = _doSubMags_T ^ io_op[0]; // @[MulAddRecFN.scala 103:42]
  assign _GEN_0 = {{1{rawC__sExp[9]}},rawC__sExp}; // @[MulAddRecFN.scala 107:42]
  assign sNatCAlignDist = $signed(sExpAlignedProd) - $signed(_GEN_0); // @[MulAddRecFN.scala 107:42]
  assign posNatCAlignDist = sNatCAlignDist[9:0]; // @[MulAddRecFN.scala 108:42]
  assign _isMinCAlign_T = rawA_isZero | rawB_isZero; // @[MulAddRecFN.scala 109:35]
  assign _isMinCAlign_T_1 = $signed(sNatCAlignDist) < 11'sh0; // @[MulAddRecFN.scala 109:69]
  assign isMinCAlign = _isMinCAlign_T | _isMinCAlign_T_1; // @[MulAddRecFN.scala 109:50]
  assign _CIsDominant_T_1 = posNatCAlignDist <= 10'h18; // @[MulAddRecFN.scala 111:60]
  assign _CIsDominant_T_2 = isMinCAlign | _CIsDominant_T_1; // @[MulAddRecFN.scala 111:39]
  assign CIsDominant = rawC_out_sig_hi_lo & _CIsDominant_T_2; // @[MulAddRecFN.scala 111:23]
  assign _CAlignDist_T = posNatCAlignDist < 10'h4a; // @[MulAddRecFN.scala 115:34]
  assign _CAlignDist_T_2 = _CAlignDist_T ? posNatCAlignDist[6:0] : 7'h4a; // @[MulAddRecFN.scala 115:16]
  assign CAlignDist = isMinCAlign ? 7'h0 : _CAlignDist_T_2; // @[MulAddRecFN.scala 113:12]
  assign mainAlignedSigC_hi = doSubMags ? ~rawC__sig : rawC__sig; // @[MulAddRecFN.scala 121:16]
  assign mainAlignedSigC_lo = doSubMags ? 53'h1fffffffffffff : 53'h0; // @[Bitwise.scala 72:12]
  assign _mainAlignedSigC_T_3 = {mainAlignedSigC_hi,mainAlignedSigC_lo}; // @[MulAddRecFN.scala 123:11]
  assign mainAlignedSigC = $signed(_mainAlignedSigC_T_3) >>> CAlignDist; // @[MulAddRecFN.scala 123:17]
  assign _reduced4CExtra_T = {rawC__sig, 2'h0}; // @[MulAddRecFN.scala 125:30]
  assign reduced4CExtra_reducedVec_0 = |_reduced4CExtra_T[3:0]; // @[primitives.scala 121:54]
  assign reduced4CExtra_reducedVec_1 = |_reduced4CExtra_T[7:4]; // @[primitives.scala 121:54]
  assign reduced4CExtra_reducedVec_2 = |_reduced4CExtra_T[11:8]; // @[primitives.scala 121:54]
  assign reduced4CExtra_reducedVec_3 = |_reduced4CExtra_T[15:12]; // @[primitives.scala 121:54]
  assign reduced4CExtra_reducedVec_4 = |_reduced4CExtra_T[19:16]; // @[primitives.scala 121:54]
  assign reduced4CExtra_reducedVec_5 = |_reduced4CExtra_T[23:20]; // @[primitives.scala 121:54]
  assign reduced4CExtra_reducedVec_6 = |_reduced4CExtra_T[26:24]; // @[primitives.scala 124:57]
  assign _reduced4CExtra_T_1 = {reduced4CExtra_reducedVec_6,reduced4CExtra_reducedVec_5,reduced4CExtra_reducedVec_4,reduced4CExtra_reducedVec_3,reduced4CExtra_reducedVec_2,reduced4CExtra_reducedVec_1,reduced4CExtra_reducedVec_0}; // @[primitives.scala 125:20]
  assign reduced4CExtra_shift = -33'sh100000000 >>> CAlignDist[6:2]; // @[primitives.scala 77:58]
  assign reduced4CExtra_hi_1 = reduced4CExtra_shift[14]; // @[Bitwise.scala 109:18]
  assign reduced4CExtra_lo_1 = reduced4CExtra_shift[15]; // @[Bitwise.scala 109:44]
  assign reduced4CExtra_hi_3 = reduced4CExtra_shift[16]; // @[Bitwise.scala 109:18]
  assign reduced4CExtra_lo_2 = reduced4CExtra_shift[17]; // @[Bitwise.scala 109:44]
  assign reduced4CExtra_hi_5 = reduced4CExtra_shift[18]; // @[Bitwise.scala 109:18]
  assign reduced4CExtra_lo_4 = reduced4CExtra_shift[19]; // @[Bitwise.scala 109:44]
  assign _reduced4CExtra_T_8 = {reduced4CExtra_hi_1,reduced4CExtra_lo_1,reduced4CExtra_hi_3,reduced4CExtra_lo_2,reduced4CExtra_hi_5,reduced4CExtra_lo_4}; // @[Cat.scala 30:58]
  assign _GEN_1 = {{1'd0}, _reduced4CExtra_T_8}; // @[MulAddRecFN.scala 125:68]
  assign _reduced4CExtra_T_9 = _reduced4CExtra_T_1 & _GEN_1; // @[MulAddRecFN.scala 125:68]
  assign reduced4CExtra = |_reduced4CExtra_T_9; // @[MulAddRecFN.scala 133:11]
  assign _alignedSigC_T_2 = &mainAlignedSigC[2:0]; // @[MulAddRecFN.scala 137:39]
  assign _alignedSigC_T_4 = _alignedSigC_T_2 & ~reduced4CExtra; // @[MulAddRecFN.scala 137:44]
  assign _alignedSigC_T_6 = |mainAlignedSigC[2:0]; // @[MulAddRecFN.scala 138:39]
  assign _alignedSigC_T_7 = _alignedSigC_T_6 | reduced4CExtra; // @[MulAddRecFN.scala 138:44]
  assign alignedSigC_lo = doSubMags ? _alignedSigC_T_4 : _alignedSigC_T_7; // @[MulAddRecFN.scala 136:16]
  assign alignedSigC_hi = mainAlignedSigC[77:3]; // @[Cat.scala 30:58]
  assign alignedSigC = {alignedSigC_hi,alignedSigC_lo}; // @[Cat.scala 30:58]
  assign _io_toPostMul_isSigNaNAny_T_2 = rawA__isNaN & ~rawA__sig[22]; // @[common.scala 81:46]
  assign _io_toPostMul_isSigNaNAny_T_5 = rawB__isNaN & ~rawB__sig[22]; // @[common.scala 81:46]
  assign _io_toPostMul_isSigNaNAny_T_6 = _io_toPostMul_isSigNaNAny_T_2 | _io_toPostMul_isSigNaNAny_T_5; // @[MulAddRecFN.scala 149:32]
  assign _io_toPostMul_isSigNaNAny_T_9 = rawC__isNaN & ~rawC__sig[22]; // @[common.scala 81:46]
  assign _io_toPostMul_sExpSum_T_2 = $signed(sExpAlignedProd) - 11'sh18; // @[MulAddRecFN.scala 161:53]
  assign _io_toPostMul_sExpSum_T_3 = CIsDominant ? $signed({{1{rawC__sExp[9]}},rawC__sExp}) : $signed(_io_toPostMul_sExpSum_T_2); // @[MulAddRecFN.scala 161:12]
  assign io_mulAddA = rawA__sig[23:0]; // @[MulAddRecFN.scala 144:16]
  assign io_mulAddB = rawB__sig[23:0]; // @[MulAddRecFN.scala 145:16]
  assign io_mulAddC = alignedSigC[48:1]; // @[MulAddRecFN.scala 146:16]
  assign io_toPostMul_isSigNaNAny = _io_toPostMul_isSigNaNAny_T_6 | _io_toPostMul_isSigNaNAny_T_9; // @[MulAddRecFN.scala 148:30]
  assign io_toPostMul_isNaNAOrB = rawA__isNaN | rawB__isNaN; // @[MulAddRecFN.scala 151:28]
  assign io_toPostMul_isInfA = rawA_isSpecial & ~rawA_exp[6]; // @[MulAddRecFN.scala 152:28]
  assign io_toPostMul_isZeroA = rawA_exp[8:6] == 3'h0; // @[MulAddRecFN.scala 153:28]
  assign io_toPostMul_isInfB = rawB_isSpecial & ~rawB_exp[6]; // @[MulAddRecFN.scala 154:28]
  assign io_toPostMul_isZeroB = rawB_exp[8:6] == 3'h0; // @[MulAddRecFN.scala 155:28]
  assign io_toPostMul_signProd = _signProd_T ^ io_op[1]; // @[MulAddRecFN.scala 156:28]
  assign io_toPostMul_isNaNC = rawC_isSpecial & rawC_exp[6]; // @[MulAddRecFN.scala 157:28]
  assign io_toPostMul_isInfC = rawC_isSpecial & ~rawC_exp[6]; // @[MulAddRecFN.scala 158:28]
  assign io_toPostMul_isZeroC = rawC_exp[8:6] == 3'h0; // @[MulAddRecFN.scala 159:28]
  assign io_toPostMul_sExpSum = _io_toPostMul_sExpSum_T_3[9:0]; // @[MulAddRecFN.scala 160:28]
  assign io_toPostMul_doSubMags = _doSubMags_T ^ io_op[0]; // @[MulAddRecFN.scala 162:28]
  assign io_toPostMul_CIsDominant = rawC_out_sig_hi_lo & _CIsDominant_T_2; // @[MulAddRecFN.scala 163:30]
  assign io_toPostMul_CDom_CAlignDist = CAlignDist[4:0]; // @[MulAddRecFN.scala 164:34]
  assign io_toPostMul_highAlignedSigC = alignedSigC[74:49]; // @[MulAddRecFN.scala 165:34]
  assign io_toPostMul_bit0AlignedSigC = alignedSigC[0]; // @[MulAddRecFN.scala 167:34]
  assign MulAddRecFNToRaw_preMul_covSum = 30'h0;
  assign io_covSum = MulAddRecFNToRaw_preMul_covSum;
  assign metaAssert = 1'h0;
endmodule
module MulAddRecFNToRaw_postMul(
  input         io_fromPreMul_isSigNaNAny,
  input         io_fromPreMul_isNaNAOrB,
  input         io_fromPreMul_isInfA,
  input         io_fromPreMul_isZeroA,
  input         io_fromPreMul_isInfB,
  input         io_fromPreMul_isZeroB,
  input         io_fromPreMul_signProd,
  input         io_fromPreMul_isNaNC,
  input         io_fromPreMul_isInfC,
  input         io_fromPreMul_isZeroC,
  input  [9:0]  io_fromPreMul_sExpSum,
  input         io_fromPreMul_doSubMags,
  input         io_fromPreMul_CIsDominant,
  input  [4:0]  io_fromPreMul_CDom_CAlignDist,
  input  [25:0] io_fromPreMul_highAlignedSigC,
  input         io_fromPreMul_bit0AlignedSigC,
  input  [48:0] io_mulAddResult,
  input  [2:0]  io_roundingMode,
  output        io_invalidExc,
  output        io_rawOut_isNaN,
  output        io_rawOut_isInf,
  output        io_rawOut_isZero,
  output        io_rawOut_sign,
  output [9:0]  io_rawOut_sExp,
  output [26:0] io_rawOut_sig,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  roundingMode_min; // @[MulAddRecFN.scala 188:45]
  wire  CDom_sign; // @[MulAddRecFN.scala 192:42]
  wire [25:0] _sigSum_T_2; // @[MulAddRecFN.scala 195:47]
  wire [25:0] sigSum_hi_hi; // @[MulAddRecFN.scala 194:16]
  wire [47:0] sigSum_hi_lo; // @[MulAddRecFN.scala 198:28]
  wire [74:0] sigSum; // @[Cat.scala 30:58]
  wire [1:0] _CDom_sExp_T; // @[MulAddRecFN.scala 205:69]
  wire [9:0] _GEN_0; // @[MulAddRecFN.scala 205:43]
  wire [9:0] CDom_sExp; // @[MulAddRecFN.scala 205:43]
  wire [1:0] CDom_absSigSum_hi_lo; // @[MulAddRecFN.scala 211:46]
  wire [46:0] CDom_absSigSum_lo; // @[MulAddRecFN.scala 212:23]
  wire [49:0] _CDom_absSigSum_T_2; // @[Cat.scala 30:58]
  wire [49:0] CDom_absSigSum; // @[MulAddRecFN.scala 207:12]
  wire  _CDom_absSigSumExtra_T_2; // @[MulAddRecFN.scala 217:36]
  wire  _CDom_absSigSumExtra_T_4; // @[MulAddRecFN.scala 218:37]
  wire  CDom_absSigSumExtra; // @[MulAddRecFN.scala 216:12]
  wire [80:0] _GEN_1; // @[MulAddRecFN.scala 221:24]
  wire [80:0] _CDom_mainSig_T; // @[MulAddRecFN.scala 221:24]
  wire [28:0] CDom_mainSig; // @[MulAddRecFN.scala 221:56]
  wire [26:0] _CDom_reduced4SigExtra_T_1; // @[MulAddRecFN.scala 224:53]
  wire  CDom_reduced4SigExtra_reducedVec_0; // @[primitives.scala 121:54]
  wire  CDom_reduced4SigExtra_reducedVec_1; // @[primitives.scala 121:54]
  wire  CDom_reduced4SigExtra_reducedVec_2; // @[primitives.scala 121:54]
  wire  CDom_reduced4SigExtra_reducedVec_3; // @[primitives.scala 121:54]
  wire  CDom_reduced4SigExtra_reducedVec_4; // @[primitives.scala 121:54]
  wire  CDom_reduced4SigExtra_reducedVec_5; // @[primitives.scala 121:54]
  wire  CDom_reduced4SigExtra_reducedVec_6; // @[primitives.scala 124:57]
  wire [6:0] _CDom_reduced4SigExtra_T_2; // @[primitives.scala 125:20]
  wire [8:0] CDom_reduced4SigExtra_shift; // @[primitives.scala 77:58]
  wire  CDom_reduced4SigExtra_hi_1; // @[Bitwise.scala 109:18]
  wire  CDom_reduced4SigExtra_lo_1; // @[Bitwise.scala 109:44]
  wire  CDom_reduced4SigExtra_hi_3; // @[Bitwise.scala 109:18]
  wire  CDom_reduced4SigExtra_lo_2; // @[Bitwise.scala 109:44]
  wire  CDom_reduced4SigExtra_hi_5; // @[Bitwise.scala 109:18]
  wire  CDom_reduced4SigExtra_lo_4; // @[Bitwise.scala 109:44]
  wire [5:0] _CDom_reduced4SigExtra_T_10; // @[Cat.scala 30:58]
  wire [6:0] _GEN_2; // @[MulAddRecFN.scala 224:72]
  wire [6:0] _CDom_reduced4SigExtra_T_11; // @[MulAddRecFN.scala 224:72]
  wire  CDom_reduced4SigExtra; // @[MulAddRecFN.scala 225:73]
  wire [25:0] CDom_sig_hi; // @[MulAddRecFN.scala 227:25]
  wire  _CDom_sig_T_1; // @[MulAddRecFN.scala 228:32]
  wire  _CDom_sig_T_2; // @[MulAddRecFN.scala 228:36]
  wire  CDom_sig_lo; // @[MulAddRecFN.scala 228:61]
  wire [26:0] CDom_sig; // @[Cat.scala 30:58]
  wire  notCDom_signSigSum; // @[MulAddRecFN.scala 234:36]
  wire [50:0] _GEN_3; // @[MulAddRecFN.scala 238:41]
  wire [50:0] _notCDom_absSigSum_T_4; // @[MulAddRecFN.scala 238:41]
  wire [50:0] notCDom_absSigSum; // @[MulAddRecFN.scala 236:12]
  wire  notCDom_reduced2AbsSigSum_reducedVec_0; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_1; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_2; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_3; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_4; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_5; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_6; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_7; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_8; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_9; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_10; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_11; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_12; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_13; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_14; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_15; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_16; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_17; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_18; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_19; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_20; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_21; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_22; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_23; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_24; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_25; // @[primitives.scala 107:57]
  wire [5:0] notCDom_reduced2AbsSigSum_lo_lo; // @[primitives.scala 108:20]
  wire [12:0] notCDom_reduced2AbsSigSum_lo; // @[primitives.scala 108:20]
  wire [5:0] notCDom_reduced2AbsSigSum_hi_lo; // @[primitives.scala 108:20]
  wire [25:0] notCDom_reduced2AbsSigSum; // @[primitives.scala 108:20]
  wire [4:0] _notCDom_normDistReduced2_T_26; // @[Mux.scala 47:69]
  wire [4:0] _notCDom_normDistReduced2_T_27; // @[Mux.scala 47:69]
  wire [4:0] _notCDom_normDistReduced2_T_28; // @[Mux.scala 47:69]
  wire [4:0] _notCDom_normDistReduced2_T_29; // @[Mux.scala 47:69]
  wire [4:0] _notCDom_normDistReduced2_T_30; // @[Mux.scala 47:69]
  wire [4:0] _notCDom_normDistReduced2_T_31; // @[Mux.scala 47:69]
  wire [4:0] _notCDom_normDistReduced2_T_32; // @[Mux.scala 47:69]
  wire [4:0] _notCDom_normDistReduced2_T_33; // @[Mux.scala 47:69]
  wire [4:0] _notCDom_normDistReduced2_T_34; // @[Mux.scala 47:69]
  wire [4:0] _notCDom_normDistReduced2_T_35; // @[Mux.scala 47:69]
  wire [4:0] _notCDom_normDistReduced2_T_36; // @[Mux.scala 47:69]
  wire [4:0] _notCDom_normDistReduced2_T_37; // @[Mux.scala 47:69]
  wire [4:0] _notCDom_normDistReduced2_T_38; // @[Mux.scala 47:69]
  wire [4:0] _notCDom_normDistReduced2_T_39; // @[Mux.scala 47:69]
  wire [4:0] _notCDom_normDistReduced2_T_40; // @[Mux.scala 47:69]
  wire [4:0] _notCDom_normDistReduced2_T_41; // @[Mux.scala 47:69]
  wire [4:0] _notCDom_normDistReduced2_T_42; // @[Mux.scala 47:69]
  wire [4:0] _notCDom_normDistReduced2_T_43; // @[Mux.scala 47:69]
  wire [4:0] _notCDom_normDistReduced2_T_44; // @[Mux.scala 47:69]
  wire [4:0] _notCDom_normDistReduced2_T_45; // @[Mux.scala 47:69]
  wire [4:0] _notCDom_normDistReduced2_T_46; // @[Mux.scala 47:69]
  wire [4:0] _notCDom_normDistReduced2_T_47; // @[Mux.scala 47:69]
  wire [4:0] _notCDom_normDistReduced2_T_48; // @[Mux.scala 47:69]
  wire [4:0] _notCDom_normDistReduced2_T_49; // @[Mux.scala 47:69]
  wire [4:0] notCDom_normDistReduced2; // @[Mux.scala 47:69]
  wire [5:0] notCDom_nearNormDist; // @[MulAddRecFN.scala 242:56]
  wire [6:0] _notCDom_sExp_T; // @[MulAddRecFN.scala 243:69]
  wire [9:0] _GEN_4; // @[MulAddRecFN.scala 243:46]
  wire [9:0] notCDom_sExp; // @[MulAddRecFN.scala 243:46]
  wire [113:0] _GEN_5; // @[MulAddRecFN.scala 245:27]
  wire [113:0] _notCDom_mainSig_T; // @[MulAddRecFN.scala 245:27]
  wire [28:0] notCDom_mainSig; // @[MulAddRecFN.scala 245:50]
  wire  notCDom_reduced4SigExtra_reducedVec_0; // @[primitives.scala 104:54]
  wire  notCDom_reduced4SigExtra_reducedVec_1; // @[primitives.scala 104:54]
  wire  notCDom_reduced4SigExtra_reducedVec_2; // @[primitives.scala 104:54]
  wire  notCDom_reduced4SigExtra_reducedVec_3; // @[primitives.scala 104:54]
  wire  notCDom_reduced4SigExtra_reducedVec_4; // @[primitives.scala 104:54]
  wire  notCDom_reduced4SigExtra_reducedVec_5; // @[primitives.scala 104:54]
  wire  notCDom_reduced4SigExtra_reducedVec_6; // @[primitives.scala 107:57]
  wire [6:0] _notCDom_reduced4SigExtra_T_2; // @[primitives.scala 108:20]
  wire [16:0] notCDom_reduced4SigExtra_shift; // @[primitives.scala 77:58]
  wire  notCDom_reduced4SigExtra_hi_1; // @[Bitwise.scala 109:18]
  wire  notCDom_reduced4SigExtra_lo_1; // @[Bitwise.scala 109:44]
  wire  notCDom_reduced4SigExtra_hi_3; // @[Bitwise.scala 109:18]
  wire  notCDom_reduced4SigExtra_lo_2; // @[Bitwise.scala 109:44]
  wire  notCDom_reduced4SigExtra_hi_5; // @[Bitwise.scala 109:18]
  wire  notCDom_reduced4SigExtra_lo_4; // @[Bitwise.scala 109:44]
  wire [5:0] _notCDom_reduced4SigExtra_T_10; // @[Cat.scala 30:58]
  wire [6:0] _GEN_6; // @[MulAddRecFN.scala 249:78]
  wire [6:0] _notCDom_reduced4SigExtra_T_11; // @[MulAddRecFN.scala 249:78]
  wire  notCDom_reduced4SigExtra; // @[MulAddRecFN.scala 251:11]
  wire [25:0] notCDom_sig_hi; // @[MulAddRecFN.scala 253:28]
  wire  _notCDom_sig_T_1; // @[MulAddRecFN.scala 254:35]
  wire  notCDom_sig_lo; // @[MulAddRecFN.scala 254:39]
  wire [26:0] notCDom_sig; // @[Cat.scala 30:58]
  wire  notCDom_completeCancellation; // @[MulAddRecFN.scala 257:50]
  wire  _notCDom_sign_T; // @[MulAddRecFN.scala 261:36]
  wire  notCDom_sign; // @[MulAddRecFN.scala 259:12]
  wire  notNaN_isInfProd; // @[MulAddRecFN.scala 266:49]
  wire  notNaN_isInfOut; // @[MulAddRecFN.scala 267:44]
  wire  _notNaN_addZeros_T; // @[MulAddRecFN.scala 269:32]
  wire  notNaN_addZeros; // @[MulAddRecFN.scala 269:58]
  wire  _io_invalidExc_T; // @[MulAddRecFN.scala 274:31]
  wire  _io_invalidExc_T_1; // @[MulAddRecFN.scala 273:35]
  wire  _io_invalidExc_T_2; // @[MulAddRecFN.scala 275:32]
  wire  _io_invalidExc_T_3; // @[MulAddRecFN.scala 274:57]
  wire  _io_invalidExc_T_6; // @[MulAddRecFN.scala 276:36]
  wire  _io_invalidExc_T_7; // @[MulAddRecFN.scala 277:61]
  wire  _io_invalidExc_T_8; // @[MulAddRecFN.scala 278:35]
  wire  _io_rawOut_isZero_T_1; // @[MulAddRecFN.scala 285:42]
  wire  _io_rawOut_sign_T; // @[MulAddRecFN.scala 287:27]
  wire  _io_rawOut_sign_T_1; // @[MulAddRecFN.scala 288:31]
  wire  _io_rawOut_sign_T_2; // @[MulAddRecFN.scala 287:54]
  wire  _io_rawOut_sign_T_4; // @[MulAddRecFN.scala 289:26]
  wire  _io_rawOut_sign_T_5; // @[MulAddRecFN.scala 289:48]
  wire  _io_rawOut_sign_T_6; // @[MulAddRecFN.scala 290:36]
  wire  _io_rawOut_sign_T_7; // @[MulAddRecFN.scala 288:43]
  wire  _io_rawOut_sign_T_8; // @[MulAddRecFN.scala 291:26]
  wire  _io_rawOut_sign_T_9; // @[MulAddRecFN.scala 292:37]
  wire  _io_rawOut_sign_T_10; // @[MulAddRecFN.scala 291:46]
  wire  _io_rawOut_sign_T_11; // @[MulAddRecFN.scala 290:48]
  wire  _io_rawOut_sign_T_14; // @[MulAddRecFN.scala 293:28]
  wire  _io_rawOut_sign_T_15; // @[MulAddRecFN.scala 294:17]
  wire  _io_rawOut_sign_T_16; // @[MulAddRecFN.scala 293:49]
  wire [29:0] MulAddRecFNToRaw_postMul_covSum;
  assign roundingMode_min = io_roundingMode == 3'h2; // @[MulAddRecFN.scala 188:45]
  assign CDom_sign = io_fromPreMul_signProd ^ io_fromPreMul_doSubMags; // @[MulAddRecFN.scala 192:42]
  assign _sigSum_T_2 = io_fromPreMul_highAlignedSigC + 26'h1; // @[MulAddRecFN.scala 195:47]
  assign sigSum_hi_hi = io_mulAddResult[48] ? _sigSum_T_2 : io_fromPreMul_highAlignedSigC; // @[MulAddRecFN.scala 194:16]
  assign sigSum_hi_lo = io_mulAddResult[47:0]; // @[MulAddRecFN.scala 198:28]
  assign sigSum = {sigSum_hi_hi,sigSum_hi_lo,io_fromPreMul_bit0AlignedSigC}; // @[Cat.scala 30:58]
  assign _CDom_sExp_T = {1'b0,$signed(io_fromPreMul_doSubMags)}; // @[MulAddRecFN.scala 205:69]
  assign _GEN_0 = {{8{_CDom_sExp_T[1]}},_CDom_sExp_T}; // @[MulAddRecFN.scala 205:43]
  assign CDom_sExp = $signed(io_fromPreMul_sExpSum) - $signed(_GEN_0); // @[MulAddRecFN.scala 205:43]
  assign CDom_absSigSum_hi_lo = io_fromPreMul_highAlignedSigC[25:24]; // @[MulAddRecFN.scala 211:46]
  assign CDom_absSigSum_lo = sigSum[72:26]; // @[MulAddRecFN.scala 212:23]
  assign _CDom_absSigSum_T_2 = {1'h0,CDom_absSigSum_hi_lo,CDom_absSigSum_lo}; // @[Cat.scala 30:58]
  assign CDom_absSigSum = io_fromPreMul_doSubMags ? ~sigSum[74:25] : _CDom_absSigSum_T_2; // @[MulAddRecFN.scala 207:12]
  assign _CDom_absSigSumExtra_T_2 = | (~sigSum[24:1]); // @[MulAddRecFN.scala 217:36]
  assign _CDom_absSigSumExtra_T_4 = |sigSum[25:1]; // @[MulAddRecFN.scala 218:37]
  assign CDom_absSigSumExtra = io_fromPreMul_doSubMags ? _CDom_absSigSumExtra_T_2 : _CDom_absSigSumExtra_T_4; // @[MulAddRecFN.scala 216:12]
  assign _GEN_1 = {{31'd0}, CDom_absSigSum}; // @[MulAddRecFN.scala 221:24]
  assign _CDom_mainSig_T = _GEN_1 << io_fromPreMul_CDom_CAlignDist; // @[MulAddRecFN.scala 221:24]
  assign CDom_mainSig = _CDom_mainSig_T[49:21]; // @[MulAddRecFN.scala 221:56]
  assign _CDom_reduced4SigExtra_T_1 = {CDom_absSigSum[23:0], 3'h0}; // @[MulAddRecFN.scala 224:53]
  assign CDom_reduced4SigExtra_reducedVec_0 = |_CDom_reduced4SigExtra_T_1[3:0]; // @[primitives.scala 121:54]
  assign CDom_reduced4SigExtra_reducedVec_1 = |_CDom_reduced4SigExtra_T_1[7:4]; // @[primitives.scala 121:54]
  assign CDom_reduced4SigExtra_reducedVec_2 = |_CDom_reduced4SigExtra_T_1[11:8]; // @[primitives.scala 121:54]
  assign CDom_reduced4SigExtra_reducedVec_3 = |_CDom_reduced4SigExtra_T_1[15:12]; // @[primitives.scala 121:54]
  assign CDom_reduced4SigExtra_reducedVec_4 = |_CDom_reduced4SigExtra_T_1[19:16]; // @[primitives.scala 121:54]
  assign CDom_reduced4SigExtra_reducedVec_5 = |_CDom_reduced4SigExtra_T_1[23:20]; // @[primitives.scala 121:54]
  assign CDom_reduced4SigExtra_reducedVec_6 = |_CDom_reduced4SigExtra_T_1[26:24]; // @[primitives.scala 124:57]
  assign _CDom_reduced4SigExtra_T_2 = {CDom_reduced4SigExtra_reducedVec_6,CDom_reduced4SigExtra_reducedVec_5,CDom_reduced4SigExtra_reducedVec_4,CDom_reduced4SigExtra_reducedVec_3,CDom_reduced4SigExtra_reducedVec_2,CDom_reduced4SigExtra_reducedVec_1,CDom_reduced4SigExtra_reducedVec_0}; // @[primitives.scala 125:20]
  assign CDom_reduced4SigExtra_shift = -9'sh100 >>> ~io_fromPreMul_CDom_CAlignDist[4:2]; // @[primitives.scala 77:58]
  assign CDom_reduced4SigExtra_hi_1 = CDom_reduced4SigExtra_shift[1]; // @[Bitwise.scala 109:18]
  assign CDom_reduced4SigExtra_lo_1 = CDom_reduced4SigExtra_shift[2]; // @[Bitwise.scala 109:44]
  assign CDom_reduced4SigExtra_hi_3 = CDom_reduced4SigExtra_shift[3]; // @[Bitwise.scala 109:18]
  assign CDom_reduced4SigExtra_lo_2 = CDom_reduced4SigExtra_shift[4]; // @[Bitwise.scala 109:44]
  assign CDom_reduced4SigExtra_hi_5 = CDom_reduced4SigExtra_shift[5]; // @[Bitwise.scala 109:18]
  assign CDom_reduced4SigExtra_lo_4 = CDom_reduced4SigExtra_shift[6]; // @[Bitwise.scala 109:44]
  assign _CDom_reduced4SigExtra_T_10 = {CDom_reduced4SigExtra_hi_1,CDom_reduced4SigExtra_lo_1,CDom_reduced4SigExtra_hi_3,CDom_reduced4SigExtra_lo_2,CDom_reduced4SigExtra_hi_5,CDom_reduced4SigExtra_lo_4}; // @[Cat.scala 30:58]
  assign _GEN_2 = {{1'd0}, _CDom_reduced4SigExtra_T_10}; // @[MulAddRecFN.scala 224:72]
  assign _CDom_reduced4SigExtra_T_11 = _CDom_reduced4SigExtra_T_2 & _GEN_2; // @[MulAddRecFN.scala 224:72]
  assign CDom_reduced4SigExtra = |_CDom_reduced4SigExtra_T_11; // @[MulAddRecFN.scala 225:73]
  assign CDom_sig_hi = CDom_mainSig[28:3]; // @[MulAddRecFN.scala 227:25]
  assign _CDom_sig_T_1 = |CDom_mainSig[2:0]; // @[MulAddRecFN.scala 228:32]
  assign _CDom_sig_T_2 = _CDom_sig_T_1 | CDom_reduced4SigExtra; // @[MulAddRecFN.scala 228:36]
  assign CDom_sig_lo = _CDom_sig_T_2 | CDom_absSigSumExtra; // @[MulAddRecFN.scala 228:61]
  assign CDom_sig = {CDom_sig_hi,CDom_sig_lo}; // @[Cat.scala 30:58]
  assign notCDom_signSigSum = sigSum[51]; // @[MulAddRecFN.scala 234:36]
  assign _GEN_3 = {{50'd0}, io_fromPreMul_doSubMags}; // @[MulAddRecFN.scala 238:41]
  assign _notCDom_absSigSum_T_4 = sigSum[50:0] + _GEN_3; // @[MulAddRecFN.scala 238:41]
  assign notCDom_absSigSum = notCDom_signSigSum ? ~sigSum[50:0] : _notCDom_absSigSum_T_4; // @[MulAddRecFN.scala 236:12]
  assign notCDom_reduced2AbsSigSum_reducedVec_0 = |notCDom_absSigSum[1:0]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_1 = |notCDom_absSigSum[3:2]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_2 = |notCDom_absSigSum[5:4]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_3 = |notCDom_absSigSum[7:6]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_4 = |notCDom_absSigSum[9:8]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_5 = |notCDom_absSigSum[11:10]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_6 = |notCDom_absSigSum[13:12]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_7 = |notCDom_absSigSum[15:14]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_8 = |notCDom_absSigSum[17:16]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_9 = |notCDom_absSigSum[19:18]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_10 = |notCDom_absSigSum[21:20]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_11 = |notCDom_absSigSum[23:22]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_12 = |notCDom_absSigSum[25:24]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_13 = |notCDom_absSigSum[27:26]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_14 = |notCDom_absSigSum[29:28]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_15 = |notCDom_absSigSum[31:30]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_16 = |notCDom_absSigSum[33:32]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_17 = |notCDom_absSigSum[35:34]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_18 = |notCDom_absSigSum[37:36]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_19 = |notCDom_absSigSum[39:38]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_20 = |notCDom_absSigSum[41:40]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_21 = |notCDom_absSigSum[43:42]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_22 = |notCDom_absSigSum[45:44]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_23 = |notCDom_absSigSum[47:46]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_24 = |notCDom_absSigSum[49:48]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_25 = |notCDom_absSigSum[50]; // @[primitives.scala 107:57]
  assign notCDom_reduced2AbsSigSum_lo_lo = {notCDom_reduced2AbsSigSum_reducedVec_5,notCDom_reduced2AbsSigSum_reducedVec_4,notCDom_reduced2AbsSigSum_reducedVec_3,notCDom_reduced2AbsSigSum_reducedVec_2,notCDom_reduced2AbsSigSum_reducedVec_1,notCDom_reduced2AbsSigSum_reducedVec_0}; // @[primitives.scala 108:20]
  assign notCDom_reduced2AbsSigSum_lo = {notCDom_reduced2AbsSigSum_reducedVec_12,notCDom_reduced2AbsSigSum_reducedVec_11,notCDom_reduced2AbsSigSum_reducedVec_10,notCDom_reduced2AbsSigSum_reducedVec_9,notCDom_reduced2AbsSigSum_reducedVec_8,notCDom_reduced2AbsSigSum_reducedVec_7,notCDom_reduced2AbsSigSum_reducedVec_6,notCDom_reduced2AbsSigSum_lo_lo}; // @[primitives.scala 108:20]
  assign notCDom_reduced2AbsSigSum_hi_lo = {notCDom_reduced2AbsSigSum_reducedVec_18,notCDom_reduced2AbsSigSum_reducedVec_17,notCDom_reduced2AbsSigSum_reducedVec_16,notCDom_reduced2AbsSigSum_reducedVec_15,notCDom_reduced2AbsSigSum_reducedVec_14,notCDom_reduced2AbsSigSum_reducedVec_13}; // @[primitives.scala 108:20]
  assign notCDom_reduced2AbsSigSum = {notCDom_reduced2AbsSigSum_reducedVec_25,notCDom_reduced2AbsSigSum_reducedVec_24,notCDom_reduced2AbsSigSum_reducedVec_23,notCDom_reduced2AbsSigSum_reducedVec_22,notCDom_reduced2AbsSigSum_reducedVec_21,notCDom_reduced2AbsSigSum_reducedVec_20,notCDom_reduced2AbsSigSum_reducedVec_19,notCDom_reduced2AbsSigSum_hi_lo,notCDom_reduced2AbsSigSum_lo}; // @[primitives.scala 108:20]
  assign _notCDom_normDistReduced2_T_26 = notCDom_reduced2AbsSigSum[1] ? 5'h18 : 5'h19; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_27 = notCDom_reduced2AbsSigSum[2] ? 5'h17 : _notCDom_normDistReduced2_T_26; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_28 = notCDom_reduced2AbsSigSum[3] ? 5'h16 : _notCDom_normDistReduced2_T_27; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_29 = notCDom_reduced2AbsSigSum[4] ? 5'h15 : _notCDom_normDistReduced2_T_28; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_30 = notCDom_reduced2AbsSigSum[5] ? 5'h14 : _notCDom_normDistReduced2_T_29; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_31 = notCDom_reduced2AbsSigSum[6] ? 5'h13 : _notCDom_normDistReduced2_T_30; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_32 = notCDom_reduced2AbsSigSum[7] ? 5'h12 : _notCDom_normDistReduced2_T_31; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_33 = notCDom_reduced2AbsSigSum[8] ? 5'h11 : _notCDom_normDistReduced2_T_32; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_34 = notCDom_reduced2AbsSigSum[9] ? 5'h10 : _notCDom_normDistReduced2_T_33; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_35 = notCDom_reduced2AbsSigSum[10] ? 5'hf : _notCDom_normDistReduced2_T_34; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_36 = notCDom_reduced2AbsSigSum[11] ? 5'he : _notCDom_normDistReduced2_T_35; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_37 = notCDom_reduced2AbsSigSum[12] ? 5'hd : _notCDom_normDistReduced2_T_36; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_38 = notCDom_reduced2AbsSigSum[13] ? 5'hc : _notCDom_normDistReduced2_T_37; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_39 = notCDom_reduced2AbsSigSum[14] ? 5'hb : _notCDom_normDistReduced2_T_38; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_40 = notCDom_reduced2AbsSigSum[15] ? 5'ha : _notCDom_normDistReduced2_T_39; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_41 = notCDom_reduced2AbsSigSum[16] ? 5'h9 : _notCDom_normDistReduced2_T_40; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_42 = notCDom_reduced2AbsSigSum[17] ? 5'h8 : _notCDom_normDistReduced2_T_41; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_43 = notCDom_reduced2AbsSigSum[18] ? 5'h7 : _notCDom_normDistReduced2_T_42; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_44 = notCDom_reduced2AbsSigSum[19] ? 5'h6 : _notCDom_normDistReduced2_T_43; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_45 = notCDom_reduced2AbsSigSum[20] ? 5'h5 : _notCDom_normDistReduced2_T_44; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_46 = notCDom_reduced2AbsSigSum[21] ? 5'h4 : _notCDom_normDistReduced2_T_45; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_47 = notCDom_reduced2AbsSigSum[22] ? 5'h3 : _notCDom_normDistReduced2_T_46; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_48 = notCDom_reduced2AbsSigSum[23] ? 5'h2 : _notCDom_normDistReduced2_T_47; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_49 = notCDom_reduced2AbsSigSum[24] ? 5'h1 : _notCDom_normDistReduced2_T_48; // @[Mux.scala 47:69]
  assign notCDom_normDistReduced2 = notCDom_reduced2AbsSigSum[25] ? 5'h0 : _notCDom_normDistReduced2_T_49; // @[Mux.scala 47:69]
  assign notCDom_nearNormDist = {notCDom_normDistReduced2, 1'h0}; // @[MulAddRecFN.scala 242:56]
  assign _notCDom_sExp_T = {1'b0,$signed(notCDom_nearNormDist)}; // @[MulAddRecFN.scala 243:69]
  assign _GEN_4 = {{3{_notCDom_sExp_T[6]}},_notCDom_sExp_T}; // @[MulAddRecFN.scala 243:46]
  assign notCDom_sExp = $signed(io_fromPreMul_sExpSum) - $signed(_GEN_4); // @[MulAddRecFN.scala 243:46]
  assign _GEN_5 = {{63'd0}, notCDom_absSigSum}; // @[MulAddRecFN.scala 245:27]
  assign _notCDom_mainSig_T = _GEN_5 << notCDom_nearNormDist; // @[MulAddRecFN.scala 245:27]
  assign notCDom_mainSig = _notCDom_mainSig_T[51:23]; // @[MulAddRecFN.scala 245:50]
  assign notCDom_reduced4SigExtra_reducedVec_0 = |notCDom_reduced2AbsSigSum[1:0]; // @[primitives.scala 104:54]
  assign notCDom_reduced4SigExtra_reducedVec_1 = |notCDom_reduced2AbsSigSum[3:2]; // @[primitives.scala 104:54]
  assign notCDom_reduced4SigExtra_reducedVec_2 = |notCDom_reduced2AbsSigSum[5:4]; // @[primitives.scala 104:54]
  assign notCDom_reduced4SigExtra_reducedVec_3 = |notCDom_reduced2AbsSigSum[7:6]; // @[primitives.scala 104:54]
  assign notCDom_reduced4SigExtra_reducedVec_4 = |notCDom_reduced2AbsSigSum[9:8]; // @[primitives.scala 104:54]
  assign notCDom_reduced4SigExtra_reducedVec_5 = |notCDom_reduced2AbsSigSum[11:10]; // @[primitives.scala 104:54]
  assign notCDom_reduced4SigExtra_reducedVec_6 = |notCDom_reduced2AbsSigSum[12]; // @[primitives.scala 107:57]
  assign _notCDom_reduced4SigExtra_T_2 = {notCDom_reduced4SigExtra_reducedVec_6,notCDom_reduced4SigExtra_reducedVec_5,notCDom_reduced4SigExtra_reducedVec_4,notCDom_reduced4SigExtra_reducedVec_3,notCDom_reduced4SigExtra_reducedVec_2,notCDom_reduced4SigExtra_reducedVec_1,notCDom_reduced4SigExtra_reducedVec_0}; // @[primitives.scala 108:20]
  assign notCDom_reduced4SigExtra_shift = -17'sh10000 >>> ~notCDom_normDistReduced2[4:1]; // @[primitives.scala 77:58]
  assign notCDom_reduced4SigExtra_hi_1 = notCDom_reduced4SigExtra_shift[1]; // @[Bitwise.scala 109:18]
  assign notCDom_reduced4SigExtra_lo_1 = notCDom_reduced4SigExtra_shift[2]; // @[Bitwise.scala 109:44]
  assign notCDom_reduced4SigExtra_hi_3 = notCDom_reduced4SigExtra_shift[3]; // @[Bitwise.scala 109:18]
  assign notCDom_reduced4SigExtra_lo_2 = notCDom_reduced4SigExtra_shift[4]; // @[Bitwise.scala 109:44]
  assign notCDom_reduced4SigExtra_hi_5 = notCDom_reduced4SigExtra_shift[5]; // @[Bitwise.scala 109:18]
  assign notCDom_reduced4SigExtra_lo_4 = notCDom_reduced4SigExtra_shift[6]; // @[Bitwise.scala 109:44]
  assign _notCDom_reduced4SigExtra_T_10 = {notCDom_reduced4SigExtra_hi_1,notCDom_reduced4SigExtra_lo_1,notCDom_reduced4SigExtra_hi_3,notCDom_reduced4SigExtra_lo_2,notCDom_reduced4SigExtra_hi_5,notCDom_reduced4SigExtra_lo_4}; // @[Cat.scala 30:58]
  assign _GEN_6 = {{1'd0}, _notCDom_reduced4SigExtra_T_10}; // @[MulAddRecFN.scala 249:78]
  assign _notCDom_reduced4SigExtra_T_11 = _notCDom_reduced4SigExtra_T_2 & _GEN_6; // @[MulAddRecFN.scala 249:78]
  assign notCDom_reduced4SigExtra = |_notCDom_reduced4SigExtra_T_11; // @[MulAddRecFN.scala 251:11]
  assign notCDom_sig_hi = notCDom_mainSig[28:3]; // @[MulAddRecFN.scala 253:28]
  assign _notCDom_sig_T_1 = |notCDom_mainSig[2:0]; // @[MulAddRecFN.scala 254:35]
  assign notCDom_sig_lo = _notCDom_sig_T_1 | notCDom_reduced4SigExtra; // @[MulAddRecFN.scala 254:39]
  assign notCDom_sig = {notCDom_sig_hi,notCDom_sig_lo}; // @[Cat.scala 30:58]
  assign notCDom_completeCancellation = notCDom_sig[26:25] == 2'h0; // @[MulAddRecFN.scala 257:50]
  assign _notCDom_sign_T = io_fromPreMul_signProd ^ notCDom_signSigSum; // @[MulAddRecFN.scala 261:36]
  assign notCDom_sign = notCDom_completeCancellation ? roundingMode_min : _notCDom_sign_T; // @[MulAddRecFN.scala 259:12]
  assign notNaN_isInfProd = io_fromPreMul_isInfA | io_fromPreMul_isInfB; // @[MulAddRecFN.scala 266:49]
  assign notNaN_isInfOut = notNaN_isInfProd | io_fromPreMul_isInfC; // @[MulAddRecFN.scala 267:44]
  assign _notNaN_addZeros_T = io_fromPreMul_isZeroA | io_fromPreMul_isZeroB; // @[MulAddRecFN.scala 269:32]
  assign notNaN_addZeros = _notNaN_addZeros_T & io_fromPreMul_isZeroC; // @[MulAddRecFN.scala 269:58]
  assign _io_invalidExc_T = io_fromPreMul_isInfA & io_fromPreMul_isZeroB; // @[MulAddRecFN.scala 274:31]
  assign _io_invalidExc_T_1 = io_fromPreMul_isSigNaNAny | _io_invalidExc_T; // @[MulAddRecFN.scala 273:35]
  assign _io_invalidExc_T_2 = io_fromPreMul_isZeroA & io_fromPreMul_isInfB; // @[MulAddRecFN.scala 275:32]
  assign _io_invalidExc_T_3 = _io_invalidExc_T_1 | _io_invalidExc_T_2; // @[MulAddRecFN.scala 274:57]
  assign _io_invalidExc_T_6 = ~io_fromPreMul_isNaNAOrB & notNaN_isInfProd; // @[MulAddRecFN.scala 276:36]
  assign _io_invalidExc_T_7 = _io_invalidExc_T_6 & io_fromPreMul_isInfC; // @[MulAddRecFN.scala 277:61]
  assign _io_invalidExc_T_8 = _io_invalidExc_T_7 & io_fromPreMul_doSubMags; // @[MulAddRecFN.scala 278:35]
  assign _io_rawOut_isZero_T_1 = ~io_fromPreMul_CIsDominant & notCDom_completeCancellation; // @[MulAddRecFN.scala 285:42]
  assign _io_rawOut_sign_T = notNaN_isInfProd & io_fromPreMul_signProd; // @[MulAddRecFN.scala 287:27]
  assign _io_rawOut_sign_T_1 = io_fromPreMul_isInfC & CDom_sign; // @[MulAddRecFN.scala 288:31]
  assign _io_rawOut_sign_T_2 = _io_rawOut_sign_T | _io_rawOut_sign_T_1; // @[MulAddRecFN.scala 287:54]
  assign _io_rawOut_sign_T_4 = notNaN_addZeros & ~roundingMode_min; // @[MulAddRecFN.scala 289:26]
  assign _io_rawOut_sign_T_5 = _io_rawOut_sign_T_4 & io_fromPreMul_signProd; // @[MulAddRecFN.scala 289:48]
  assign _io_rawOut_sign_T_6 = _io_rawOut_sign_T_5 & CDom_sign; // @[MulAddRecFN.scala 290:36]
  assign _io_rawOut_sign_T_7 = _io_rawOut_sign_T_2 | _io_rawOut_sign_T_6; // @[MulAddRecFN.scala 288:43]
  assign _io_rawOut_sign_T_8 = notNaN_addZeros & roundingMode_min; // @[MulAddRecFN.scala 291:26]
  assign _io_rawOut_sign_T_9 = io_fromPreMul_signProd | CDom_sign; // @[MulAddRecFN.scala 292:37]
  assign _io_rawOut_sign_T_10 = _io_rawOut_sign_T_8 & _io_rawOut_sign_T_9; // @[MulAddRecFN.scala 291:46]
  assign _io_rawOut_sign_T_11 = _io_rawOut_sign_T_7 | _io_rawOut_sign_T_10; // @[MulAddRecFN.scala 290:48]
  assign _io_rawOut_sign_T_14 = ~notNaN_isInfOut & ~notNaN_addZeros; // @[MulAddRecFN.scala 293:28]
  assign _io_rawOut_sign_T_15 = io_fromPreMul_CIsDominant ? CDom_sign : notCDom_sign; // @[MulAddRecFN.scala 294:17]
  assign _io_rawOut_sign_T_16 = _io_rawOut_sign_T_14 & _io_rawOut_sign_T_15; // @[MulAddRecFN.scala 293:49]
  assign io_invalidExc = _io_invalidExc_T_3 | _io_invalidExc_T_8; // @[MulAddRecFN.scala 272:19]
  assign io_rawOut_isNaN = io_fromPreMul_isNaNAOrB | io_fromPreMul_isNaNC; // @[MulAddRecFN.scala 280:21]
  assign io_rawOut_isInf = notNaN_isInfProd | io_fromPreMul_isInfC; // @[MulAddRecFN.scala 281:21]
  assign io_rawOut_isZero = notNaN_addZeros | _io_rawOut_isZero_T_1; // @[MulAddRecFN.scala 283:22]
  assign io_rawOut_sign = _io_rawOut_sign_T_11 | _io_rawOut_sign_T_16; // @[MulAddRecFN.scala 286:20]
  assign io_rawOut_sExp = io_fromPreMul_CIsDominant ? $signed(CDom_sExp) : $signed(notCDom_sExp); // @[MulAddRecFN.scala 295:20]
  assign io_rawOut_sig = io_fromPreMul_CIsDominant ? CDom_sig : notCDom_sig; // @[MulAddRecFN.scala 296:19]
  assign MulAddRecFNToRaw_postMul_covSum = 30'h0;
  assign io_covSum = MulAddRecFNToRaw_postMul_covSum;
  assign metaAssert = 1'h0;
endmodule
module RoundAnyRawFNToRecFN_1(
  input         io_in_isZero,
  input         io_in_sign,
  input  [8:0]  io_in_sExp,
  input  [64:0] io_in_sig,
  input  [2:0]  io_roundingMode,
  output [32:0] io_out,
  output [4:0]  io_exceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  roundingMode_near_even; // @[RoundAnyRawFNToRecFN.scala 88:53]
  wire  roundingMode_min; // @[RoundAnyRawFNToRecFN.scala 90:53]
  wire  roundingMode_max; // @[RoundAnyRawFNToRecFN.scala 91:53]
  wire  roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 92:53]
  wire  roundingMode_odd; // @[RoundAnyRawFNToRecFN.scala 93:53]
  wire  _roundMagUp_T; // @[RoundAnyRawFNToRecFN.scala 96:27]
  wire  _roundMagUp_T_2; // @[RoundAnyRawFNToRecFN.scala 96:63]
  wire  roundMagUp; // @[RoundAnyRawFNToRecFN.scala 96:42]
  wire [9:0] _sAdjustedExp_T; // @[RoundAnyRawFNToRecFN.scala 102:25]
  wire [9:0] sAdjustedExp; // @[RoundAnyRawFNToRecFN.scala 104:31]
  wire [25:0] adjustedSig_hi; // @[RoundAnyRawFNToRecFN.scala 114:26]
  wire  adjustedSig_lo; // @[RoundAnyRawFNToRecFN.scala 115:60]
  wire [26:0] adjustedSig; // @[Cat.scala 30:58]
  wire [26:0] _roundPosBit_T; // @[RoundAnyRawFNToRecFN.scala 162:40]
  wire  roundPosBit; // @[RoundAnyRawFNToRecFN.scala 162:56]
  wire [26:0] _anyRoundExtra_T; // @[RoundAnyRawFNToRecFN.scala 163:42]
  wire  anyRoundExtra; // @[RoundAnyRawFNToRecFN.scala 163:62]
  wire  anyRound; // @[RoundAnyRawFNToRecFN.scala 164:36]
  wire  _roundIncr_T; // @[RoundAnyRawFNToRecFN.scala 167:38]
  wire  _roundIncr_T_1; // @[RoundAnyRawFNToRecFN.scala 167:67]
  wire  _roundIncr_T_2; // @[RoundAnyRawFNToRecFN.scala 169:29]
  wire  roundIncr; // @[RoundAnyRawFNToRecFN.scala 168:31]
  wire [26:0] _roundedSig_T; // @[RoundAnyRawFNToRecFN.scala 172:32]
  wire [25:0] _roundedSig_T_2; // @[RoundAnyRawFNToRecFN.scala 172:49]
  wire  _roundedSig_T_3; // @[RoundAnyRawFNToRecFN.scala 173:49]
  wire  _roundedSig_T_5; // @[RoundAnyRawFNToRecFN.scala 173:64]
  wire [25:0] _roundedSig_T_7; // @[RoundAnyRawFNToRecFN.scala 173:25]
  wire [25:0] _roundedSig_T_9; // @[RoundAnyRawFNToRecFN.scala 172:61]
  wire [26:0] _roundedSig_T_11; // @[RoundAnyRawFNToRecFN.scala 178:30]
  wire  _roundedSig_T_13; // @[RoundAnyRawFNToRecFN.scala 179:42]
  wire [25:0] _roundedSig_T_15; // @[RoundAnyRawFNToRecFN.scala 179:24]
  wire [25:0] _GEN_0; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [25:0] _roundedSig_T_16; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [25:0] roundedSig; // @[RoundAnyRawFNToRecFN.scala 171:16]
  wire [2:0] _sRoundedExp_T_1; // @[RoundAnyRawFNToRecFN.scala 183:69]
  wire [9:0] _GEN_1; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [10:0] sRoundedExp; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [8:0] common_expOut; // @[RoundAnyRawFNToRecFN.scala 185:37]
  wire [22:0] common_fractOut; // @[RoundAnyRawFNToRecFN.scala 189:27]
  wire  commonCase; // @[RoundAnyRawFNToRecFN.scala 235:64]
  wire  inexact; // @[RoundAnyRawFNToRecFN.scala 238:43]
  wire [8:0] _expOut_T_1; // @[RoundAnyRawFNToRecFN.scala 251:18]
  wire [8:0] expOut; // @[RoundAnyRawFNToRecFN.scala 250:24]
  wire [22:0] fractOut; // @[RoundAnyRawFNToRecFN.scala 278:12]
  wire [9:0] io_out_hi; // @[Cat.scala 30:58]
  wire [1:0] io_exceptionFlags_lo; // @[Cat.scala 30:58]
  wire [29:0] RoundAnyRawFNToRecFN_1_covSum;
  assign roundingMode_near_even = io_roundingMode == 3'h0; // @[RoundAnyRawFNToRecFN.scala 88:53]
  assign roundingMode_min = io_roundingMode == 3'h2; // @[RoundAnyRawFNToRecFN.scala 90:53]
  assign roundingMode_max = io_roundingMode == 3'h3; // @[RoundAnyRawFNToRecFN.scala 91:53]
  assign roundingMode_near_maxMag = io_roundingMode == 3'h4; // @[RoundAnyRawFNToRecFN.scala 92:53]
  assign roundingMode_odd = io_roundingMode == 3'h6; // @[RoundAnyRawFNToRecFN.scala 93:53]
  assign _roundMagUp_T = roundingMode_min & io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:27]
  assign _roundMagUp_T_2 = roundingMode_max & ~io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:63]
  assign roundMagUp = _roundMagUp_T | _roundMagUp_T_2; // @[RoundAnyRawFNToRecFN.scala 96:42]
  assign _sAdjustedExp_T = $signed(io_in_sExp) + 9'sh80; // @[RoundAnyRawFNToRecFN.scala 102:25]
  assign sAdjustedExp = {1'b0,$signed(_sAdjustedExp_T[8:0])}; // @[RoundAnyRawFNToRecFN.scala 104:31]
  assign adjustedSig_hi = io_in_sig[64:39]; // @[RoundAnyRawFNToRecFN.scala 114:26]
  assign adjustedSig_lo = |io_in_sig[38:0]; // @[RoundAnyRawFNToRecFN.scala 115:60]
  assign adjustedSig = {adjustedSig_hi,adjustedSig_lo}; // @[Cat.scala 30:58]
  assign _roundPosBit_T = adjustedSig & 27'h2; // @[RoundAnyRawFNToRecFN.scala 162:40]
  assign roundPosBit = |_roundPosBit_T; // @[RoundAnyRawFNToRecFN.scala 162:56]
  assign _anyRoundExtra_T = adjustedSig & 27'h1; // @[RoundAnyRawFNToRecFN.scala 163:42]
  assign anyRoundExtra = |_anyRoundExtra_T; // @[RoundAnyRawFNToRecFN.scala 163:62]
  assign anyRound = roundPosBit | anyRoundExtra; // @[RoundAnyRawFNToRecFN.scala 164:36]
  assign _roundIncr_T = roundingMode_near_even | roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 167:38]
  assign _roundIncr_T_1 = _roundIncr_T & roundPosBit; // @[RoundAnyRawFNToRecFN.scala 167:67]
  assign _roundIncr_T_2 = roundMagUp & anyRound; // @[RoundAnyRawFNToRecFN.scala 169:29]
  assign roundIncr = _roundIncr_T_1 | _roundIncr_T_2; // @[RoundAnyRawFNToRecFN.scala 168:31]
  assign _roundedSig_T = adjustedSig | 27'h3; // @[RoundAnyRawFNToRecFN.scala 172:32]
  assign _roundedSig_T_2 = _roundedSig_T[26:2] + 25'h1; // @[RoundAnyRawFNToRecFN.scala 172:49]
  assign _roundedSig_T_3 = roundingMode_near_even & roundPosBit; // @[RoundAnyRawFNToRecFN.scala 173:49]
  assign _roundedSig_T_5 = _roundedSig_T_3 & ~anyRoundExtra; // @[RoundAnyRawFNToRecFN.scala 173:64]
  assign _roundedSig_T_7 = _roundedSig_T_5 ? 26'h1 : 26'h0; // @[RoundAnyRawFNToRecFN.scala 173:25]
  assign _roundedSig_T_9 = _roundedSig_T_2 & ~_roundedSig_T_7; // @[RoundAnyRawFNToRecFN.scala 172:61]
  assign _roundedSig_T_11 = adjustedSig & 27'h7fffffc; // @[RoundAnyRawFNToRecFN.scala 178:30]
  assign _roundedSig_T_13 = roundingMode_odd & anyRound; // @[RoundAnyRawFNToRecFN.scala 179:42]
  assign _roundedSig_T_15 = _roundedSig_T_13 ? 26'h1 : 26'h0; // @[RoundAnyRawFNToRecFN.scala 179:24]
  assign _GEN_0 = {{1'd0}, _roundedSig_T_11[26:2]}; // @[RoundAnyRawFNToRecFN.scala 178:47]
  assign _roundedSig_T_16 = _GEN_0 | _roundedSig_T_15; // @[RoundAnyRawFNToRecFN.scala 178:47]
  assign roundedSig = roundIncr ? _roundedSig_T_9 : _roundedSig_T_16; // @[RoundAnyRawFNToRecFN.scala 171:16]
  assign _sRoundedExp_T_1 = {1'b0,$signed(roundedSig[25:24])}; // @[RoundAnyRawFNToRecFN.scala 183:69]
  assign _GEN_1 = {{7{_sRoundedExp_T_1[2]}},_sRoundedExp_T_1}; // @[RoundAnyRawFNToRecFN.scala 183:40]
  assign sRoundedExp = $signed(sAdjustedExp) + $signed(_GEN_1); // @[RoundAnyRawFNToRecFN.scala 183:40]
  assign common_expOut = sRoundedExp[8:0]; // @[RoundAnyRawFNToRecFN.scala 185:37]
  assign common_fractOut = roundedSig[22:0]; // @[RoundAnyRawFNToRecFN.scala 189:27]
  assign commonCase = ~io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 235:64]
  assign inexact = commonCase & anyRound; // @[RoundAnyRawFNToRecFN.scala 238:43]
  assign _expOut_T_1 = io_in_isZero ? 9'h1c0 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 251:18]
  assign expOut = common_expOut & ~_expOut_T_1; // @[RoundAnyRawFNToRecFN.scala 250:24]
  assign fractOut = io_in_isZero ? 23'h0 : common_fractOut; // @[RoundAnyRawFNToRecFN.scala 278:12]
  assign io_out_hi = {io_in_sign,expOut}; // @[Cat.scala 30:58]
  assign io_exceptionFlags_lo = {1'h0,inexact}; // @[Cat.scala 30:58]
  assign io_out = {io_out_hi,fractOut}; // @[RoundAnyRawFNToRecFN.scala 284:12]
  assign io_exceptionFlags = {3'h0,io_exceptionFlags_lo}; // @[RoundAnyRawFNToRecFN.scala 285:23]
  assign RoundAnyRawFNToRecFN_1_covSum = 30'h0;
  assign io_covSum = RoundAnyRawFNToRecFN_1_covSum;
  assign metaAssert = 1'h0;
endmodule
module RoundAnyRawFNToRecFN_2(
  input         io_in_isZero,
  input         io_in_sign,
  input  [8:0]  io_in_sExp,
  input  [64:0] io_in_sig,
  input  [2:0]  io_roundingMode,
  output [64:0] io_out,
  output [4:0]  io_exceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  roundingMode_near_even; // @[RoundAnyRawFNToRecFN.scala 88:53]
  wire  roundingMode_min; // @[RoundAnyRawFNToRecFN.scala 90:53]
  wire  roundingMode_max; // @[RoundAnyRawFNToRecFN.scala 91:53]
  wire  roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 92:53]
  wire  roundingMode_odd; // @[RoundAnyRawFNToRecFN.scala 93:53]
  wire  _roundMagUp_T; // @[RoundAnyRawFNToRecFN.scala 96:27]
  wire  _roundMagUp_T_2; // @[RoundAnyRawFNToRecFN.scala 96:63]
  wire  roundMagUp; // @[RoundAnyRawFNToRecFN.scala 96:42]
  wire [11:0] _GEN_0; // @[RoundAnyRawFNToRecFN.scala 102:25]
  wire [12:0] _sAdjustedExp_T; // @[RoundAnyRawFNToRecFN.scala 102:25]
  wire [12:0] sAdjustedExp; // @[RoundAnyRawFNToRecFN.scala 104:31]
  wire [54:0] adjustedSig_hi; // @[RoundAnyRawFNToRecFN.scala 114:26]
  wire  adjustedSig_lo; // @[RoundAnyRawFNToRecFN.scala 115:60]
  wire [55:0] adjustedSig; // @[Cat.scala 30:58]
  wire [55:0] _roundPosBit_T; // @[RoundAnyRawFNToRecFN.scala 162:40]
  wire  roundPosBit; // @[RoundAnyRawFNToRecFN.scala 162:56]
  wire [55:0] _anyRoundExtra_T; // @[RoundAnyRawFNToRecFN.scala 163:42]
  wire  anyRoundExtra; // @[RoundAnyRawFNToRecFN.scala 163:62]
  wire  anyRound; // @[RoundAnyRawFNToRecFN.scala 164:36]
  wire  _roundIncr_T; // @[RoundAnyRawFNToRecFN.scala 167:38]
  wire  _roundIncr_T_1; // @[RoundAnyRawFNToRecFN.scala 167:67]
  wire  _roundIncr_T_2; // @[RoundAnyRawFNToRecFN.scala 169:29]
  wire  roundIncr; // @[RoundAnyRawFNToRecFN.scala 168:31]
  wire [55:0] _roundedSig_T; // @[RoundAnyRawFNToRecFN.scala 172:32]
  wire [54:0] _roundedSig_T_2; // @[RoundAnyRawFNToRecFN.scala 172:49]
  wire  _roundedSig_T_3; // @[RoundAnyRawFNToRecFN.scala 173:49]
  wire  _roundedSig_T_5; // @[RoundAnyRawFNToRecFN.scala 173:64]
  wire [54:0] _roundedSig_T_7; // @[RoundAnyRawFNToRecFN.scala 173:25]
  wire [54:0] _roundedSig_T_9; // @[RoundAnyRawFNToRecFN.scala 172:61]
  wire [55:0] _roundedSig_T_11; // @[RoundAnyRawFNToRecFN.scala 178:30]
  wire  _roundedSig_T_13; // @[RoundAnyRawFNToRecFN.scala 179:42]
  wire [54:0] _roundedSig_T_15; // @[RoundAnyRawFNToRecFN.scala 179:24]
  wire [54:0] _GEN_1; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [54:0] _roundedSig_T_16; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [54:0] roundedSig; // @[RoundAnyRawFNToRecFN.scala 171:16]
  wire [2:0] _sRoundedExp_T_1; // @[RoundAnyRawFNToRecFN.scala 183:69]
  wire [12:0] _GEN_2; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [13:0] sRoundedExp; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [11:0] common_expOut; // @[RoundAnyRawFNToRecFN.scala 185:37]
  wire [51:0] common_fractOut; // @[RoundAnyRawFNToRecFN.scala 189:27]
  wire  commonCase; // @[RoundAnyRawFNToRecFN.scala 235:64]
  wire  inexact; // @[RoundAnyRawFNToRecFN.scala 238:43]
  wire [11:0] _expOut_T_1; // @[RoundAnyRawFNToRecFN.scala 251:18]
  wire [11:0] expOut; // @[RoundAnyRawFNToRecFN.scala 250:24]
  wire [51:0] fractOut; // @[RoundAnyRawFNToRecFN.scala 278:12]
  wire [12:0] io_out_hi; // @[Cat.scala 30:58]
  wire [1:0] io_exceptionFlags_lo; // @[Cat.scala 30:58]
  wire [29:0] RoundAnyRawFNToRecFN_2_covSum;
  assign roundingMode_near_even = io_roundingMode == 3'h0; // @[RoundAnyRawFNToRecFN.scala 88:53]
  assign roundingMode_min = io_roundingMode == 3'h2; // @[RoundAnyRawFNToRecFN.scala 90:53]
  assign roundingMode_max = io_roundingMode == 3'h3; // @[RoundAnyRawFNToRecFN.scala 91:53]
  assign roundingMode_near_maxMag = io_roundingMode == 3'h4; // @[RoundAnyRawFNToRecFN.scala 92:53]
  assign roundingMode_odd = io_roundingMode == 3'h6; // @[RoundAnyRawFNToRecFN.scala 93:53]
  assign _roundMagUp_T = roundingMode_min & io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:27]
  assign _roundMagUp_T_2 = roundingMode_max & ~io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:63]
  assign roundMagUp = _roundMagUp_T | _roundMagUp_T_2; // @[RoundAnyRawFNToRecFN.scala 96:42]
  assign _GEN_0 = {{3{io_in_sExp[8]}},io_in_sExp}; // @[RoundAnyRawFNToRecFN.scala 102:25]
  assign _sAdjustedExp_T = $signed(_GEN_0) + 12'sh780; // @[RoundAnyRawFNToRecFN.scala 102:25]
  assign sAdjustedExp = {1'b0,$signed(_sAdjustedExp_T[11:0])}; // @[RoundAnyRawFNToRecFN.scala 104:31]
  assign adjustedSig_hi = io_in_sig[64:10]; // @[RoundAnyRawFNToRecFN.scala 114:26]
  assign adjustedSig_lo = |io_in_sig[9:0]; // @[RoundAnyRawFNToRecFN.scala 115:60]
  assign adjustedSig = {adjustedSig_hi,adjustedSig_lo}; // @[Cat.scala 30:58]
  assign _roundPosBit_T = adjustedSig & 56'h2; // @[RoundAnyRawFNToRecFN.scala 162:40]
  assign roundPosBit = |_roundPosBit_T; // @[RoundAnyRawFNToRecFN.scala 162:56]
  assign _anyRoundExtra_T = adjustedSig & 56'h1; // @[RoundAnyRawFNToRecFN.scala 163:42]
  assign anyRoundExtra = |_anyRoundExtra_T; // @[RoundAnyRawFNToRecFN.scala 163:62]
  assign anyRound = roundPosBit | anyRoundExtra; // @[RoundAnyRawFNToRecFN.scala 164:36]
  assign _roundIncr_T = roundingMode_near_even | roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 167:38]
  assign _roundIncr_T_1 = _roundIncr_T & roundPosBit; // @[RoundAnyRawFNToRecFN.scala 167:67]
  assign _roundIncr_T_2 = roundMagUp & anyRound; // @[RoundAnyRawFNToRecFN.scala 169:29]
  assign roundIncr = _roundIncr_T_1 | _roundIncr_T_2; // @[RoundAnyRawFNToRecFN.scala 168:31]
  assign _roundedSig_T = adjustedSig | 56'h3; // @[RoundAnyRawFNToRecFN.scala 172:32]
  assign _roundedSig_T_2 = _roundedSig_T[55:2] + 54'h1; // @[RoundAnyRawFNToRecFN.scala 172:49]
  assign _roundedSig_T_3 = roundingMode_near_even & roundPosBit; // @[RoundAnyRawFNToRecFN.scala 173:49]
  assign _roundedSig_T_5 = _roundedSig_T_3 & ~anyRoundExtra; // @[RoundAnyRawFNToRecFN.scala 173:64]
  assign _roundedSig_T_7 = _roundedSig_T_5 ? 55'h1 : 55'h0; // @[RoundAnyRawFNToRecFN.scala 173:25]
  assign _roundedSig_T_9 = _roundedSig_T_2 & ~_roundedSig_T_7; // @[RoundAnyRawFNToRecFN.scala 172:61]
  assign _roundedSig_T_11 = adjustedSig & 56'hfffffffffffffc; // @[RoundAnyRawFNToRecFN.scala 178:30]
  assign _roundedSig_T_13 = roundingMode_odd & anyRound; // @[RoundAnyRawFNToRecFN.scala 179:42]
  assign _roundedSig_T_15 = _roundedSig_T_13 ? 55'h1 : 55'h0; // @[RoundAnyRawFNToRecFN.scala 179:24]
  assign _GEN_1 = {{1'd0}, _roundedSig_T_11[55:2]}; // @[RoundAnyRawFNToRecFN.scala 178:47]
  assign _roundedSig_T_16 = _GEN_1 | _roundedSig_T_15; // @[RoundAnyRawFNToRecFN.scala 178:47]
  assign roundedSig = roundIncr ? _roundedSig_T_9 : _roundedSig_T_16; // @[RoundAnyRawFNToRecFN.scala 171:16]
  assign _sRoundedExp_T_1 = {1'b0,$signed(roundedSig[54:53])}; // @[RoundAnyRawFNToRecFN.scala 183:69]
  assign _GEN_2 = {{10{_sRoundedExp_T_1[2]}},_sRoundedExp_T_1}; // @[RoundAnyRawFNToRecFN.scala 183:40]
  assign sRoundedExp = $signed(sAdjustedExp) + $signed(_GEN_2); // @[RoundAnyRawFNToRecFN.scala 183:40]
  assign common_expOut = sRoundedExp[11:0]; // @[RoundAnyRawFNToRecFN.scala 185:37]
  assign common_fractOut = roundedSig[51:0]; // @[RoundAnyRawFNToRecFN.scala 189:27]
  assign commonCase = ~io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 235:64]
  assign inexact = commonCase & anyRound; // @[RoundAnyRawFNToRecFN.scala 238:43]
  assign _expOut_T_1 = io_in_isZero ? 12'he00 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 251:18]
  assign expOut = common_expOut & ~_expOut_T_1; // @[RoundAnyRawFNToRecFN.scala 250:24]
  assign fractOut = io_in_isZero ? 52'h0 : common_fractOut; // @[RoundAnyRawFNToRecFN.scala 278:12]
  assign io_out_hi = {io_in_sign,expOut}; // @[Cat.scala 30:58]
  assign io_exceptionFlags_lo = {1'h0,inexact}; // @[Cat.scala 30:58]
  assign io_out = {io_out_hi,fractOut}; // @[RoundAnyRawFNToRecFN.scala 284:12]
  assign io_exceptionFlags = {3'h0,io_exceptionFlags_lo}; // @[RoundAnyRawFNToRecFN.scala 285:23]
  assign RoundAnyRawFNToRecFN_2_covSum = 30'h0;
  assign io_covSum = RoundAnyRawFNToRecFN_2_covSum;
  assign metaAssert = 1'h0;
endmodule
module RoundAnyRawFNToRecFN_3(
  input         io_invalidExc,
  input         io_in_isNaN,
  input         io_in_isInf,
  input         io_in_isZero,
  input         io_in_sign,
  input  [12:0] io_in_sExp,
  input  [53:0] io_in_sig,
  input  [2:0]  io_roundingMode,
  output [32:0] io_out,
  output [4:0]  io_exceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  roundingMode_near_even; // @[RoundAnyRawFNToRecFN.scala 88:53]
  wire  roundingMode_min; // @[RoundAnyRawFNToRecFN.scala 90:53]
  wire  roundingMode_max; // @[RoundAnyRawFNToRecFN.scala 91:53]
  wire  roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 92:53]
  wire  roundingMode_odd; // @[RoundAnyRawFNToRecFN.scala 93:53]
  wire  _roundMagUp_T; // @[RoundAnyRawFNToRecFN.scala 96:27]
  wire  _roundMagUp_T_2; // @[RoundAnyRawFNToRecFN.scala 96:63]
  wire  roundMagUp; // @[RoundAnyRawFNToRecFN.scala 96:42]
  wire [13:0] sAdjustedExp; // @[RoundAnyRawFNToRecFN.scala 108:24]
  wire [25:0] adjustedSig_hi; // @[RoundAnyRawFNToRecFN.scala 114:26]
  wire  adjustedSig_lo; // @[RoundAnyRawFNToRecFN.scala 115:60]
  wire [26:0] adjustedSig; // @[Cat.scala 30:58]
  wire  roundMask_msb; // @[primitives.scala 57:25]
  wire [7:0] roundMask_lsbs; // @[primitives.scala 58:26]
  wire  roundMask_msb_1; // @[primitives.scala 57:25]
  wire [6:0] roundMask_lsbs_1; // @[primitives.scala 58:26]
  wire  roundMask_msb_2; // @[primitives.scala 57:25]
  wire [5:0] roundMask_lsbs_2; // @[primitives.scala 58:26]
  wire [64:0] roundMask_shift; // @[primitives.scala 77:58]
  wire [15:0] _roundMask_T_7; // @[Bitwise.scala 103:31]
  wire [15:0] _roundMask_T_9; // @[Bitwise.scala 103:65]
  wire [15:0] _roundMask_T_11; // @[Bitwise.scala 103:75]
  wire [15:0] _roundMask_T_12; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_0; // @[Bitwise.scala 103:31]
  wire [15:0] _roundMask_T_17; // @[Bitwise.scala 103:31]
  wire [15:0] _roundMask_T_19; // @[Bitwise.scala 103:65]
  wire [15:0] _roundMask_T_21; // @[Bitwise.scala 103:75]
  wire [15:0] _roundMask_T_22; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_1; // @[Bitwise.scala 103:31]
  wire [15:0] _roundMask_T_27; // @[Bitwise.scala 103:31]
  wire [15:0] _roundMask_T_29; // @[Bitwise.scala 103:65]
  wire [15:0] _roundMask_T_31; // @[Bitwise.scala 103:75]
  wire [15:0] _roundMask_T_32; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_2; // @[Bitwise.scala 103:31]
  wire [15:0] _roundMask_T_37; // @[Bitwise.scala 103:31]
  wire [15:0] _roundMask_T_39; // @[Bitwise.scala 103:65]
  wire [15:0] _roundMask_T_41; // @[Bitwise.scala 103:75]
  wire [15:0] roundMask_hi; // @[Bitwise.scala 103:39]
  wire  roundMask_hi_1; // @[Bitwise.scala 109:18]
  wire  roundMask_lo; // @[Bitwise.scala 109:44]
  wire  roundMask_hi_3; // @[Bitwise.scala 109:18]
  wire  roundMask_lo_1; // @[Bitwise.scala 109:44]
  wire  roundMask_hi_5; // @[Bitwise.scala 109:18]
  wire  roundMask_lo_3; // @[Bitwise.scala 109:44]
  wire [21:0] _roundMask_T_47; // @[Cat.scala 30:58]
  wire [21:0] _roundMask_T_49; // @[primitives.scala 74:21]
  wire [21:0] roundMask_hi_6; // @[primitives.scala 74:17]
  wire [24:0] _roundMask_T_50; // @[Cat.scala 30:58]
  wire  roundMask_hi_7; // @[Bitwise.scala 109:18]
  wire  roundMask_lo_6; // @[Bitwise.scala 109:44]
  wire  roundMask_lo_7; // @[Bitwise.scala 109:44]
  wire [2:0] _roundMask_T_53; // @[Cat.scala 30:58]
  wire [2:0] _roundMask_T_54; // @[primitives.scala 61:24]
  wire [24:0] _roundMask_T_55; // @[primitives.scala 66:24]
  wire [24:0] roundMask_hi_9; // @[primitives.scala 61:24]
  wire [26:0] roundMask; // @[Cat.scala 30:58]
  wire [25:0] shiftedRoundMask_lo; // @[RoundAnyRawFNToRecFN.scala 160:57]
  wire [26:0] shiftedRoundMask; // @[Cat.scala 30:58]
  wire [26:0] roundPosMask; // @[RoundAnyRawFNToRecFN.scala 161:46]
  wire [26:0] _roundPosBit_T; // @[RoundAnyRawFNToRecFN.scala 162:40]
  wire  roundPosBit; // @[RoundAnyRawFNToRecFN.scala 162:56]
  wire [26:0] _anyRoundExtra_T; // @[RoundAnyRawFNToRecFN.scala 163:42]
  wire  anyRoundExtra; // @[RoundAnyRawFNToRecFN.scala 163:62]
  wire  anyRound; // @[RoundAnyRawFNToRecFN.scala 164:36]
  wire  _roundIncr_T; // @[RoundAnyRawFNToRecFN.scala 167:38]
  wire  _roundIncr_T_1; // @[RoundAnyRawFNToRecFN.scala 167:67]
  wire  _roundIncr_T_2; // @[RoundAnyRawFNToRecFN.scala 169:29]
  wire  roundIncr; // @[RoundAnyRawFNToRecFN.scala 168:31]
  wire [26:0] _roundedSig_T; // @[RoundAnyRawFNToRecFN.scala 172:32]
  wire [25:0] _roundedSig_T_2; // @[RoundAnyRawFNToRecFN.scala 172:49]
  wire  _roundedSig_T_3; // @[RoundAnyRawFNToRecFN.scala 173:49]
  wire  _roundedSig_T_5; // @[RoundAnyRawFNToRecFN.scala 173:64]
  wire [25:0] _roundedSig_T_7; // @[RoundAnyRawFNToRecFN.scala 173:25]
  wire [25:0] _roundedSig_T_9; // @[RoundAnyRawFNToRecFN.scala 172:61]
  wire [26:0] _roundedSig_T_11; // @[RoundAnyRawFNToRecFN.scala 178:30]
  wire  _roundedSig_T_13; // @[RoundAnyRawFNToRecFN.scala 179:42]
  wire [25:0] _roundedSig_T_15; // @[RoundAnyRawFNToRecFN.scala 179:24]
  wire [25:0] _GEN_3; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [25:0] _roundedSig_T_16; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [25:0] roundedSig; // @[RoundAnyRawFNToRecFN.scala 171:16]
  wire [2:0] _sRoundedExp_T_1; // @[RoundAnyRawFNToRecFN.scala 183:69]
  wire [13:0] _GEN_4; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [14:0] sRoundedExp; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [8:0] common_expOut; // @[RoundAnyRawFNToRecFN.scala 185:37]
  wire [22:0] common_fractOut; // @[RoundAnyRawFNToRecFN.scala 189:27]
  wire [7:0] _common_overflow_T; // @[RoundAnyRawFNToRecFN.scala 194:30]
  wire  common_overflow; // @[RoundAnyRawFNToRecFN.scala 194:50]
  wire  common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 198:31]
  wire  unboundedRange_roundPosBit; // @[RoundAnyRawFNToRecFN.scala 201:61]
  wire  unboundedRange_anyRound; // @[RoundAnyRawFNToRecFN.scala 203:70]
  wire  _unboundedRange_roundIncr_T_1; // @[RoundAnyRawFNToRecFN.scala 205:67]
  wire  _unboundedRange_roundIncr_T_2; // @[RoundAnyRawFNToRecFN.scala 207:29]
  wire  unboundedRange_roundIncr; // @[RoundAnyRawFNToRecFN.scala 206:46]
  wire  roundCarry; // @[RoundAnyRawFNToRecFN.scala 211:27]
  wire [5:0] _common_underflow_T; // @[RoundAnyRawFNToRecFN.scala 218:48]
  wire  _common_underflow_T_1; // @[RoundAnyRawFNToRecFN.scala 218:62]
  wire  _common_underflow_T_2; // @[RoundAnyRawFNToRecFN.scala 218:32]
  wire  _common_underflow_T_6; // @[RoundAnyRawFNToRecFN.scala 218:74]
  wire  _common_underflow_T_13; // @[RoundAnyRawFNToRecFN.scala 224:38]
  wire  _common_underflow_T_14; // @[RoundAnyRawFNToRecFN.scala 225:45]
  wire  _common_underflow_T_15; // @[RoundAnyRawFNToRecFN.scala 225:60]
  wire  _common_underflow_T_17; // @[RoundAnyRawFNToRecFN.scala 219:76]
  wire  common_underflow; // @[RoundAnyRawFNToRecFN.scala 215:40]
  wire  common_inexact; // @[RoundAnyRawFNToRecFN.scala 228:49]
  wire  isNaNOut; // @[RoundAnyRawFNToRecFN.scala 233:34]
  wire  _commonCase_T_2; // @[RoundAnyRawFNToRecFN.scala 235:33]
  wire  commonCase; // @[RoundAnyRawFNToRecFN.scala 235:61]
  wire  overflow; // @[RoundAnyRawFNToRecFN.scala 236:32]
  wire  underflow; // @[RoundAnyRawFNToRecFN.scala 237:32]
  wire  _inexact_T; // @[RoundAnyRawFNToRecFN.scala 238:43]
  wire  inexact; // @[RoundAnyRawFNToRecFN.scala 238:28]
  wire  overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 241:60]
  wire  _pegMinNonzeroMagOut_T; // @[RoundAnyRawFNToRecFN.scala 243:20]
  wire  _pegMinNonzeroMagOut_T_1; // @[RoundAnyRawFNToRecFN.scala 243:60]
  wire  pegMinNonzeroMagOut; // @[RoundAnyRawFNToRecFN.scala 243:45]
  wire  pegMaxFiniteMagOut; // @[RoundAnyRawFNToRecFN.scala 244:39]
  wire  _notNaN_isInfOut_T; // @[RoundAnyRawFNToRecFN.scala 246:45]
  wire  notNaN_isInfOut; // @[RoundAnyRawFNToRecFN.scala 246:32]
  wire  signOut; // @[RoundAnyRawFNToRecFN.scala 248:22]
  wire  _expOut_T; // @[RoundAnyRawFNToRecFN.scala 251:32]
  wire [8:0] _expOut_T_1; // @[RoundAnyRawFNToRecFN.scala 251:18]
  wire [8:0] _expOut_T_3; // @[RoundAnyRawFNToRecFN.scala 250:24]
  wire [8:0] _expOut_T_5; // @[RoundAnyRawFNToRecFN.scala 255:18]
  wire [8:0] _expOut_T_7; // @[RoundAnyRawFNToRecFN.scala 254:17]
  wire [8:0] _expOut_T_8; // @[RoundAnyRawFNToRecFN.scala 259:18]
  wire [8:0] _expOut_T_10; // @[RoundAnyRawFNToRecFN.scala 258:17]
  wire [8:0] _expOut_T_11; // @[RoundAnyRawFNToRecFN.scala 263:18]
  wire [8:0] _expOut_T_13; // @[RoundAnyRawFNToRecFN.scala 262:17]
  wire [8:0] _expOut_T_14; // @[RoundAnyRawFNToRecFN.scala 267:16]
  wire [8:0] _expOut_T_15; // @[RoundAnyRawFNToRecFN.scala 266:18]
  wire [8:0] _expOut_T_16; // @[RoundAnyRawFNToRecFN.scala 271:16]
  wire [8:0] _expOut_T_17; // @[RoundAnyRawFNToRecFN.scala 270:15]
  wire [8:0] _expOut_T_18; // @[RoundAnyRawFNToRecFN.scala 275:16]
  wire [8:0] _expOut_T_19; // @[RoundAnyRawFNToRecFN.scala 274:15]
  wire [8:0] _expOut_T_20; // @[RoundAnyRawFNToRecFN.scala 276:16]
  wire [8:0] expOut; // @[RoundAnyRawFNToRecFN.scala 275:77]
  wire  _fractOut_T; // @[RoundAnyRawFNToRecFN.scala 278:22]
  wire  _fractOut_T_1; // @[RoundAnyRawFNToRecFN.scala 278:38]
  wire [22:0] _fractOut_T_2; // @[RoundAnyRawFNToRecFN.scala 279:16]
  wire [22:0] _fractOut_T_3; // @[RoundAnyRawFNToRecFN.scala 278:12]
  wire [22:0] _fractOut_T_5; // @[Bitwise.scala 72:12]
  wire [22:0] fractOut; // @[RoundAnyRawFNToRecFN.scala 281:11]
  wire [9:0] io_out_hi; // @[Cat.scala 30:58]
  wire [1:0] io_exceptionFlags_lo; // @[Cat.scala 30:58]
  wire [2:0] io_exceptionFlags_hi; // @[Cat.scala 30:58]
  wire [29:0] RoundAnyRawFNToRecFN_3_covSum;
  assign roundingMode_near_even = io_roundingMode == 3'h0; // @[RoundAnyRawFNToRecFN.scala 88:53]
  assign roundingMode_min = io_roundingMode == 3'h2; // @[RoundAnyRawFNToRecFN.scala 90:53]
  assign roundingMode_max = io_roundingMode == 3'h3; // @[RoundAnyRawFNToRecFN.scala 91:53]
  assign roundingMode_near_maxMag = io_roundingMode == 3'h4; // @[RoundAnyRawFNToRecFN.scala 92:53]
  assign roundingMode_odd = io_roundingMode == 3'h6; // @[RoundAnyRawFNToRecFN.scala 93:53]
  assign _roundMagUp_T = roundingMode_min & io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:27]
  assign _roundMagUp_T_2 = roundingMode_max & ~io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:63]
  assign roundMagUp = _roundMagUp_T | _roundMagUp_T_2; // @[RoundAnyRawFNToRecFN.scala 96:42]
  assign sAdjustedExp = $signed(io_in_sExp) + $signed(-13'sh700); // @[RoundAnyRawFNToRecFN.scala 108:24]
  assign adjustedSig_hi = io_in_sig[53:28]; // @[RoundAnyRawFNToRecFN.scala 114:26]
  assign adjustedSig_lo = |io_in_sig[27:0]; // @[RoundAnyRawFNToRecFN.scala 115:60]
  assign adjustedSig = {adjustedSig_hi,adjustedSig_lo}; // @[Cat.scala 30:58]
  assign roundMask_msb = ~sAdjustedExp[8]; // @[primitives.scala 57:25]
  assign roundMask_lsbs = ~sAdjustedExp[7:0]; // @[primitives.scala 58:26]
  assign roundMask_msb_1 = roundMask_lsbs[7]; // @[primitives.scala 57:25]
  assign roundMask_lsbs_1 = roundMask_lsbs[6:0]; // @[primitives.scala 58:26]
  assign roundMask_msb_2 = roundMask_lsbs_1[6]; // @[primitives.scala 57:25]
  assign roundMask_lsbs_2 = roundMask_lsbs_1[5:0]; // @[primitives.scala 58:26]
  assign roundMask_shift = -65'sh10000000000000000 >>> roundMask_lsbs_2; // @[primitives.scala 77:58]
  assign _roundMask_T_7 = {{8'd0}, roundMask_shift[57:50]}; // @[Bitwise.scala 103:31]
  assign _roundMask_T_9 = {roundMask_shift[49:42], 8'h0}; // @[Bitwise.scala 103:65]
  assign _roundMask_T_11 = _roundMask_T_9 & 16'hff00; // @[Bitwise.scala 103:75]
  assign _roundMask_T_12 = _roundMask_T_7 | _roundMask_T_11; // @[Bitwise.scala 103:39]
  assign _GEN_0 = {{4'd0}, _roundMask_T_12[15:4]}; // @[Bitwise.scala 103:31]
  assign _roundMask_T_17 = _GEN_0 & 16'hf0f; // @[Bitwise.scala 103:31]
  assign _roundMask_T_19 = {_roundMask_T_12[11:0], 4'h0}; // @[Bitwise.scala 103:65]
  assign _roundMask_T_21 = _roundMask_T_19 & 16'hf0f0; // @[Bitwise.scala 103:75]
  assign _roundMask_T_22 = _roundMask_T_17 | _roundMask_T_21; // @[Bitwise.scala 103:39]
  assign _GEN_1 = {{2'd0}, _roundMask_T_22[15:2]}; // @[Bitwise.scala 103:31]
  assign _roundMask_T_27 = _GEN_1 & 16'h3333; // @[Bitwise.scala 103:31]
  assign _roundMask_T_29 = {_roundMask_T_22[13:0], 2'h0}; // @[Bitwise.scala 103:65]
  assign _roundMask_T_31 = _roundMask_T_29 & 16'hcccc; // @[Bitwise.scala 103:75]
  assign _roundMask_T_32 = _roundMask_T_27 | _roundMask_T_31; // @[Bitwise.scala 103:39]
  assign _GEN_2 = {{1'd0}, _roundMask_T_32[15:1]}; // @[Bitwise.scala 103:31]
  assign _roundMask_T_37 = _GEN_2 & 16'h5555; // @[Bitwise.scala 103:31]
  assign _roundMask_T_39 = {_roundMask_T_32[14:0], 1'h0}; // @[Bitwise.scala 103:65]
  assign _roundMask_T_41 = _roundMask_T_39 & 16'haaaa; // @[Bitwise.scala 103:75]
  assign roundMask_hi = _roundMask_T_37 | _roundMask_T_41; // @[Bitwise.scala 103:39]
  assign roundMask_hi_1 = roundMask_shift[58]; // @[Bitwise.scala 109:18]
  assign roundMask_lo = roundMask_shift[59]; // @[Bitwise.scala 109:44]
  assign roundMask_hi_3 = roundMask_shift[60]; // @[Bitwise.scala 109:18]
  assign roundMask_lo_1 = roundMask_shift[61]; // @[Bitwise.scala 109:44]
  assign roundMask_hi_5 = roundMask_shift[62]; // @[Bitwise.scala 109:18]
  assign roundMask_lo_3 = roundMask_shift[63]; // @[Bitwise.scala 109:44]
  assign _roundMask_T_47 = {roundMask_hi,roundMask_hi_1,roundMask_lo,roundMask_hi_3,roundMask_lo_1,roundMask_hi_5,roundMask_lo_3}; // @[Cat.scala 30:58]
  assign _roundMask_T_49 = roundMask_msb_2 ? 22'h0 : ~_roundMask_T_47; // @[primitives.scala 74:21]
  assign roundMask_hi_6 = ~_roundMask_T_49; // @[primitives.scala 74:17]
  assign _roundMask_T_50 = {roundMask_hi_6,3'h7}; // @[Cat.scala 30:58]
  assign roundMask_hi_7 = roundMask_shift[0]; // @[Bitwise.scala 109:18]
  assign roundMask_lo_6 = roundMask_shift[1]; // @[Bitwise.scala 109:44]
  assign roundMask_lo_7 = roundMask_shift[2]; // @[Bitwise.scala 109:44]
  assign _roundMask_T_53 = {roundMask_hi_7,roundMask_lo_6,roundMask_lo_7}; // @[Cat.scala 30:58]
  assign _roundMask_T_54 = roundMask_msb_2 ? _roundMask_T_53 : 3'h0; // @[primitives.scala 61:24]
  assign _roundMask_T_55 = roundMask_msb_1 ? _roundMask_T_50 : {{22'd0}, _roundMask_T_54}; // @[primitives.scala 66:24]
  assign roundMask_hi_9 = roundMask_msb ? _roundMask_T_55 : 25'h0; // @[primitives.scala 61:24]
  assign roundMask = {roundMask_hi_9,2'h3}; // @[Cat.scala 30:58]
  assign shiftedRoundMask_lo = roundMask[26:1]; // @[RoundAnyRawFNToRecFN.scala 160:57]
  assign shiftedRoundMask = {1'h0,shiftedRoundMask_lo}; // @[Cat.scala 30:58]
  assign roundPosMask = ~shiftedRoundMask & roundMask; // @[RoundAnyRawFNToRecFN.scala 161:46]
  assign _roundPosBit_T = adjustedSig & roundPosMask; // @[RoundAnyRawFNToRecFN.scala 162:40]
  assign roundPosBit = |_roundPosBit_T; // @[RoundAnyRawFNToRecFN.scala 162:56]
  assign _anyRoundExtra_T = adjustedSig & shiftedRoundMask; // @[RoundAnyRawFNToRecFN.scala 163:42]
  assign anyRoundExtra = |_anyRoundExtra_T; // @[RoundAnyRawFNToRecFN.scala 163:62]
  assign anyRound = roundPosBit | anyRoundExtra; // @[RoundAnyRawFNToRecFN.scala 164:36]
  assign _roundIncr_T = roundingMode_near_even | roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 167:38]
  assign _roundIncr_T_1 = _roundIncr_T & roundPosBit; // @[RoundAnyRawFNToRecFN.scala 167:67]
  assign _roundIncr_T_2 = roundMagUp & anyRound; // @[RoundAnyRawFNToRecFN.scala 169:29]
  assign roundIncr = _roundIncr_T_1 | _roundIncr_T_2; // @[RoundAnyRawFNToRecFN.scala 168:31]
  assign _roundedSig_T = adjustedSig | roundMask; // @[RoundAnyRawFNToRecFN.scala 172:32]
  assign _roundedSig_T_2 = _roundedSig_T[26:2] + 25'h1; // @[RoundAnyRawFNToRecFN.scala 172:49]
  assign _roundedSig_T_3 = roundingMode_near_even & roundPosBit; // @[RoundAnyRawFNToRecFN.scala 173:49]
  assign _roundedSig_T_5 = _roundedSig_T_3 & ~anyRoundExtra; // @[RoundAnyRawFNToRecFN.scala 173:64]
  assign _roundedSig_T_7 = _roundedSig_T_5 ? shiftedRoundMask_lo : 26'h0; // @[RoundAnyRawFNToRecFN.scala 173:25]
  assign _roundedSig_T_9 = _roundedSig_T_2 & ~_roundedSig_T_7; // @[RoundAnyRawFNToRecFN.scala 172:61]
  assign _roundedSig_T_11 = adjustedSig & ~roundMask; // @[RoundAnyRawFNToRecFN.scala 178:30]
  assign _roundedSig_T_13 = roundingMode_odd & anyRound; // @[RoundAnyRawFNToRecFN.scala 179:42]
  assign _roundedSig_T_15 = _roundedSig_T_13 ? roundPosMask[26:1] : 26'h0; // @[RoundAnyRawFNToRecFN.scala 179:24]
  assign _GEN_3 = {{1'd0}, _roundedSig_T_11[26:2]}; // @[RoundAnyRawFNToRecFN.scala 178:47]
  assign _roundedSig_T_16 = _GEN_3 | _roundedSig_T_15; // @[RoundAnyRawFNToRecFN.scala 178:47]
  assign roundedSig = roundIncr ? _roundedSig_T_9 : _roundedSig_T_16; // @[RoundAnyRawFNToRecFN.scala 171:16]
  assign _sRoundedExp_T_1 = {1'b0,$signed(roundedSig[25:24])}; // @[RoundAnyRawFNToRecFN.scala 183:69]
  assign _GEN_4 = {{11{_sRoundedExp_T_1[2]}},_sRoundedExp_T_1}; // @[RoundAnyRawFNToRecFN.scala 183:40]
  assign sRoundedExp = $signed(sAdjustedExp) + $signed(_GEN_4); // @[RoundAnyRawFNToRecFN.scala 183:40]
  assign common_expOut = sRoundedExp[8:0]; // @[RoundAnyRawFNToRecFN.scala 185:37]
  assign common_fractOut = roundedSig[22:0]; // @[RoundAnyRawFNToRecFN.scala 189:27]
  assign _common_overflow_T = sRoundedExp[14:7]; // @[RoundAnyRawFNToRecFN.scala 194:30]
  assign common_overflow = $signed(_common_overflow_T) >= 8'sh3; // @[RoundAnyRawFNToRecFN.scala 194:50]
  assign common_totalUnderflow = $signed(sRoundedExp) < 15'sh6b; // @[RoundAnyRawFNToRecFN.scala 198:31]
  assign unboundedRange_roundPosBit = adjustedSig[1]; // @[RoundAnyRawFNToRecFN.scala 201:61]
  assign unboundedRange_anyRound = |adjustedSig[1:0]; // @[RoundAnyRawFNToRecFN.scala 203:70]
  assign _unboundedRange_roundIncr_T_1 = _roundIncr_T & unboundedRange_roundPosBit; // @[RoundAnyRawFNToRecFN.scala 205:67]
  assign _unboundedRange_roundIncr_T_2 = roundMagUp & unboundedRange_anyRound; // @[RoundAnyRawFNToRecFN.scala 207:29]
  assign unboundedRange_roundIncr = _unboundedRange_roundIncr_T_1 | _unboundedRange_roundIncr_T_2; // @[RoundAnyRawFNToRecFN.scala 206:46]
  assign roundCarry = roundedSig[24]; // @[RoundAnyRawFNToRecFN.scala 211:27]
  assign _common_underflow_T = sAdjustedExp[13:8]; // @[RoundAnyRawFNToRecFN.scala 218:48]
  assign _common_underflow_T_1 = $signed(_common_underflow_T) <= 6'sh0; // @[RoundAnyRawFNToRecFN.scala 218:62]
  assign _common_underflow_T_2 = anyRound & _common_underflow_T_1; // @[RoundAnyRawFNToRecFN.scala 218:32]
  assign _common_underflow_T_6 = _common_underflow_T_2 & roundMask[2]; // @[RoundAnyRawFNToRecFN.scala 218:74]
  assign _common_underflow_T_13 = ~roundMask[3] & roundCarry; // @[RoundAnyRawFNToRecFN.scala 224:38]
  assign _common_underflow_T_14 = _common_underflow_T_13 & roundPosBit; // @[RoundAnyRawFNToRecFN.scala 225:45]
  assign _common_underflow_T_15 = _common_underflow_T_14 & unboundedRange_roundIncr; // @[RoundAnyRawFNToRecFN.scala 225:60]
  assign _common_underflow_T_17 = _common_underflow_T_6 & ~_common_underflow_T_15; // @[RoundAnyRawFNToRecFN.scala 219:76]
  assign common_underflow = common_totalUnderflow | _common_underflow_T_17; // @[RoundAnyRawFNToRecFN.scala 215:40]
  assign common_inexact = common_totalUnderflow | anyRound; // @[RoundAnyRawFNToRecFN.scala 228:49]
  assign isNaNOut = io_invalidExc | io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 233:34]
  assign _commonCase_T_2 = ~isNaNOut & ~io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 235:33]
  assign commonCase = _commonCase_T_2 & ~io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 235:61]
  assign overflow = commonCase & common_overflow; // @[RoundAnyRawFNToRecFN.scala 236:32]
  assign underflow = commonCase & common_underflow; // @[RoundAnyRawFNToRecFN.scala 237:32]
  assign _inexact_T = commonCase & common_inexact; // @[RoundAnyRawFNToRecFN.scala 238:43]
  assign inexact = overflow | _inexact_T; // @[RoundAnyRawFNToRecFN.scala 238:28]
  assign overflow_roundMagUp = _roundIncr_T | roundMagUp; // @[RoundAnyRawFNToRecFN.scala 241:60]
  assign _pegMinNonzeroMagOut_T = commonCase & common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 243:20]
  assign _pegMinNonzeroMagOut_T_1 = roundMagUp | roundingMode_odd; // @[RoundAnyRawFNToRecFN.scala 243:60]
  assign pegMinNonzeroMagOut = _pegMinNonzeroMagOut_T & _pegMinNonzeroMagOut_T_1; // @[RoundAnyRawFNToRecFN.scala 243:45]
  assign pegMaxFiniteMagOut = overflow & ~overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 244:39]
  assign _notNaN_isInfOut_T = overflow & overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 246:45]
  assign notNaN_isInfOut = io_in_isInf | _notNaN_isInfOut_T; // @[RoundAnyRawFNToRecFN.scala 246:32]
  assign signOut = isNaNOut ? 1'h0 : io_in_sign; // @[RoundAnyRawFNToRecFN.scala 248:22]
  assign _expOut_T = io_in_isZero | common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 251:32]
  assign _expOut_T_1 = _expOut_T ? 9'h1c0 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 251:18]
  assign _expOut_T_3 = common_expOut & ~_expOut_T_1; // @[RoundAnyRawFNToRecFN.scala 250:24]
  assign _expOut_T_5 = pegMinNonzeroMagOut ? 9'h194 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 255:18]
  assign _expOut_T_7 = _expOut_T_3 & ~_expOut_T_5; // @[RoundAnyRawFNToRecFN.scala 254:17]
  assign _expOut_T_8 = pegMaxFiniteMagOut ? 9'h80 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 259:18]
  assign _expOut_T_10 = _expOut_T_7 & ~_expOut_T_8; // @[RoundAnyRawFNToRecFN.scala 258:17]
  assign _expOut_T_11 = notNaN_isInfOut ? 9'h40 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 263:18]
  assign _expOut_T_13 = _expOut_T_10 & ~_expOut_T_11; // @[RoundAnyRawFNToRecFN.scala 262:17]
  assign _expOut_T_14 = pegMinNonzeroMagOut ? 9'h6b : 9'h0; // @[RoundAnyRawFNToRecFN.scala 267:16]
  assign _expOut_T_15 = _expOut_T_13 | _expOut_T_14; // @[RoundAnyRawFNToRecFN.scala 266:18]
  assign _expOut_T_16 = pegMaxFiniteMagOut ? 9'h17f : 9'h0; // @[RoundAnyRawFNToRecFN.scala 271:16]
  assign _expOut_T_17 = _expOut_T_15 | _expOut_T_16; // @[RoundAnyRawFNToRecFN.scala 270:15]
  assign _expOut_T_18 = notNaN_isInfOut ? 9'h180 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 275:16]
  assign _expOut_T_19 = _expOut_T_17 | _expOut_T_18; // @[RoundAnyRawFNToRecFN.scala 274:15]
  assign _expOut_T_20 = isNaNOut ? 9'h1c0 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 276:16]
  assign expOut = _expOut_T_19 | _expOut_T_20; // @[RoundAnyRawFNToRecFN.scala 275:77]
  assign _fractOut_T = isNaNOut | io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 278:22]
  assign _fractOut_T_1 = _fractOut_T | common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 278:38]
  assign _fractOut_T_2 = isNaNOut ? 23'h400000 : 23'h0; // @[RoundAnyRawFNToRecFN.scala 279:16]
  assign _fractOut_T_3 = _fractOut_T_1 ? _fractOut_T_2 : common_fractOut; // @[RoundAnyRawFNToRecFN.scala 278:12]
  assign _fractOut_T_5 = pegMaxFiniteMagOut ? 23'h7fffff : 23'h0; // @[Bitwise.scala 72:12]
  assign fractOut = _fractOut_T_3 | _fractOut_T_5; // @[RoundAnyRawFNToRecFN.scala 281:11]
  assign io_out_hi = {signOut,expOut}; // @[Cat.scala 30:58]
  assign io_exceptionFlags_lo = {underflow,inexact}; // @[Cat.scala 30:58]
  assign io_exceptionFlags_hi = {io_invalidExc,1'h0,overflow}; // @[Cat.scala 30:58]
  assign io_out = {io_out_hi,fractOut}; // @[RoundAnyRawFNToRecFN.scala 284:12]
  assign io_exceptionFlags = {io_exceptionFlags_hi,io_exceptionFlags_lo}; // @[RoundAnyRawFNToRecFN.scala 285:23]
  assign RoundAnyRawFNToRecFN_3_covSum = 30'h0;
  assign io_covSum = RoundAnyRawFNToRecFN_3_covSum;
  assign metaAssert = 1'h0;
endmodule
module MulAddRecFNToRaw_preMul_1(
  input  [1:0]   io_op,
  input  [64:0]  io_a,
  input  [64:0]  io_b,
  input  [64:0]  io_c,
  output [52:0]  io_mulAddA,
  output [52:0]  io_mulAddB,
  output [105:0] io_mulAddC,
  output         io_toPostMul_isSigNaNAny,
  output         io_toPostMul_isNaNAOrB,
  output         io_toPostMul_isInfA,
  output         io_toPostMul_isZeroA,
  output         io_toPostMul_isInfB,
  output         io_toPostMul_isZeroB,
  output         io_toPostMul_signProd,
  output         io_toPostMul_isNaNC,
  output         io_toPostMul_isInfC,
  output         io_toPostMul_isZeroC,
  output [12:0]  io_toPostMul_sExpSum,
  output         io_toPostMul_doSubMags,
  output         io_toPostMul_CIsDominant,
  output [5:0]   io_toPostMul_CDom_CAlignDist,
  output [54:0]  io_toPostMul_highAlignedSigC,
  output         io_toPostMul_bit0AlignedSigC,
  output [29:0]  io_covSum,
  output         metaAssert
);
  wire [11:0] rawA_exp; // @[rawFloatFromRecFN.scala 50:21]
  wire  rawA_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  rawA_isSpecial; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawA__isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawA__sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [12:0] rawA__sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire  rawA_out_sig_hi_lo; // @[rawFloatFromRecFN.scala 60:39]
  wire [51:0] rawA_out_sig_lo; // @[rawFloatFromRecFN.scala 60:51]
  wire [53:0] rawA__sig; // @[Cat.scala 30:58]
  wire [11:0] rawB_exp; // @[rawFloatFromRecFN.scala 50:21]
  wire  rawB_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  rawB_isSpecial; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawB__isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawB__sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [12:0] rawB__sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire  rawB_out_sig_hi_lo; // @[rawFloatFromRecFN.scala 60:39]
  wire [51:0] rawB_out_sig_lo; // @[rawFloatFromRecFN.scala 60:51]
  wire [53:0] rawB__sig; // @[Cat.scala 30:58]
  wire [11:0] rawC_exp; // @[rawFloatFromRecFN.scala 50:21]
  wire  rawC_isZero; // @[rawFloatFromRecFN.scala 51:54]
  wire  rawC_isSpecial; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawC__isNaN; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawC__sign; // @[rawFloatFromRecFN.scala 58:25]
  wire [12:0] rawC__sExp; // @[rawFloatFromRecFN.scala 59:27]
  wire  rawC_out_sig_hi_lo; // @[rawFloatFromRecFN.scala 60:39]
  wire [51:0] rawC_out_sig_lo; // @[rawFloatFromRecFN.scala 60:51]
  wire [53:0] rawC__sig; // @[Cat.scala 30:58]
  wire  _signProd_T; // @[MulAddRecFN.scala 98:30]
  wire  signProd; // @[MulAddRecFN.scala 98:42]
  wire [13:0] _sExpAlignedProd_T; // @[MulAddRecFN.scala 101:19]
  wire [13:0] sExpAlignedProd; // @[MulAddRecFN.scala 101:32]
  wire  _doSubMags_T; // @[MulAddRecFN.scala 103:30]
  wire  doSubMags; // @[MulAddRecFN.scala 103:42]
  wire [13:0] _GEN_0; // @[MulAddRecFN.scala 107:42]
  wire [13:0] sNatCAlignDist; // @[MulAddRecFN.scala 107:42]
  wire [12:0] posNatCAlignDist; // @[MulAddRecFN.scala 108:42]
  wire  _isMinCAlign_T; // @[MulAddRecFN.scala 109:35]
  wire  _isMinCAlign_T_1; // @[MulAddRecFN.scala 109:69]
  wire  isMinCAlign; // @[MulAddRecFN.scala 109:50]
  wire  _CIsDominant_T_1; // @[MulAddRecFN.scala 111:60]
  wire  _CIsDominant_T_2; // @[MulAddRecFN.scala 111:39]
  wire  CIsDominant; // @[MulAddRecFN.scala 111:23]
  wire  _CAlignDist_T; // @[MulAddRecFN.scala 115:34]
  wire [7:0] _CAlignDist_T_2; // @[MulAddRecFN.scala 115:16]
  wire [7:0] CAlignDist; // @[MulAddRecFN.scala 113:12]
  wire [53:0] mainAlignedSigC_hi; // @[MulAddRecFN.scala 121:16]
  wire [110:0] mainAlignedSigC_lo; // @[Bitwise.scala 72:12]
  wire [164:0] _mainAlignedSigC_T_3; // @[MulAddRecFN.scala 123:11]
  wire [164:0] mainAlignedSigC; // @[MulAddRecFN.scala 123:17]
  wire  reduced4CExtra_reducedVec_0; // @[primitives.scala 121:54]
  wire  reduced4CExtra_reducedVec_1; // @[primitives.scala 121:54]
  wire  reduced4CExtra_reducedVec_2; // @[primitives.scala 121:54]
  wire  reduced4CExtra_reducedVec_3; // @[primitives.scala 121:54]
  wire  reduced4CExtra_reducedVec_4; // @[primitives.scala 121:54]
  wire  reduced4CExtra_reducedVec_5; // @[primitives.scala 121:54]
  wire  reduced4CExtra_reducedVec_6; // @[primitives.scala 121:54]
  wire  reduced4CExtra_reducedVec_7; // @[primitives.scala 121:54]
  wire  reduced4CExtra_reducedVec_8; // @[primitives.scala 121:54]
  wire  reduced4CExtra_reducedVec_9; // @[primitives.scala 121:54]
  wire  reduced4CExtra_reducedVec_10; // @[primitives.scala 121:54]
  wire  reduced4CExtra_reducedVec_11; // @[primitives.scala 121:54]
  wire  reduced4CExtra_reducedVec_12; // @[primitives.scala 121:54]
  wire  reduced4CExtra_reducedVec_13; // @[primitives.scala 124:57]
  wire [6:0] reduced4CExtra_lo; // @[primitives.scala 125:20]
  wire [13:0] _reduced4CExtra_T_1; // @[primitives.scala 125:20]
  wire [64:0] reduced4CExtra_shift; // @[primitives.scala 77:58]
  wire [7:0] _reduced4CExtra_T_8; // @[Bitwise.scala 103:31]
  wire [7:0] _reduced4CExtra_T_10; // @[Bitwise.scala 103:65]
  wire [7:0] _reduced4CExtra_T_12; // @[Bitwise.scala 103:75]
  wire [7:0] _reduced4CExtra_T_13; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_1; // @[Bitwise.scala 103:31]
  wire [7:0] _reduced4CExtra_T_18; // @[Bitwise.scala 103:31]
  wire [7:0] _reduced4CExtra_T_20; // @[Bitwise.scala 103:65]
  wire [7:0] _reduced4CExtra_T_22; // @[Bitwise.scala 103:75]
  wire [7:0] _reduced4CExtra_T_23; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_2; // @[Bitwise.scala 103:31]
  wire [7:0] _reduced4CExtra_T_28; // @[Bitwise.scala 103:31]
  wire [7:0] _reduced4CExtra_T_30; // @[Bitwise.scala 103:65]
  wire [7:0] _reduced4CExtra_T_32; // @[Bitwise.scala 103:75]
  wire [7:0] reduced4CExtra_hi_1; // @[Bitwise.scala 103:39]
  wire  reduced4CExtra_hi_2; // @[Bitwise.scala 109:18]
  wire  reduced4CExtra_lo_1; // @[Bitwise.scala 109:44]
  wire  reduced4CExtra_hi_4; // @[Bitwise.scala 109:18]
  wire  reduced4CExtra_lo_2; // @[Bitwise.scala 109:44]
  wire  reduced4CExtra_lo_4; // @[Bitwise.scala 109:44]
  wire [12:0] _reduced4CExtra_T_37; // @[Cat.scala 30:58]
  wire [13:0] _GEN_3; // @[MulAddRecFN.scala 125:68]
  wire [13:0] _reduced4CExtra_T_38; // @[MulAddRecFN.scala 125:68]
  wire  reduced4CExtra; // @[MulAddRecFN.scala 133:11]
  wire  _alignedSigC_T_2; // @[MulAddRecFN.scala 137:39]
  wire  _alignedSigC_T_4; // @[MulAddRecFN.scala 137:44]
  wire  _alignedSigC_T_6; // @[MulAddRecFN.scala 138:39]
  wire  _alignedSigC_T_7; // @[MulAddRecFN.scala 138:44]
  wire  alignedSigC_lo; // @[MulAddRecFN.scala 136:16]
  wire [161:0] alignedSigC_hi; // @[Cat.scala 30:58]
  wire [162:0] alignedSigC; // @[Cat.scala 30:58]
  wire  _io_toPostMul_isSigNaNAny_T_2; // @[common.scala 81:46]
  wire  _io_toPostMul_isSigNaNAny_T_5; // @[common.scala 81:46]
  wire  _io_toPostMul_isSigNaNAny_T_6; // @[MulAddRecFN.scala 149:32]
  wire  _io_toPostMul_isSigNaNAny_T_9; // @[common.scala 81:46]
  wire [13:0] _io_toPostMul_sExpSum_T_2; // @[MulAddRecFN.scala 161:53]
  wire [13:0] _io_toPostMul_sExpSum_T_3; // @[MulAddRecFN.scala 161:12]
  wire [29:0] MulAddRecFNToRaw_preMul_1_covSum;
  assign rawA_exp = io_a[63:52]; // @[rawFloatFromRecFN.scala 50:21]
  assign rawA_isZero = rawA_exp[11:9] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign rawA_isSpecial = rawA_exp[11:10] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawA__isNaN = rawA_isSpecial & rawA_exp[9]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawA__sign = io_a[64]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawA__sExp = {1'b0,$signed(rawA_exp)}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawA_out_sig_hi_lo = ~rawA_isZero; // @[rawFloatFromRecFN.scala 60:39]
  assign rawA_out_sig_lo = io_a[51:0]; // @[rawFloatFromRecFN.scala 60:51]
  assign rawA__sig = {1'h0,rawA_out_sig_hi_lo,rawA_out_sig_lo}; // @[Cat.scala 30:58]
  assign rawB_exp = io_b[63:52]; // @[rawFloatFromRecFN.scala 50:21]
  assign rawB_isZero = rawB_exp[11:9] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign rawB_isSpecial = rawB_exp[11:10] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawB__isNaN = rawB_isSpecial & rawB_exp[9]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawB__sign = io_b[64]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawB__sExp = {1'b0,$signed(rawB_exp)}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawB_out_sig_hi_lo = ~rawB_isZero; // @[rawFloatFromRecFN.scala 60:39]
  assign rawB_out_sig_lo = io_b[51:0]; // @[rawFloatFromRecFN.scala 60:51]
  assign rawB__sig = {1'h0,rawB_out_sig_hi_lo,rawB_out_sig_lo}; // @[Cat.scala 30:58]
  assign rawC_exp = io_c[63:52]; // @[rawFloatFromRecFN.scala 50:21]
  assign rawC_isZero = rawC_exp[11:9] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign rawC_isSpecial = rawC_exp[11:10] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  assign rawC__isNaN = rawC_isSpecial & rawC_exp[9]; // @[rawFloatFromRecFN.scala 55:33]
  assign rawC__sign = io_c[64]; // @[rawFloatFromRecFN.scala 58:25]
  assign rawC__sExp = {1'b0,$signed(rawC_exp)}; // @[rawFloatFromRecFN.scala 59:27]
  assign rawC_out_sig_hi_lo = ~rawC_isZero; // @[rawFloatFromRecFN.scala 60:39]
  assign rawC_out_sig_lo = io_c[51:0]; // @[rawFloatFromRecFN.scala 60:51]
  assign rawC__sig = {1'h0,rawC_out_sig_hi_lo,rawC_out_sig_lo}; // @[Cat.scala 30:58]
  assign _signProd_T = rawA__sign ^ rawB__sign; // @[MulAddRecFN.scala 98:30]
  assign signProd = _signProd_T ^ io_op[1]; // @[MulAddRecFN.scala 98:42]
  assign _sExpAlignedProd_T = $signed(rawA__sExp) + $signed(rawB__sExp); // @[MulAddRecFN.scala 101:19]
  assign sExpAlignedProd = $signed(_sExpAlignedProd_T) + -14'sh7c8; // @[MulAddRecFN.scala 101:32]
  assign _doSubMags_T = signProd ^ rawC__sign; // @[MulAddRecFN.scala 103:30]
  assign doSubMags = _doSubMags_T ^ io_op[0]; // @[MulAddRecFN.scala 103:42]
  assign _GEN_0 = {{1{rawC__sExp[12]}},rawC__sExp}; // @[MulAddRecFN.scala 107:42]
  assign sNatCAlignDist = $signed(sExpAlignedProd) - $signed(_GEN_0); // @[MulAddRecFN.scala 107:42]
  assign posNatCAlignDist = sNatCAlignDist[12:0]; // @[MulAddRecFN.scala 108:42]
  assign _isMinCAlign_T = rawA_isZero | rawB_isZero; // @[MulAddRecFN.scala 109:35]
  assign _isMinCAlign_T_1 = $signed(sNatCAlignDist) < 14'sh0; // @[MulAddRecFN.scala 109:69]
  assign isMinCAlign = _isMinCAlign_T | _isMinCAlign_T_1; // @[MulAddRecFN.scala 109:50]
  assign _CIsDominant_T_1 = posNatCAlignDist <= 13'h35; // @[MulAddRecFN.scala 111:60]
  assign _CIsDominant_T_2 = isMinCAlign | _CIsDominant_T_1; // @[MulAddRecFN.scala 111:39]
  assign CIsDominant = rawC_out_sig_hi_lo & _CIsDominant_T_2; // @[MulAddRecFN.scala 111:23]
  assign _CAlignDist_T = posNatCAlignDist < 13'ha1; // @[MulAddRecFN.scala 115:34]
  assign _CAlignDist_T_2 = _CAlignDist_T ? posNatCAlignDist[7:0] : 8'ha1; // @[MulAddRecFN.scala 115:16]
  assign CAlignDist = isMinCAlign ? 8'h0 : _CAlignDist_T_2; // @[MulAddRecFN.scala 113:12]
  assign mainAlignedSigC_hi = doSubMags ? ~rawC__sig : rawC__sig; // @[MulAddRecFN.scala 121:16]
  assign mainAlignedSigC_lo = doSubMags ? 111'h7fffffffffffffffffffffffffff : 111'h0; // @[Bitwise.scala 72:12]
  assign _mainAlignedSigC_T_3 = {mainAlignedSigC_hi,mainAlignedSigC_lo}; // @[MulAddRecFN.scala 123:11]
  assign mainAlignedSigC = $signed(_mainAlignedSigC_T_3) >>> CAlignDist; // @[MulAddRecFN.scala 123:17]
  assign reduced4CExtra_reducedVec_0 = |rawC__sig[3:0]; // @[primitives.scala 121:54]
  assign reduced4CExtra_reducedVec_1 = |rawC__sig[7:4]; // @[primitives.scala 121:54]
  assign reduced4CExtra_reducedVec_2 = |rawC__sig[11:8]; // @[primitives.scala 121:54]
  assign reduced4CExtra_reducedVec_3 = |rawC__sig[15:12]; // @[primitives.scala 121:54]
  assign reduced4CExtra_reducedVec_4 = |rawC__sig[19:16]; // @[primitives.scala 121:54]
  assign reduced4CExtra_reducedVec_5 = |rawC__sig[23:20]; // @[primitives.scala 121:54]
  assign reduced4CExtra_reducedVec_6 = |rawC__sig[27:24]; // @[primitives.scala 121:54]
  assign reduced4CExtra_reducedVec_7 = |rawC__sig[31:28]; // @[primitives.scala 121:54]
  assign reduced4CExtra_reducedVec_8 = |rawC__sig[35:32]; // @[primitives.scala 121:54]
  assign reduced4CExtra_reducedVec_9 = |rawC__sig[39:36]; // @[primitives.scala 121:54]
  assign reduced4CExtra_reducedVec_10 = |rawC__sig[43:40]; // @[primitives.scala 121:54]
  assign reduced4CExtra_reducedVec_11 = |rawC__sig[47:44]; // @[primitives.scala 121:54]
  assign reduced4CExtra_reducedVec_12 = |rawC__sig[51:48]; // @[primitives.scala 121:54]
  assign reduced4CExtra_reducedVec_13 = |rawC__sig[53:52]; // @[primitives.scala 124:57]
  assign reduced4CExtra_lo = {reduced4CExtra_reducedVec_6,reduced4CExtra_reducedVec_5,reduced4CExtra_reducedVec_4,reduced4CExtra_reducedVec_3,reduced4CExtra_reducedVec_2,reduced4CExtra_reducedVec_1,reduced4CExtra_reducedVec_0}; // @[primitives.scala 125:20]
  assign _reduced4CExtra_T_1 = {reduced4CExtra_reducedVec_13,reduced4CExtra_reducedVec_12,reduced4CExtra_reducedVec_11,reduced4CExtra_reducedVec_10,reduced4CExtra_reducedVec_9,reduced4CExtra_reducedVec_8,reduced4CExtra_reducedVec_7,reduced4CExtra_lo}; // @[primitives.scala 125:20]
  assign reduced4CExtra_shift = -65'sh10000000000000000 >>> CAlignDist[7:2]; // @[primitives.scala 77:58]
  assign _reduced4CExtra_T_8 = {{4'd0}, reduced4CExtra_shift[31:28]}; // @[Bitwise.scala 103:31]
  assign _reduced4CExtra_T_10 = {reduced4CExtra_shift[27:24], 4'h0}; // @[Bitwise.scala 103:65]
  assign _reduced4CExtra_T_12 = _reduced4CExtra_T_10 & 8'hf0; // @[Bitwise.scala 103:75]
  assign _reduced4CExtra_T_13 = _reduced4CExtra_T_8 | _reduced4CExtra_T_12; // @[Bitwise.scala 103:39]
  assign _GEN_1 = {{2'd0}, _reduced4CExtra_T_13[7:2]}; // @[Bitwise.scala 103:31]
  assign _reduced4CExtra_T_18 = _GEN_1 & 8'h33; // @[Bitwise.scala 103:31]
  assign _reduced4CExtra_T_20 = {_reduced4CExtra_T_13[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  assign _reduced4CExtra_T_22 = _reduced4CExtra_T_20 & 8'hcc; // @[Bitwise.scala 103:75]
  assign _reduced4CExtra_T_23 = _reduced4CExtra_T_18 | _reduced4CExtra_T_22; // @[Bitwise.scala 103:39]
  assign _GEN_2 = {{1'd0}, _reduced4CExtra_T_23[7:1]}; // @[Bitwise.scala 103:31]
  assign _reduced4CExtra_T_28 = _GEN_2 & 8'h55; // @[Bitwise.scala 103:31]
  assign _reduced4CExtra_T_30 = {_reduced4CExtra_T_23[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  assign _reduced4CExtra_T_32 = _reduced4CExtra_T_30 & 8'haa; // @[Bitwise.scala 103:75]
  assign reduced4CExtra_hi_1 = _reduced4CExtra_T_28 | _reduced4CExtra_T_32; // @[Bitwise.scala 103:39]
  assign reduced4CExtra_hi_2 = reduced4CExtra_shift[32]; // @[Bitwise.scala 109:18]
  assign reduced4CExtra_lo_1 = reduced4CExtra_shift[33]; // @[Bitwise.scala 109:44]
  assign reduced4CExtra_hi_4 = reduced4CExtra_shift[34]; // @[Bitwise.scala 109:18]
  assign reduced4CExtra_lo_2 = reduced4CExtra_shift[35]; // @[Bitwise.scala 109:44]
  assign reduced4CExtra_lo_4 = reduced4CExtra_shift[36]; // @[Bitwise.scala 109:44]
  assign _reduced4CExtra_T_37 = {reduced4CExtra_hi_1,reduced4CExtra_hi_2,reduced4CExtra_lo_1,reduced4CExtra_hi_4,reduced4CExtra_lo_2,reduced4CExtra_lo_4}; // @[Cat.scala 30:58]
  assign _GEN_3 = {{1'd0}, _reduced4CExtra_T_37}; // @[MulAddRecFN.scala 125:68]
  assign _reduced4CExtra_T_38 = _reduced4CExtra_T_1 & _GEN_3; // @[MulAddRecFN.scala 125:68]
  assign reduced4CExtra = |_reduced4CExtra_T_38; // @[MulAddRecFN.scala 133:11]
  assign _alignedSigC_T_2 = &mainAlignedSigC[2:0]; // @[MulAddRecFN.scala 137:39]
  assign _alignedSigC_T_4 = _alignedSigC_T_2 & ~reduced4CExtra; // @[MulAddRecFN.scala 137:44]
  assign _alignedSigC_T_6 = |mainAlignedSigC[2:0]; // @[MulAddRecFN.scala 138:39]
  assign _alignedSigC_T_7 = _alignedSigC_T_6 | reduced4CExtra; // @[MulAddRecFN.scala 138:44]
  assign alignedSigC_lo = doSubMags ? _alignedSigC_T_4 : _alignedSigC_T_7; // @[MulAddRecFN.scala 136:16]
  assign alignedSigC_hi = mainAlignedSigC[164:3]; // @[Cat.scala 30:58]
  assign alignedSigC = {alignedSigC_hi,alignedSigC_lo}; // @[Cat.scala 30:58]
  assign _io_toPostMul_isSigNaNAny_T_2 = rawA__isNaN & ~rawA__sig[51]; // @[common.scala 81:46]
  assign _io_toPostMul_isSigNaNAny_T_5 = rawB__isNaN & ~rawB__sig[51]; // @[common.scala 81:46]
  assign _io_toPostMul_isSigNaNAny_T_6 = _io_toPostMul_isSigNaNAny_T_2 | _io_toPostMul_isSigNaNAny_T_5; // @[MulAddRecFN.scala 149:32]
  assign _io_toPostMul_isSigNaNAny_T_9 = rawC__isNaN & ~rawC__sig[51]; // @[common.scala 81:46]
  assign _io_toPostMul_sExpSum_T_2 = $signed(sExpAlignedProd) - 14'sh35; // @[MulAddRecFN.scala 161:53]
  assign _io_toPostMul_sExpSum_T_3 = CIsDominant ? $signed({{1{rawC__sExp[12]}},rawC__sExp}) : $signed(_io_toPostMul_sExpSum_T_2); // @[MulAddRecFN.scala 161:12]
  assign io_mulAddA = rawA__sig[52:0]; // @[MulAddRecFN.scala 144:16]
  assign io_mulAddB = rawB__sig[52:0]; // @[MulAddRecFN.scala 145:16]
  assign io_mulAddC = alignedSigC[106:1]; // @[MulAddRecFN.scala 146:16]
  assign io_toPostMul_isSigNaNAny = _io_toPostMul_isSigNaNAny_T_6 | _io_toPostMul_isSigNaNAny_T_9; // @[MulAddRecFN.scala 148:30]
  assign io_toPostMul_isNaNAOrB = rawA__isNaN | rawB__isNaN; // @[MulAddRecFN.scala 151:28]
  assign io_toPostMul_isInfA = rawA_isSpecial & ~rawA_exp[9]; // @[MulAddRecFN.scala 152:28]
  assign io_toPostMul_isZeroA = rawA_exp[11:9] == 3'h0; // @[MulAddRecFN.scala 153:28]
  assign io_toPostMul_isInfB = rawB_isSpecial & ~rawB_exp[9]; // @[MulAddRecFN.scala 154:28]
  assign io_toPostMul_isZeroB = rawB_exp[11:9] == 3'h0; // @[MulAddRecFN.scala 155:28]
  assign io_toPostMul_signProd = _signProd_T ^ io_op[1]; // @[MulAddRecFN.scala 156:28]
  assign io_toPostMul_isNaNC = rawC_isSpecial & rawC_exp[9]; // @[MulAddRecFN.scala 157:28]
  assign io_toPostMul_isInfC = rawC_isSpecial & ~rawC_exp[9]; // @[MulAddRecFN.scala 158:28]
  assign io_toPostMul_isZeroC = rawC_exp[11:9] == 3'h0; // @[MulAddRecFN.scala 159:28]
  assign io_toPostMul_sExpSum = _io_toPostMul_sExpSum_T_3[12:0]; // @[MulAddRecFN.scala 160:28]
  assign io_toPostMul_doSubMags = _doSubMags_T ^ io_op[0]; // @[MulAddRecFN.scala 162:28]
  assign io_toPostMul_CIsDominant = rawC_out_sig_hi_lo & _CIsDominant_T_2; // @[MulAddRecFN.scala 163:30]
  assign io_toPostMul_CDom_CAlignDist = CAlignDist[5:0]; // @[MulAddRecFN.scala 164:34]
  assign io_toPostMul_highAlignedSigC = alignedSigC[161:107]; // @[MulAddRecFN.scala 165:34]
  assign io_toPostMul_bit0AlignedSigC = alignedSigC[0]; // @[MulAddRecFN.scala 167:34]
  assign MulAddRecFNToRaw_preMul_1_covSum = 30'h0;
  assign io_covSum = MulAddRecFNToRaw_preMul_1_covSum;
  assign metaAssert = 1'h0;
endmodule
module MulAddRecFNToRaw_postMul_1(
  input          io_fromPreMul_isSigNaNAny,
  input          io_fromPreMul_isNaNAOrB,
  input          io_fromPreMul_isInfA,
  input          io_fromPreMul_isZeroA,
  input          io_fromPreMul_isInfB,
  input          io_fromPreMul_isZeroB,
  input          io_fromPreMul_signProd,
  input          io_fromPreMul_isNaNC,
  input          io_fromPreMul_isInfC,
  input          io_fromPreMul_isZeroC,
  input  [12:0]  io_fromPreMul_sExpSum,
  input          io_fromPreMul_doSubMags,
  input          io_fromPreMul_CIsDominant,
  input  [5:0]   io_fromPreMul_CDom_CAlignDist,
  input  [54:0]  io_fromPreMul_highAlignedSigC,
  input          io_fromPreMul_bit0AlignedSigC,
  input  [106:0] io_mulAddResult,
  input  [2:0]   io_roundingMode,
  output         io_invalidExc,
  output         io_rawOut_isNaN,
  output         io_rawOut_isInf,
  output         io_rawOut_isZero,
  output         io_rawOut_sign,
  output [12:0]  io_rawOut_sExp,
  output [55:0]  io_rawOut_sig,
  output [29:0]  io_covSum,
  output         metaAssert
);
  wire  roundingMode_min; // @[MulAddRecFN.scala 188:45]
  wire  CDom_sign; // @[MulAddRecFN.scala 192:42]
  wire [54:0] _sigSum_T_2; // @[MulAddRecFN.scala 195:47]
  wire [54:0] sigSum_hi_hi; // @[MulAddRecFN.scala 194:16]
  wire [105:0] sigSum_hi_lo; // @[MulAddRecFN.scala 198:28]
  wire [161:0] sigSum; // @[Cat.scala 30:58]
  wire [1:0] _CDom_sExp_T; // @[MulAddRecFN.scala 205:69]
  wire [12:0] _GEN_0; // @[MulAddRecFN.scala 205:43]
  wire [12:0] CDom_sExp; // @[MulAddRecFN.scala 205:43]
  wire [1:0] CDom_absSigSum_hi_lo; // @[MulAddRecFN.scala 211:46]
  wire [104:0] CDom_absSigSum_lo; // @[MulAddRecFN.scala 212:23]
  wire [107:0] _CDom_absSigSum_T_2; // @[Cat.scala 30:58]
  wire [107:0] CDom_absSigSum; // @[MulAddRecFN.scala 207:12]
  wire  _CDom_absSigSumExtra_T_2; // @[MulAddRecFN.scala 217:36]
  wire  _CDom_absSigSumExtra_T_4; // @[MulAddRecFN.scala 218:37]
  wire  CDom_absSigSumExtra; // @[MulAddRecFN.scala 216:12]
  wire [170:0] _GEN_1; // @[MulAddRecFN.scala 221:24]
  wire [170:0] _CDom_mainSig_T; // @[MulAddRecFN.scala 221:24]
  wire [57:0] CDom_mainSig; // @[MulAddRecFN.scala 221:56]
  wire [54:0] _CDom_reduced4SigExtra_T_1; // @[MulAddRecFN.scala 224:53]
  wire  CDom_reduced4SigExtra_reducedVec_0; // @[primitives.scala 121:54]
  wire  CDom_reduced4SigExtra_reducedVec_1; // @[primitives.scala 121:54]
  wire  CDom_reduced4SigExtra_reducedVec_2; // @[primitives.scala 121:54]
  wire  CDom_reduced4SigExtra_reducedVec_3; // @[primitives.scala 121:54]
  wire  CDom_reduced4SigExtra_reducedVec_4; // @[primitives.scala 121:54]
  wire  CDom_reduced4SigExtra_reducedVec_5; // @[primitives.scala 121:54]
  wire  CDom_reduced4SigExtra_reducedVec_6; // @[primitives.scala 121:54]
  wire  CDom_reduced4SigExtra_reducedVec_7; // @[primitives.scala 121:54]
  wire  CDom_reduced4SigExtra_reducedVec_8; // @[primitives.scala 121:54]
  wire  CDom_reduced4SigExtra_reducedVec_9; // @[primitives.scala 121:54]
  wire  CDom_reduced4SigExtra_reducedVec_10; // @[primitives.scala 121:54]
  wire  CDom_reduced4SigExtra_reducedVec_11; // @[primitives.scala 121:54]
  wire  CDom_reduced4SigExtra_reducedVec_12; // @[primitives.scala 121:54]
  wire  CDom_reduced4SigExtra_reducedVec_13; // @[primitives.scala 124:57]
  wire [6:0] CDom_reduced4SigExtra_lo; // @[primitives.scala 125:20]
  wire [13:0] _CDom_reduced4SigExtra_T_2; // @[primitives.scala 125:20]
  wire [16:0] CDom_reduced4SigExtra_shift; // @[primitives.scala 77:58]
  wire [7:0] _CDom_reduced4SigExtra_T_10; // @[Bitwise.scala 103:31]
  wire [7:0] _CDom_reduced4SigExtra_T_12; // @[Bitwise.scala 103:65]
  wire [7:0] _CDom_reduced4SigExtra_T_14; // @[Bitwise.scala 103:75]
  wire [7:0] _CDom_reduced4SigExtra_T_15; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_2; // @[Bitwise.scala 103:31]
  wire [7:0] _CDom_reduced4SigExtra_T_20; // @[Bitwise.scala 103:31]
  wire [7:0] _CDom_reduced4SigExtra_T_22; // @[Bitwise.scala 103:65]
  wire [7:0] _CDom_reduced4SigExtra_T_24; // @[Bitwise.scala 103:75]
  wire [7:0] _CDom_reduced4SigExtra_T_25; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_3; // @[Bitwise.scala 103:31]
  wire [7:0] _CDom_reduced4SigExtra_T_30; // @[Bitwise.scala 103:31]
  wire [7:0] _CDom_reduced4SigExtra_T_32; // @[Bitwise.scala 103:65]
  wire [7:0] _CDom_reduced4SigExtra_T_34; // @[Bitwise.scala 103:75]
  wire [7:0] CDom_reduced4SigExtra_hi_1; // @[Bitwise.scala 103:39]
  wire  CDom_reduced4SigExtra_hi_2; // @[Bitwise.scala 109:18]
  wire  CDom_reduced4SigExtra_lo_1; // @[Bitwise.scala 109:44]
  wire  CDom_reduced4SigExtra_hi_4; // @[Bitwise.scala 109:18]
  wire  CDom_reduced4SigExtra_lo_2; // @[Bitwise.scala 109:44]
  wire  CDom_reduced4SigExtra_lo_4; // @[Bitwise.scala 109:44]
  wire [12:0] _CDom_reduced4SigExtra_T_39; // @[Cat.scala 30:58]
  wire [13:0] _GEN_4; // @[MulAddRecFN.scala 224:72]
  wire [13:0] _CDom_reduced4SigExtra_T_40; // @[MulAddRecFN.scala 224:72]
  wire  CDom_reduced4SigExtra; // @[MulAddRecFN.scala 225:73]
  wire [54:0] CDom_sig_hi; // @[MulAddRecFN.scala 227:25]
  wire  _CDom_sig_T_1; // @[MulAddRecFN.scala 228:32]
  wire  _CDom_sig_T_2; // @[MulAddRecFN.scala 228:36]
  wire  CDom_sig_lo; // @[MulAddRecFN.scala 228:61]
  wire [55:0] CDom_sig; // @[Cat.scala 30:58]
  wire  notCDom_signSigSum; // @[MulAddRecFN.scala 234:36]
  wire [108:0] _GEN_5; // @[MulAddRecFN.scala 238:41]
  wire [108:0] _notCDom_absSigSum_T_4; // @[MulAddRecFN.scala 238:41]
  wire [108:0] notCDom_absSigSum; // @[MulAddRecFN.scala 236:12]
  wire  notCDom_reduced2AbsSigSum_reducedVec_0; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_1; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_2; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_3; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_4; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_5; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_6; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_7; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_8; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_9; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_10; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_11; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_12; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_13; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_14; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_15; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_16; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_17; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_18; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_19; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_20; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_21; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_22; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_23; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_24; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_25; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_26; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_27; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_28; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_29; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_30; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_31; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_32; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_33; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_34; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_35; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_36; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_37; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_38; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_39; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_40; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_41; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_42; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_43; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_44; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_45; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_46; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_47; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_48; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_49; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_50; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_51; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_52; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_53; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_54; // @[primitives.scala 107:57]
  wire [5:0] notCDom_reduced2AbsSigSum_lo_lo_lo; // @[primitives.scala 108:20]
  wire [12:0] notCDom_reduced2AbsSigSum_lo_lo; // @[primitives.scala 108:20]
  wire [6:0] notCDom_reduced2AbsSigSum_lo_hi_lo; // @[primitives.scala 108:20]
  wire [26:0] notCDom_reduced2AbsSigSum_lo; // @[primitives.scala 108:20]
  wire [6:0] notCDom_reduced2AbsSigSum_hi_lo_lo; // @[primitives.scala 108:20]
  wire [13:0] notCDom_reduced2AbsSigSum_hi_lo; // @[primitives.scala 108:20]
  wire [6:0] notCDom_reduced2AbsSigSum_hi_hi_lo; // @[primitives.scala 108:20]
  wire [54:0] notCDom_reduced2AbsSigSum; // @[primitives.scala 108:20]
  wire [5:0] _notCDom_normDistReduced2_T_55; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_56; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_57; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_58; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_59; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_60; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_61; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_62; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_63; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_64; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_65; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_66; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_67; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_68; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_69; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_70; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_71; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_72; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_73; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_74; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_75; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_76; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_77; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_78; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_79; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_80; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_81; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_82; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_83; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_84; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_85; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_86; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_87; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_88; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_89; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_90; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_91; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_92; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_93; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_94; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_95; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_96; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_97; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_98; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_99; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_100; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_101; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_102; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_103; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_104; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_105; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_106; // @[Mux.scala 47:69]
  wire [5:0] _notCDom_normDistReduced2_T_107; // @[Mux.scala 47:69]
  wire [5:0] notCDom_normDistReduced2; // @[Mux.scala 47:69]
  wire [6:0] notCDom_nearNormDist; // @[MulAddRecFN.scala 242:56]
  wire [7:0] _notCDom_sExp_T; // @[MulAddRecFN.scala 243:69]
  wire [12:0] _GEN_6; // @[MulAddRecFN.scala 243:46]
  wire [12:0] notCDom_sExp; // @[MulAddRecFN.scala 243:46]
  wire [235:0] _GEN_7; // @[MulAddRecFN.scala 245:27]
  wire [235:0] _notCDom_mainSig_T; // @[MulAddRecFN.scala 245:27]
  wire [57:0] notCDom_mainSig; // @[MulAddRecFN.scala 245:50]
  wire  notCDom_reduced4SigExtra_reducedVec_0; // @[primitives.scala 104:54]
  wire  notCDom_reduced4SigExtra_reducedVec_1; // @[primitives.scala 104:54]
  wire  notCDom_reduced4SigExtra_reducedVec_2; // @[primitives.scala 104:54]
  wire  notCDom_reduced4SigExtra_reducedVec_3; // @[primitives.scala 104:54]
  wire  notCDom_reduced4SigExtra_reducedVec_4; // @[primitives.scala 104:54]
  wire  notCDom_reduced4SigExtra_reducedVec_5; // @[primitives.scala 104:54]
  wire  notCDom_reduced4SigExtra_reducedVec_6; // @[primitives.scala 104:54]
  wire  notCDom_reduced4SigExtra_reducedVec_7; // @[primitives.scala 104:54]
  wire  notCDom_reduced4SigExtra_reducedVec_8; // @[primitives.scala 104:54]
  wire  notCDom_reduced4SigExtra_reducedVec_9; // @[primitives.scala 104:54]
  wire  notCDom_reduced4SigExtra_reducedVec_10; // @[primitives.scala 104:54]
  wire  notCDom_reduced4SigExtra_reducedVec_11; // @[primitives.scala 104:54]
  wire  notCDom_reduced4SigExtra_reducedVec_12; // @[primitives.scala 104:54]
  wire  notCDom_reduced4SigExtra_reducedVec_13; // @[primitives.scala 107:57]
  wire [6:0] notCDom_reduced4SigExtra_lo; // @[primitives.scala 108:20]
  wire [13:0] _notCDom_reduced4SigExtra_T_2; // @[primitives.scala 108:20]
  wire [32:0] notCDom_reduced4SigExtra_shift; // @[primitives.scala 77:58]
  wire [7:0] _notCDom_reduced4SigExtra_T_10; // @[Bitwise.scala 103:31]
  wire [7:0] _notCDom_reduced4SigExtra_T_12; // @[Bitwise.scala 103:65]
  wire [7:0] _notCDom_reduced4SigExtra_T_14; // @[Bitwise.scala 103:75]
  wire [7:0] _notCDom_reduced4SigExtra_T_15; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_8; // @[Bitwise.scala 103:31]
  wire [7:0] _notCDom_reduced4SigExtra_T_20; // @[Bitwise.scala 103:31]
  wire [7:0] _notCDom_reduced4SigExtra_T_22; // @[Bitwise.scala 103:65]
  wire [7:0] _notCDom_reduced4SigExtra_T_24; // @[Bitwise.scala 103:75]
  wire [7:0] _notCDom_reduced4SigExtra_T_25; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_9; // @[Bitwise.scala 103:31]
  wire [7:0] _notCDom_reduced4SigExtra_T_30; // @[Bitwise.scala 103:31]
  wire [7:0] _notCDom_reduced4SigExtra_T_32; // @[Bitwise.scala 103:65]
  wire [7:0] _notCDom_reduced4SigExtra_T_34; // @[Bitwise.scala 103:75]
  wire [7:0] notCDom_reduced4SigExtra_hi_1; // @[Bitwise.scala 103:39]
  wire  notCDom_reduced4SigExtra_hi_2; // @[Bitwise.scala 109:18]
  wire  notCDom_reduced4SigExtra_lo_1; // @[Bitwise.scala 109:44]
  wire  notCDom_reduced4SigExtra_hi_4; // @[Bitwise.scala 109:18]
  wire  notCDom_reduced4SigExtra_lo_2; // @[Bitwise.scala 109:44]
  wire  notCDom_reduced4SigExtra_lo_4; // @[Bitwise.scala 109:44]
  wire [12:0] _notCDom_reduced4SigExtra_T_39; // @[Cat.scala 30:58]
  wire [13:0] _GEN_10; // @[MulAddRecFN.scala 249:78]
  wire [13:0] _notCDom_reduced4SigExtra_T_40; // @[MulAddRecFN.scala 249:78]
  wire  notCDom_reduced4SigExtra; // @[MulAddRecFN.scala 251:11]
  wire [54:0] notCDom_sig_hi; // @[MulAddRecFN.scala 253:28]
  wire  _notCDom_sig_T_1; // @[MulAddRecFN.scala 254:35]
  wire  notCDom_sig_lo; // @[MulAddRecFN.scala 254:39]
  wire [55:0] notCDom_sig; // @[Cat.scala 30:58]
  wire  notCDom_completeCancellation; // @[MulAddRecFN.scala 257:50]
  wire  _notCDom_sign_T; // @[MulAddRecFN.scala 261:36]
  wire  notCDom_sign; // @[MulAddRecFN.scala 259:12]
  wire  notNaN_isInfProd; // @[MulAddRecFN.scala 266:49]
  wire  notNaN_isInfOut; // @[MulAddRecFN.scala 267:44]
  wire  _notNaN_addZeros_T; // @[MulAddRecFN.scala 269:32]
  wire  notNaN_addZeros; // @[MulAddRecFN.scala 269:58]
  wire  _io_invalidExc_T; // @[MulAddRecFN.scala 274:31]
  wire  _io_invalidExc_T_1; // @[MulAddRecFN.scala 273:35]
  wire  _io_invalidExc_T_2; // @[MulAddRecFN.scala 275:32]
  wire  _io_invalidExc_T_3; // @[MulAddRecFN.scala 274:57]
  wire  _io_invalidExc_T_6; // @[MulAddRecFN.scala 276:36]
  wire  _io_invalidExc_T_7; // @[MulAddRecFN.scala 277:61]
  wire  _io_invalidExc_T_8; // @[MulAddRecFN.scala 278:35]
  wire  _io_rawOut_isZero_T_1; // @[MulAddRecFN.scala 285:42]
  wire  _io_rawOut_sign_T; // @[MulAddRecFN.scala 287:27]
  wire  _io_rawOut_sign_T_1; // @[MulAddRecFN.scala 288:31]
  wire  _io_rawOut_sign_T_2; // @[MulAddRecFN.scala 287:54]
  wire  _io_rawOut_sign_T_4; // @[MulAddRecFN.scala 289:26]
  wire  _io_rawOut_sign_T_5; // @[MulAddRecFN.scala 289:48]
  wire  _io_rawOut_sign_T_6; // @[MulAddRecFN.scala 290:36]
  wire  _io_rawOut_sign_T_7; // @[MulAddRecFN.scala 288:43]
  wire  _io_rawOut_sign_T_8; // @[MulAddRecFN.scala 291:26]
  wire  _io_rawOut_sign_T_9; // @[MulAddRecFN.scala 292:37]
  wire  _io_rawOut_sign_T_10; // @[MulAddRecFN.scala 291:46]
  wire  _io_rawOut_sign_T_11; // @[MulAddRecFN.scala 290:48]
  wire  _io_rawOut_sign_T_14; // @[MulAddRecFN.scala 293:28]
  wire  _io_rawOut_sign_T_15; // @[MulAddRecFN.scala 294:17]
  wire  _io_rawOut_sign_T_16; // @[MulAddRecFN.scala 293:49]
  wire [29:0] MulAddRecFNToRaw_postMul_1_covSum;
  assign roundingMode_min = io_roundingMode == 3'h2; // @[MulAddRecFN.scala 188:45]
  assign CDom_sign = io_fromPreMul_signProd ^ io_fromPreMul_doSubMags; // @[MulAddRecFN.scala 192:42]
  assign _sigSum_T_2 = io_fromPreMul_highAlignedSigC + 55'h1; // @[MulAddRecFN.scala 195:47]
  assign sigSum_hi_hi = io_mulAddResult[106] ? _sigSum_T_2 : io_fromPreMul_highAlignedSigC; // @[MulAddRecFN.scala 194:16]
  assign sigSum_hi_lo = io_mulAddResult[105:0]; // @[MulAddRecFN.scala 198:28]
  assign sigSum = {sigSum_hi_hi,sigSum_hi_lo,io_fromPreMul_bit0AlignedSigC}; // @[Cat.scala 30:58]
  assign _CDom_sExp_T = {1'b0,$signed(io_fromPreMul_doSubMags)}; // @[MulAddRecFN.scala 205:69]
  assign _GEN_0 = {{11{_CDom_sExp_T[1]}},_CDom_sExp_T}; // @[MulAddRecFN.scala 205:43]
  assign CDom_sExp = $signed(io_fromPreMul_sExpSum) - $signed(_GEN_0); // @[MulAddRecFN.scala 205:43]
  assign CDom_absSigSum_hi_lo = io_fromPreMul_highAlignedSigC[54:53]; // @[MulAddRecFN.scala 211:46]
  assign CDom_absSigSum_lo = sigSum[159:55]; // @[MulAddRecFN.scala 212:23]
  assign _CDom_absSigSum_T_2 = {1'h0,CDom_absSigSum_hi_lo,CDom_absSigSum_lo}; // @[Cat.scala 30:58]
  assign CDom_absSigSum = io_fromPreMul_doSubMags ? ~sigSum[161:54] : _CDom_absSigSum_T_2; // @[MulAddRecFN.scala 207:12]
  assign _CDom_absSigSumExtra_T_2 = |(~sigSum[53:1]); // @[MulAddRecFN.scala 217:36]
  assign _CDom_absSigSumExtra_T_4 = |sigSum[54:1]; // @[MulAddRecFN.scala 218:37]
  assign CDom_absSigSumExtra = io_fromPreMul_doSubMags ? _CDom_absSigSumExtra_T_2 : _CDom_absSigSumExtra_T_4; // @[MulAddRecFN.scala 216:12]
  assign _GEN_1 = {{63'd0}, CDom_absSigSum}; // @[MulAddRecFN.scala 221:24]
  assign _CDom_mainSig_T = _GEN_1 << io_fromPreMul_CDom_CAlignDist; // @[MulAddRecFN.scala 221:24]
  assign CDom_mainSig = _CDom_mainSig_T[107:50]; // @[MulAddRecFN.scala 221:56]
  assign _CDom_reduced4SigExtra_T_1 = {CDom_absSigSum[52:0], 2'h0}; // @[MulAddRecFN.scala 224:53]
  assign CDom_reduced4SigExtra_reducedVec_0 = |_CDom_reduced4SigExtra_T_1[3:0]; // @[primitives.scala 121:54]
  assign CDom_reduced4SigExtra_reducedVec_1 = |_CDom_reduced4SigExtra_T_1[7:4]; // @[primitives.scala 121:54]
  assign CDom_reduced4SigExtra_reducedVec_2 = |_CDom_reduced4SigExtra_T_1[11:8]; // @[primitives.scala 121:54]
  assign CDom_reduced4SigExtra_reducedVec_3 = |_CDom_reduced4SigExtra_T_1[15:12]; // @[primitives.scala 121:54]
  assign CDom_reduced4SigExtra_reducedVec_4 = |_CDom_reduced4SigExtra_T_1[19:16]; // @[primitives.scala 121:54]
  assign CDom_reduced4SigExtra_reducedVec_5 = |_CDom_reduced4SigExtra_T_1[23:20]; // @[primitives.scala 121:54]
  assign CDom_reduced4SigExtra_reducedVec_6 = |_CDom_reduced4SigExtra_T_1[27:24]; // @[primitives.scala 121:54]
  assign CDom_reduced4SigExtra_reducedVec_7 = |_CDom_reduced4SigExtra_T_1[31:28]; // @[primitives.scala 121:54]
  assign CDom_reduced4SigExtra_reducedVec_8 = |_CDom_reduced4SigExtra_T_1[35:32]; // @[primitives.scala 121:54]
  assign CDom_reduced4SigExtra_reducedVec_9 = |_CDom_reduced4SigExtra_T_1[39:36]; // @[primitives.scala 121:54]
  assign CDom_reduced4SigExtra_reducedVec_10 = |_CDom_reduced4SigExtra_T_1[43:40]; // @[primitives.scala 121:54]
  assign CDom_reduced4SigExtra_reducedVec_11 = |_CDom_reduced4SigExtra_T_1[47:44]; // @[primitives.scala 121:54]
  assign CDom_reduced4SigExtra_reducedVec_12 = |_CDom_reduced4SigExtra_T_1[51:48]; // @[primitives.scala 121:54]
  assign CDom_reduced4SigExtra_reducedVec_13 = |_CDom_reduced4SigExtra_T_1[54:52]; // @[primitives.scala 124:57]
  assign CDom_reduced4SigExtra_lo = {CDom_reduced4SigExtra_reducedVec_6,CDom_reduced4SigExtra_reducedVec_5,CDom_reduced4SigExtra_reducedVec_4,CDom_reduced4SigExtra_reducedVec_3,CDom_reduced4SigExtra_reducedVec_2,CDom_reduced4SigExtra_reducedVec_1,CDom_reduced4SigExtra_reducedVec_0}; // @[primitives.scala 125:20]
  assign _CDom_reduced4SigExtra_T_2 = {CDom_reduced4SigExtra_reducedVec_13,CDom_reduced4SigExtra_reducedVec_12,CDom_reduced4SigExtra_reducedVec_11,CDom_reduced4SigExtra_reducedVec_10,CDom_reduced4SigExtra_reducedVec_9,CDom_reduced4SigExtra_reducedVec_8,CDom_reduced4SigExtra_reducedVec_7,CDom_reduced4SigExtra_lo}; // @[primitives.scala 125:20]
  assign CDom_reduced4SigExtra_shift = -17'sh10000 >>> ~io_fromPreMul_CDom_CAlignDist[5:2]; // @[primitives.scala 77:58]
  assign _CDom_reduced4SigExtra_T_10 = {{4'd0}, CDom_reduced4SigExtra_shift[8:5]}; // @[Bitwise.scala 103:31]
  assign _CDom_reduced4SigExtra_T_12 = {CDom_reduced4SigExtra_shift[4:1], 4'h0}; // @[Bitwise.scala 103:65]
  assign _CDom_reduced4SigExtra_T_14 = _CDom_reduced4SigExtra_T_12 & 8'hf0; // @[Bitwise.scala 103:75]
  assign _CDom_reduced4SigExtra_T_15 = _CDom_reduced4SigExtra_T_10 | _CDom_reduced4SigExtra_T_14; // @[Bitwise.scala 103:39]
  assign _GEN_2 = {{2'd0}, _CDom_reduced4SigExtra_T_15[7:2]}; // @[Bitwise.scala 103:31]
  assign _CDom_reduced4SigExtra_T_20 = _GEN_2 & 8'h33; // @[Bitwise.scala 103:31]
  assign _CDom_reduced4SigExtra_T_22 = {_CDom_reduced4SigExtra_T_15[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  assign _CDom_reduced4SigExtra_T_24 = _CDom_reduced4SigExtra_T_22 & 8'hcc; // @[Bitwise.scala 103:75]
  assign _CDom_reduced4SigExtra_T_25 = _CDom_reduced4SigExtra_T_20 | _CDom_reduced4SigExtra_T_24; // @[Bitwise.scala 103:39]
  assign _GEN_3 = {{1'd0}, _CDom_reduced4SigExtra_T_25[7:1]}; // @[Bitwise.scala 103:31]
  assign _CDom_reduced4SigExtra_T_30 = _GEN_3 & 8'h55; // @[Bitwise.scala 103:31]
  assign _CDom_reduced4SigExtra_T_32 = {_CDom_reduced4SigExtra_T_25[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  assign _CDom_reduced4SigExtra_T_34 = _CDom_reduced4SigExtra_T_32 & 8'haa; // @[Bitwise.scala 103:75]
  assign CDom_reduced4SigExtra_hi_1 = _CDom_reduced4SigExtra_T_30 | _CDom_reduced4SigExtra_T_34; // @[Bitwise.scala 103:39]
  assign CDom_reduced4SigExtra_hi_2 = CDom_reduced4SigExtra_shift[9]; // @[Bitwise.scala 109:18]
  assign CDom_reduced4SigExtra_lo_1 = CDom_reduced4SigExtra_shift[10]; // @[Bitwise.scala 109:44]
  assign CDom_reduced4SigExtra_hi_4 = CDom_reduced4SigExtra_shift[11]; // @[Bitwise.scala 109:18]
  assign CDom_reduced4SigExtra_lo_2 = CDom_reduced4SigExtra_shift[12]; // @[Bitwise.scala 109:44]
  assign CDom_reduced4SigExtra_lo_4 = CDom_reduced4SigExtra_shift[13]; // @[Bitwise.scala 109:44]
  assign _CDom_reduced4SigExtra_T_39 = {CDom_reduced4SigExtra_hi_1,CDom_reduced4SigExtra_hi_2,CDom_reduced4SigExtra_lo_1,CDom_reduced4SigExtra_hi_4,CDom_reduced4SigExtra_lo_2,CDom_reduced4SigExtra_lo_4}; // @[Cat.scala 30:58]
  assign _GEN_4 = {{1'd0}, _CDom_reduced4SigExtra_T_39}; // @[MulAddRecFN.scala 224:72]
  assign _CDom_reduced4SigExtra_T_40 = _CDom_reduced4SigExtra_T_2 & _GEN_4; // @[MulAddRecFN.scala 224:72]
  assign CDom_reduced4SigExtra = |_CDom_reduced4SigExtra_T_40; // @[MulAddRecFN.scala 225:73]
  assign CDom_sig_hi = CDom_mainSig[57:3]; // @[MulAddRecFN.scala 227:25]
  assign _CDom_sig_T_1 = |CDom_mainSig[2:0]; // @[MulAddRecFN.scala 228:32]
  assign _CDom_sig_T_2 = _CDom_sig_T_1 | CDom_reduced4SigExtra; // @[MulAddRecFN.scala 228:36]
  assign CDom_sig_lo = _CDom_sig_T_2 | CDom_absSigSumExtra; // @[MulAddRecFN.scala 228:61]
  assign CDom_sig = {CDom_sig_hi,CDom_sig_lo}; // @[Cat.scala 30:58]
  assign notCDom_signSigSum = sigSum[109]; // @[MulAddRecFN.scala 234:36]
  assign _GEN_5 = {{108'd0}, io_fromPreMul_doSubMags}; // @[MulAddRecFN.scala 238:41]
  assign _notCDom_absSigSum_T_4 = sigSum[108:0] + _GEN_5; // @[MulAddRecFN.scala 238:41]
  assign notCDom_absSigSum = notCDom_signSigSum ? ~sigSum[108:0] : _notCDom_absSigSum_T_4; // @[MulAddRecFN.scala 236:12]
  assign notCDom_reduced2AbsSigSum_reducedVec_0 = |notCDom_absSigSum[1:0]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_1 = |notCDom_absSigSum[3:2]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_2 = |notCDom_absSigSum[5:4]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_3 = |notCDom_absSigSum[7:6]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_4 = |notCDom_absSigSum[9:8]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_5 = |notCDom_absSigSum[11:10]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_6 = |notCDom_absSigSum[13:12]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_7 = |notCDom_absSigSum[15:14]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_8 = |notCDom_absSigSum[17:16]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_9 = |notCDom_absSigSum[19:18]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_10 = |notCDom_absSigSum[21:20]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_11 = |notCDom_absSigSum[23:22]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_12 = |notCDom_absSigSum[25:24]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_13 = |notCDom_absSigSum[27:26]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_14 = |notCDom_absSigSum[29:28]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_15 = |notCDom_absSigSum[31:30]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_16 = |notCDom_absSigSum[33:32]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_17 = |notCDom_absSigSum[35:34]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_18 = |notCDom_absSigSum[37:36]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_19 = |notCDom_absSigSum[39:38]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_20 = |notCDom_absSigSum[41:40]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_21 = |notCDom_absSigSum[43:42]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_22 = |notCDom_absSigSum[45:44]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_23 = |notCDom_absSigSum[47:46]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_24 = |notCDom_absSigSum[49:48]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_25 = |notCDom_absSigSum[51:50]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_26 = |notCDom_absSigSum[53:52]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_27 = |notCDom_absSigSum[55:54]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_28 = |notCDom_absSigSum[57:56]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_29 = |notCDom_absSigSum[59:58]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_30 = |notCDom_absSigSum[61:60]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_31 = |notCDom_absSigSum[63:62]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_32 = |notCDom_absSigSum[65:64]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_33 = |notCDom_absSigSum[67:66]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_34 = |notCDom_absSigSum[69:68]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_35 = |notCDom_absSigSum[71:70]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_36 = |notCDom_absSigSum[73:72]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_37 = |notCDom_absSigSum[75:74]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_38 = |notCDom_absSigSum[77:76]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_39 = |notCDom_absSigSum[79:78]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_40 = |notCDom_absSigSum[81:80]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_41 = |notCDom_absSigSum[83:82]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_42 = |notCDom_absSigSum[85:84]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_43 = |notCDom_absSigSum[87:86]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_44 = |notCDom_absSigSum[89:88]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_45 = |notCDom_absSigSum[91:90]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_46 = |notCDom_absSigSum[93:92]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_47 = |notCDom_absSigSum[95:94]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_48 = |notCDom_absSigSum[97:96]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_49 = |notCDom_absSigSum[99:98]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_50 = |notCDom_absSigSum[101:100]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_51 = |notCDom_absSigSum[103:102]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_52 = |notCDom_absSigSum[105:104]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_53 = |notCDom_absSigSum[107:106]; // @[primitives.scala 104:54]
  assign notCDom_reduced2AbsSigSum_reducedVec_54 = |notCDom_absSigSum[108]; // @[primitives.scala 107:57]
  assign notCDom_reduced2AbsSigSum_lo_lo_lo = {notCDom_reduced2AbsSigSum_reducedVec_5,notCDom_reduced2AbsSigSum_reducedVec_4,notCDom_reduced2AbsSigSum_reducedVec_3,notCDom_reduced2AbsSigSum_reducedVec_2,notCDom_reduced2AbsSigSum_reducedVec_1,notCDom_reduced2AbsSigSum_reducedVec_0}; // @[primitives.scala 108:20]
  assign notCDom_reduced2AbsSigSum_lo_lo = {notCDom_reduced2AbsSigSum_reducedVec_12,notCDom_reduced2AbsSigSum_reducedVec_11,notCDom_reduced2AbsSigSum_reducedVec_10,notCDom_reduced2AbsSigSum_reducedVec_9,notCDom_reduced2AbsSigSum_reducedVec_8,notCDom_reduced2AbsSigSum_reducedVec_7,notCDom_reduced2AbsSigSum_reducedVec_6,notCDom_reduced2AbsSigSum_lo_lo_lo}; // @[primitives.scala 108:20]
  assign notCDom_reduced2AbsSigSum_lo_hi_lo = {notCDom_reduced2AbsSigSum_reducedVec_19,notCDom_reduced2AbsSigSum_reducedVec_18,notCDom_reduced2AbsSigSum_reducedVec_17,notCDom_reduced2AbsSigSum_reducedVec_16,notCDom_reduced2AbsSigSum_reducedVec_15,notCDom_reduced2AbsSigSum_reducedVec_14,notCDom_reduced2AbsSigSum_reducedVec_13}; // @[primitives.scala 108:20]
  assign notCDom_reduced2AbsSigSum_lo = {notCDom_reduced2AbsSigSum_reducedVec_26,notCDom_reduced2AbsSigSum_reducedVec_25,notCDom_reduced2AbsSigSum_reducedVec_24,notCDom_reduced2AbsSigSum_reducedVec_23,notCDom_reduced2AbsSigSum_reducedVec_22,notCDom_reduced2AbsSigSum_reducedVec_21,notCDom_reduced2AbsSigSum_reducedVec_20,notCDom_reduced2AbsSigSum_lo_hi_lo,notCDom_reduced2AbsSigSum_lo_lo}; // @[primitives.scala 108:20]
  assign notCDom_reduced2AbsSigSum_hi_lo_lo = {notCDom_reduced2AbsSigSum_reducedVec_33,notCDom_reduced2AbsSigSum_reducedVec_32,notCDom_reduced2AbsSigSum_reducedVec_31,notCDom_reduced2AbsSigSum_reducedVec_30,notCDom_reduced2AbsSigSum_reducedVec_29,notCDom_reduced2AbsSigSum_reducedVec_28,notCDom_reduced2AbsSigSum_reducedVec_27}; // @[primitives.scala 108:20]
  assign notCDom_reduced2AbsSigSum_hi_lo = {notCDom_reduced2AbsSigSum_reducedVec_40,notCDom_reduced2AbsSigSum_reducedVec_39,notCDom_reduced2AbsSigSum_reducedVec_38,notCDom_reduced2AbsSigSum_reducedVec_37,notCDom_reduced2AbsSigSum_reducedVec_36,notCDom_reduced2AbsSigSum_reducedVec_35,notCDom_reduced2AbsSigSum_reducedVec_34,notCDom_reduced2AbsSigSum_hi_lo_lo}; // @[primitives.scala 108:20]
  assign notCDom_reduced2AbsSigSum_hi_hi_lo = {notCDom_reduced2AbsSigSum_reducedVec_47,notCDom_reduced2AbsSigSum_reducedVec_46,notCDom_reduced2AbsSigSum_reducedVec_45,notCDom_reduced2AbsSigSum_reducedVec_44,notCDom_reduced2AbsSigSum_reducedVec_43,notCDom_reduced2AbsSigSum_reducedVec_42,notCDom_reduced2AbsSigSum_reducedVec_41}; // @[primitives.scala 108:20]
  assign notCDom_reduced2AbsSigSum = {notCDom_reduced2AbsSigSum_reducedVec_54,notCDom_reduced2AbsSigSum_reducedVec_53,notCDom_reduced2AbsSigSum_reducedVec_52,notCDom_reduced2AbsSigSum_reducedVec_51,notCDom_reduced2AbsSigSum_reducedVec_50,notCDom_reduced2AbsSigSum_reducedVec_49,notCDom_reduced2AbsSigSum_reducedVec_48,notCDom_reduced2AbsSigSum_hi_hi_lo,notCDom_reduced2AbsSigSum_hi_lo,notCDom_reduced2AbsSigSum_lo}; // @[primitives.scala 108:20]
  assign _notCDom_normDistReduced2_T_55 = notCDom_reduced2AbsSigSum[1] ? 6'h35 : 6'h36; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_56 = notCDom_reduced2AbsSigSum[2] ? 6'h34 : _notCDom_normDistReduced2_T_55; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_57 = notCDom_reduced2AbsSigSum[3] ? 6'h33 : _notCDom_normDistReduced2_T_56; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_58 = notCDom_reduced2AbsSigSum[4] ? 6'h32 : _notCDom_normDistReduced2_T_57; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_59 = notCDom_reduced2AbsSigSum[5] ? 6'h31 : _notCDom_normDistReduced2_T_58; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_60 = notCDom_reduced2AbsSigSum[6] ? 6'h30 : _notCDom_normDistReduced2_T_59; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_61 = notCDom_reduced2AbsSigSum[7] ? 6'h2f : _notCDom_normDistReduced2_T_60; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_62 = notCDom_reduced2AbsSigSum[8] ? 6'h2e : _notCDom_normDistReduced2_T_61; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_63 = notCDom_reduced2AbsSigSum[9] ? 6'h2d : _notCDom_normDistReduced2_T_62; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_64 = notCDom_reduced2AbsSigSum[10] ? 6'h2c : _notCDom_normDistReduced2_T_63; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_65 = notCDom_reduced2AbsSigSum[11] ? 6'h2b : _notCDom_normDistReduced2_T_64; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_66 = notCDom_reduced2AbsSigSum[12] ? 6'h2a : _notCDom_normDistReduced2_T_65; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_67 = notCDom_reduced2AbsSigSum[13] ? 6'h29 : _notCDom_normDistReduced2_T_66; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_68 = notCDom_reduced2AbsSigSum[14] ? 6'h28 : _notCDom_normDistReduced2_T_67; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_69 = notCDom_reduced2AbsSigSum[15] ? 6'h27 : _notCDom_normDistReduced2_T_68; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_70 = notCDom_reduced2AbsSigSum[16] ? 6'h26 : _notCDom_normDistReduced2_T_69; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_71 = notCDom_reduced2AbsSigSum[17] ? 6'h25 : _notCDom_normDistReduced2_T_70; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_72 = notCDom_reduced2AbsSigSum[18] ? 6'h24 : _notCDom_normDistReduced2_T_71; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_73 = notCDom_reduced2AbsSigSum[19] ? 6'h23 : _notCDom_normDistReduced2_T_72; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_74 = notCDom_reduced2AbsSigSum[20] ? 6'h22 : _notCDom_normDistReduced2_T_73; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_75 = notCDom_reduced2AbsSigSum[21] ? 6'h21 : _notCDom_normDistReduced2_T_74; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_76 = notCDom_reduced2AbsSigSum[22] ? 6'h20 : _notCDom_normDistReduced2_T_75; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_77 = notCDom_reduced2AbsSigSum[23] ? 6'h1f : _notCDom_normDistReduced2_T_76; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_78 = notCDom_reduced2AbsSigSum[24] ? 6'h1e : _notCDom_normDistReduced2_T_77; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_79 = notCDom_reduced2AbsSigSum[25] ? 6'h1d : _notCDom_normDistReduced2_T_78; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_80 = notCDom_reduced2AbsSigSum[26] ? 6'h1c : _notCDom_normDistReduced2_T_79; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_81 = notCDom_reduced2AbsSigSum[27] ? 6'h1b : _notCDom_normDistReduced2_T_80; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_82 = notCDom_reduced2AbsSigSum[28] ? 6'h1a : _notCDom_normDistReduced2_T_81; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_83 = notCDom_reduced2AbsSigSum[29] ? 6'h19 : _notCDom_normDistReduced2_T_82; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_84 = notCDom_reduced2AbsSigSum[30] ? 6'h18 : _notCDom_normDistReduced2_T_83; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_85 = notCDom_reduced2AbsSigSum[31] ? 6'h17 : _notCDom_normDistReduced2_T_84; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_86 = notCDom_reduced2AbsSigSum[32] ? 6'h16 : _notCDom_normDistReduced2_T_85; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_87 = notCDom_reduced2AbsSigSum[33] ? 6'h15 : _notCDom_normDistReduced2_T_86; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_88 = notCDom_reduced2AbsSigSum[34] ? 6'h14 : _notCDom_normDistReduced2_T_87; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_89 = notCDom_reduced2AbsSigSum[35] ? 6'h13 : _notCDom_normDistReduced2_T_88; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_90 = notCDom_reduced2AbsSigSum[36] ? 6'h12 : _notCDom_normDistReduced2_T_89; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_91 = notCDom_reduced2AbsSigSum[37] ? 6'h11 : _notCDom_normDistReduced2_T_90; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_92 = notCDom_reduced2AbsSigSum[38] ? 6'h10 : _notCDom_normDistReduced2_T_91; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_93 = notCDom_reduced2AbsSigSum[39] ? 6'hf : _notCDom_normDistReduced2_T_92; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_94 = notCDom_reduced2AbsSigSum[40] ? 6'he : _notCDom_normDistReduced2_T_93; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_95 = notCDom_reduced2AbsSigSum[41] ? 6'hd : _notCDom_normDistReduced2_T_94; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_96 = notCDom_reduced2AbsSigSum[42] ? 6'hc : _notCDom_normDistReduced2_T_95; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_97 = notCDom_reduced2AbsSigSum[43] ? 6'hb : _notCDom_normDistReduced2_T_96; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_98 = notCDom_reduced2AbsSigSum[44] ? 6'ha : _notCDom_normDistReduced2_T_97; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_99 = notCDom_reduced2AbsSigSum[45] ? 6'h9 : _notCDom_normDistReduced2_T_98; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_100 = notCDom_reduced2AbsSigSum[46] ? 6'h8 : _notCDom_normDistReduced2_T_99; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_101 = notCDom_reduced2AbsSigSum[47] ? 6'h7 : _notCDom_normDistReduced2_T_100; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_102 = notCDom_reduced2AbsSigSum[48] ? 6'h6 : _notCDom_normDistReduced2_T_101; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_103 = notCDom_reduced2AbsSigSum[49] ? 6'h5 : _notCDom_normDistReduced2_T_102; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_104 = notCDom_reduced2AbsSigSum[50] ? 6'h4 : _notCDom_normDistReduced2_T_103; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_105 = notCDom_reduced2AbsSigSum[51] ? 6'h3 : _notCDom_normDistReduced2_T_104; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_106 = notCDom_reduced2AbsSigSum[52] ? 6'h2 : _notCDom_normDistReduced2_T_105; // @[Mux.scala 47:69]
  assign _notCDom_normDistReduced2_T_107 = notCDom_reduced2AbsSigSum[53] ? 6'h1 : _notCDom_normDistReduced2_T_106; // @[Mux.scala 47:69]
  assign notCDom_normDistReduced2 = notCDom_reduced2AbsSigSum[54] ? 6'h0 : _notCDom_normDistReduced2_T_107; // @[Mux.scala 47:69]
  assign notCDom_nearNormDist = {notCDom_normDistReduced2, 1'h0}; // @[MulAddRecFN.scala 242:56]
  assign _notCDom_sExp_T = {1'b0,$signed(notCDom_nearNormDist)}; // @[MulAddRecFN.scala 243:69]
  assign _GEN_6 = {{5{_notCDom_sExp_T[7]}},_notCDom_sExp_T}; // @[MulAddRecFN.scala 243:46]
  assign notCDom_sExp = $signed(io_fromPreMul_sExpSum) - $signed(_GEN_6); // @[MulAddRecFN.scala 243:46]
  assign _GEN_7 = {{127'd0}, notCDom_absSigSum}; // @[MulAddRecFN.scala 245:27]
  assign _notCDom_mainSig_T = _GEN_7 << notCDom_nearNormDist; // @[MulAddRecFN.scala 245:27]
  assign notCDom_mainSig = _notCDom_mainSig_T[109:52]; // @[MulAddRecFN.scala 245:50]
  assign notCDom_reduced4SigExtra_reducedVec_0 = |notCDom_reduced2AbsSigSum[1:0]; // @[primitives.scala 104:54]
  assign notCDom_reduced4SigExtra_reducedVec_1 = |notCDom_reduced2AbsSigSum[3:2]; // @[primitives.scala 104:54]
  assign notCDom_reduced4SigExtra_reducedVec_2 = |notCDom_reduced2AbsSigSum[5:4]; // @[primitives.scala 104:54]
  assign notCDom_reduced4SigExtra_reducedVec_3 = |notCDom_reduced2AbsSigSum[7:6]; // @[primitives.scala 104:54]
  assign notCDom_reduced4SigExtra_reducedVec_4 = |notCDom_reduced2AbsSigSum[9:8]; // @[primitives.scala 104:54]
  assign notCDom_reduced4SigExtra_reducedVec_5 = |notCDom_reduced2AbsSigSum[11:10]; // @[primitives.scala 104:54]
  assign notCDom_reduced4SigExtra_reducedVec_6 = |notCDom_reduced2AbsSigSum[13:12]; // @[primitives.scala 104:54]
  assign notCDom_reduced4SigExtra_reducedVec_7 = |notCDom_reduced2AbsSigSum[15:14]; // @[primitives.scala 104:54]
  assign notCDom_reduced4SigExtra_reducedVec_8 = |notCDom_reduced2AbsSigSum[17:16]; // @[primitives.scala 104:54]
  assign notCDom_reduced4SigExtra_reducedVec_9 = |notCDom_reduced2AbsSigSum[19:18]; // @[primitives.scala 104:54]
  assign notCDom_reduced4SigExtra_reducedVec_10 = |notCDom_reduced2AbsSigSum[21:20]; // @[primitives.scala 104:54]
  assign notCDom_reduced4SigExtra_reducedVec_11 = |notCDom_reduced2AbsSigSum[23:22]; // @[primitives.scala 104:54]
  assign notCDom_reduced4SigExtra_reducedVec_12 = |notCDom_reduced2AbsSigSum[25:24]; // @[primitives.scala 104:54]
  assign notCDom_reduced4SigExtra_reducedVec_13 = |notCDom_reduced2AbsSigSum[26]; // @[primitives.scala 107:57]
  assign notCDom_reduced4SigExtra_lo = {notCDom_reduced4SigExtra_reducedVec_6,notCDom_reduced4SigExtra_reducedVec_5,notCDom_reduced4SigExtra_reducedVec_4,notCDom_reduced4SigExtra_reducedVec_3,notCDom_reduced4SigExtra_reducedVec_2,notCDom_reduced4SigExtra_reducedVec_1,notCDom_reduced4SigExtra_reducedVec_0}; // @[primitives.scala 108:20]
  assign _notCDom_reduced4SigExtra_T_2 = {notCDom_reduced4SigExtra_reducedVec_13,notCDom_reduced4SigExtra_reducedVec_12,notCDom_reduced4SigExtra_reducedVec_11,notCDom_reduced4SigExtra_reducedVec_10,notCDom_reduced4SigExtra_reducedVec_9,notCDom_reduced4SigExtra_reducedVec_8,notCDom_reduced4SigExtra_reducedVec_7,notCDom_reduced4SigExtra_lo}; // @[primitives.scala 108:20]
  assign notCDom_reduced4SigExtra_shift = -33'sh100000000 >>> ~notCDom_normDistReduced2[5:1]; // @[primitives.scala 77:58]
  assign _notCDom_reduced4SigExtra_T_10 = {{4'd0}, notCDom_reduced4SigExtra_shift[8:5]}; // @[Bitwise.scala 103:31]
  assign _notCDom_reduced4SigExtra_T_12 = {notCDom_reduced4SigExtra_shift[4:1], 4'h0}; // @[Bitwise.scala 103:65]
  assign _notCDom_reduced4SigExtra_T_14 = _notCDom_reduced4SigExtra_T_12 & 8'hf0; // @[Bitwise.scala 103:75]
  assign _notCDom_reduced4SigExtra_T_15 = _notCDom_reduced4SigExtra_T_10 | _notCDom_reduced4SigExtra_T_14; // @[Bitwise.scala 103:39]
  assign _GEN_8 = {{2'd0}, _notCDom_reduced4SigExtra_T_15[7:2]}; // @[Bitwise.scala 103:31]
  assign _notCDom_reduced4SigExtra_T_20 = _GEN_8 & 8'h33; // @[Bitwise.scala 103:31]
  assign _notCDom_reduced4SigExtra_T_22 = {_notCDom_reduced4SigExtra_T_15[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  assign _notCDom_reduced4SigExtra_T_24 = _notCDom_reduced4SigExtra_T_22 & 8'hcc; // @[Bitwise.scala 103:75]
  assign _notCDom_reduced4SigExtra_T_25 = _notCDom_reduced4SigExtra_T_20 | _notCDom_reduced4SigExtra_T_24; // @[Bitwise.scala 103:39]
  assign _GEN_9 = {{1'd0}, _notCDom_reduced4SigExtra_T_25[7:1]}; // @[Bitwise.scala 103:31]
  assign _notCDom_reduced4SigExtra_T_30 = _GEN_9 & 8'h55; // @[Bitwise.scala 103:31]
  assign _notCDom_reduced4SigExtra_T_32 = {_notCDom_reduced4SigExtra_T_25[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  assign _notCDom_reduced4SigExtra_T_34 = _notCDom_reduced4SigExtra_T_32 & 8'haa; // @[Bitwise.scala 103:75]
  assign notCDom_reduced4SigExtra_hi_1 = _notCDom_reduced4SigExtra_T_30 | _notCDom_reduced4SigExtra_T_34; // @[Bitwise.scala 103:39]
  assign notCDom_reduced4SigExtra_hi_2 = notCDom_reduced4SigExtra_shift[9]; // @[Bitwise.scala 109:18]
  assign notCDom_reduced4SigExtra_lo_1 = notCDom_reduced4SigExtra_shift[10]; // @[Bitwise.scala 109:44]
  assign notCDom_reduced4SigExtra_hi_4 = notCDom_reduced4SigExtra_shift[11]; // @[Bitwise.scala 109:18]
  assign notCDom_reduced4SigExtra_lo_2 = notCDom_reduced4SigExtra_shift[12]; // @[Bitwise.scala 109:44]
  assign notCDom_reduced4SigExtra_lo_4 = notCDom_reduced4SigExtra_shift[13]; // @[Bitwise.scala 109:44]
  assign _notCDom_reduced4SigExtra_T_39 = {notCDom_reduced4SigExtra_hi_1,notCDom_reduced4SigExtra_hi_2,notCDom_reduced4SigExtra_lo_1,notCDom_reduced4SigExtra_hi_4,notCDom_reduced4SigExtra_lo_2,notCDom_reduced4SigExtra_lo_4}; // @[Cat.scala 30:58]
  assign _GEN_10 = {{1'd0}, _notCDom_reduced4SigExtra_T_39}; // @[MulAddRecFN.scala 249:78]
  assign _notCDom_reduced4SigExtra_T_40 = _notCDom_reduced4SigExtra_T_2 & _GEN_10; // @[MulAddRecFN.scala 249:78]
  assign notCDom_reduced4SigExtra = |_notCDom_reduced4SigExtra_T_40; // @[MulAddRecFN.scala 251:11]
  assign notCDom_sig_hi = notCDom_mainSig[57:3]; // @[MulAddRecFN.scala 253:28]
  assign _notCDom_sig_T_1 = |notCDom_mainSig[2:0]; // @[MulAddRecFN.scala 254:35]
  assign notCDom_sig_lo = _notCDom_sig_T_1 | notCDom_reduced4SigExtra; // @[MulAddRecFN.scala 254:39]
  assign notCDom_sig = {notCDom_sig_hi,notCDom_sig_lo}; // @[Cat.scala 30:58]
  assign notCDom_completeCancellation = notCDom_sig[55:54] == 2'h0; // @[MulAddRecFN.scala 257:50]
  assign _notCDom_sign_T = io_fromPreMul_signProd ^ notCDom_signSigSum; // @[MulAddRecFN.scala 261:36]
  assign notCDom_sign = notCDom_completeCancellation ? roundingMode_min : _notCDom_sign_T; // @[MulAddRecFN.scala 259:12]
  assign notNaN_isInfProd = io_fromPreMul_isInfA | io_fromPreMul_isInfB; // @[MulAddRecFN.scala 266:49]
  assign notNaN_isInfOut = notNaN_isInfProd | io_fromPreMul_isInfC; // @[MulAddRecFN.scala 267:44]
  assign _notNaN_addZeros_T = io_fromPreMul_isZeroA | io_fromPreMul_isZeroB; // @[MulAddRecFN.scala 269:32]
  assign notNaN_addZeros = _notNaN_addZeros_T & io_fromPreMul_isZeroC; // @[MulAddRecFN.scala 269:58]
  assign _io_invalidExc_T = io_fromPreMul_isInfA & io_fromPreMul_isZeroB; // @[MulAddRecFN.scala 274:31]
  assign _io_invalidExc_T_1 = io_fromPreMul_isSigNaNAny | _io_invalidExc_T; // @[MulAddRecFN.scala 273:35]
  assign _io_invalidExc_T_2 = io_fromPreMul_isZeroA & io_fromPreMul_isInfB; // @[MulAddRecFN.scala 275:32]
  assign _io_invalidExc_T_3 = _io_invalidExc_T_1 | _io_invalidExc_T_2; // @[MulAddRecFN.scala 274:57]
  assign _io_invalidExc_T_6 = ~io_fromPreMul_isNaNAOrB & notNaN_isInfProd; // @[MulAddRecFN.scala 276:36]
  assign _io_invalidExc_T_7 = _io_invalidExc_T_6 & io_fromPreMul_isInfC; // @[MulAddRecFN.scala 277:61]
  assign _io_invalidExc_T_8 = _io_invalidExc_T_7 & io_fromPreMul_doSubMags; // @[MulAddRecFN.scala 278:35]
  assign _io_rawOut_isZero_T_1 = ~io_fromPreMul_CIsDominant & notCDom_completeCancellation; // @[MulAddRecFN.scala 285:42]
  assign _io_rawOut_sign_T = notNaN_isInfProd & io_fromPreMul_signProd; // @[MulAddRecFN.scala 287:27]
  assign _io_rawOut_sign_T_1 = io_fromPreMul_isInfC & CDom_sign; // @[MulAddRecFN.scala 288:31]
  assign _io_rawOut_sign_T_2 = _io_rawOut_sign_T | _io_rawOut_sign_T_1; // @[MulAddRecFN.scala 287:54]
  assign _io_rawOut_sign_T_4 = notNaN_addZeros & ~roundingMode_min; // @[MulAddRecFN.scala 289:26]
  assign _io_rawOut_sign_T_5 = _io_rawOut_sign_T_4 & io_fromPreMul_signProd; // @[MulAddRecFN.scala 289:48]
  assign _io_rawOut_sign_T_6 = _io_rawOut_sign_T_5 & CDom_sign; // @[MulAddRecFN.scala 290:36]
  assign _io_rawOut_sign_T_7 = _io_rawOut_sign_T_2 | _io_rawOut_sign_T_6; // @[MulAddRecFN.scala 288:43]
  assign _io_rawOut_sign_T_8 = notNaN_addZeros & roundingMode_min; // @[MulAddRecFN.scala 291:26]
  assign _io_rawOut_sign_T_9 = io_fromPreMul_signProd | CDom_sign; // @[MulAddRecFN.scala 292:37]
  assign _io_rawOut_sign_T_10 = _io_rawOut_sign_T_8 & _io_rawOut_sign_T_9; // @[MulAddRecFN.scala 291:46]
  assign _io_rawOut_sign_T_11 = _io_rawOut_sign_T_7 | _io_rawOut_sign_T_10; // @[MulAddRecFN.scala 290:48]
  assign _io_rawOut_sign_T_14 = ~notNaN_isInfOut & ~notNaN_addZeros; // @[MulAddRecFN.scala 293:28]
  assign _io_rawOut_sign_T_15 = io_fromPreMul_CIsDominant ? CDom_sign : notCDom_sign; // @[MulAddRecFN.scala 294:17]
  assign _io_rawOut_sign_T_16 = _io_rawOut_sign_T_14 & _io_rawOut_sign_T_15; // @[MulAddRecFN.scala 293:49]
  assign io_invalidExc = _io_invalidExc_T_3 | _io_invalidExc_T_8; // @[MulAddRecFN.scala 272:19]
  assign io_rawOut_isNaN = io_fromPreMul_isNaNAOrB | io_fromPreMul_isNaNC; // @[MulAddRecFN.scala 280:21]
  assign io_rawOut_isInf = notNaN_isInfProd | io_fromPreMul_isInfC; // @[MulAddRecFN.scala 281:21]
  assign io_rawOut_isZero = notNaN_addZeros | _io_rawOut_isZero_T_1; // @[MulAddRecFN.scala 283:22]
  assign io_rawOut_sign = _io_rawOut_sign_T_11 | _io_rawOut_sign_T_16; // @[MulAddRecFN.scala 286:20]
  assign io_rawOut_sExp = io_fromPreMul_CIsDominant ? $signed(CDom_sExp) : $signed(notCDom_sExp); // @[MulAddRecFN.scala 295:20]
  assign io_rawOut_sig = io_fromPreMul_CIsDominant ? CDom_sig : notCDom_sig; // @[MulAddRecFN.scala 296:19]
  assign MulAddRecFNToRaw_postMul_1_covSum = 30'h0;
  assign io_covSum = MulAddRecFNToRaw_postMul_1_covSum;
  assign metaAssert = 1'h0;
endmodule
module DivSqrtRawFN_small(
  input         clock,
  input         reset,
  output        io_inReady,
  input         io_inValid,
  input         io_sqrtOp,
  input         io_a_isNaN,
  input         io_a_isInf,
  input         io_a_isZero,
  input         io_a_sign,
  input  [9:0]  io_a_sExp,
  input  [24:0] io_a_sig,
  input         io_b_isNaN,
  input         io_b_isInf,
  input         io_b_isZero,
  input         io_b_sign,
  input  [9:0]  io_b_sExp,
  input  [24:0] io_b_sig,
  input  [2:0]  io_roundingMode,
  output        io_rawOutValid_div,
  output        io_rawOutValid_sqrt,
  output [2:0]  io_roundingModeOut,
  output        io_invalidExc,
  output        io_infiniteExc,
  output        io_rawOut_isNaN,
  output        io_rawOut_isInf,
  output        io_rawOut_isZero,
  output        io_rawOut_sign,
  output [9:0]  io_rawOut_sExp,
  output [26:0] io_rawOut_sig,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  reg [26:0] cycleNum; // @[DivSqrtRecFN_small.scala 223:33]
  reg [31:0] _RAND_0;
  reg  sqrtOp_Z; // @[DivSqrtRecFN_small.scala 225:29]
  reg [31:0] _RAND_1;
  reg  majorExc_Z; // @[DivSqrtRecFN_small.scala 226:29]
  reg [31:0] _RAND_2;
  reg  isNaN_Z; // @[DivSqrtRecFN_small.scala 228:29]
  reg [31:0] _RAND_3;
  reg  isInf_Z; // @[DivSqrtRecFN_small.scala 229:29]
  reg [31:0] _RAND_4;
  reg  isZero_Z; // @[DivSqrtRecFN_small.scala 230:29]
  reg [31:0] _RAND_5;
  reg  sign_Z; // @[DivSqrtRecFN_small.scala 231:29]
  reg [31:0] _RAND_6;
  reg [9:0] sExp_Z; // @[DivSqrtRecFN_small.scala 232:29]
  reg [31:0] _RAND_7;
  reg [22:0] fractB_Z; // @[DivSqrtRecFN_small.scala 233:29]
  reg [31:0] _RAND_8;
  reg [2:0] roundingMode_Z; // @[DivSqrtRecFN_small.scala 234:29]
  reg [31:0] _RAND_9;
  reg [25:0] rem_Z; // @[DivSqrtRecFN_small.scala 240:29]
  reg [31:0] _RAND_10;
  reg  notZeroRem_Z; // @[DivSqrtRecFN_small.scala 241:29]
  reg [31:0] _RAND_11;
  reg [25:0] sigX_Z; // @[DivSqrtRecFN_small.scala 242:29]
  reg [31:0] _RAND_12;
  wire  _notSigNaNIn_invalidExc_S_div_T; // @[DivSqrtRecFN_small.scala 251:24]
  wire  _notSigNaNIn_invalidExc_S_div_T_1; // @[DivSqrtRecFN_small.scala 251:59]
  wire  notSigNaNIn_invalidExc_S_div; // @[DivSqrtRecFN_small.scala 251:42]
  wire  _notSigNaNIn_invalidExc_S_sqrt_T_2; // @[DivSqrtRecFN_small.scala 253:24]
  wire  notSigNaNIn_invalidExc_S_sqrt; // @[DivSqrtRecFN_small.scala 253:43]
  wire  _majorExc_S_T_2; // @[common.scala 81:46]
  wire  _majorExc_S_T_3; // @[DivSqrtRecFN_small.scala 256:38]
  wire  _majorExc_S_T_9; // @[common.scala 81:46]
  wire  _majorExc_S_T_10; // @[DivSqrtRecFN_small.scala 257:38]
  wire  _majorExc_S_T_11; // @[DivSqrtRecFN_small.scala 257:66]
  wire  _majorExc_S_T_14; // @[DivSqrtRecFN_small.scala 259:33]
  wire  _majorExc_S_T_15; // @[DivSqrtRecFN_small.scala 259:51]
  wire  _majorExc_S_T_16; // @[DivSqrtRecFN_small.scala 258:46]
  wire  _isNaN_S_T; // @[DivSqrtRecFN_small.scala 263:26]
  wire  _isNaN_S_T_1; // @[DivSqrtRecFN_small.scala 264:26]
  wire  _isNaN_S_T_2; // @[DivSqrtRecFN_small.scala 264:42]
  wire  _isInf_S_T; // @[DivSqrtRecFN_small.scala 266:63]
  wire  _isZero_S_T; // @[DivSqrtRecFN_small.scala 267:64]
  wire  _sign_S_T_1; // @[DivSqrtRecFN_small.scala 268:45]
  wire  sign_S; // @[DivSqrtRecFN_small.scala 268:30]
  wire  _specialCaseA_S_T; // @[DivSqrtRecFN_small.scala 270:39]
  wire  specialCaseA_S; // @[DivSqrtRecFN_small.scala 270:55]
  wire  _specialCaseB_S_T; // @[DivSqrtRecFN_small.scala 271:39]
  wire  specialCaseB_S; // @[DivSqrtRecFN_small.scala 271:55]
  wire  normalCase_S_div; // @[DivSqrtRecFN_small.scala 272:45]
  wire  normalCase_S_sqrt; // @[DivSqrtRecFN_small.scala 273:46]
  wire  normalCase_S; // @[DivSqrtRecFN_small.scala 274:27]
  wire  sExpQuot_S_div_hi; // @[DivSqrtRecFN_small.scala 278:28]
  wire [7:0] sExpQuot_S_div_lo; // @[DivSqrtRecFN_small.scala 278:40]
  wire [8:0] _sExpQuot_S_div_T_2; // @[DivSqrtRecFN_small.scala 278:71]
  wire [9:0] _GEN_13; // @[DivSqrtRecFN_small.scala 277:21]
  wire [10:0] sExpQuot_S_div; // @[DivSqrtRecFN_small.scala 277:21]
  wire  _sSatExpQuot_S_div_T; // @[DivSqrtRecFN_small.scala 281:48]
  wire [3:0] sSatExpQuot_S_div_hi; // @[DivSqrtRecFN_small.scala 281:16]
  wire [5:0] sSatExpQuot_S_div_lo; // @[DivSqrtRecFN_small.scala 285:27]
  wire [9:0] sSatExpQuot_S_div; // @[DivSqrtRecFN_small.scala 286:11]
  wire  evenSqrt_S; // @[DivSqrtRecFN_small.scala 288:32]
  wire  oddSqrt_S; // @[DivSqrtRecFN_small.scala 289:32]
  wire  idle; // @[DivSqrtRecFN_small.scala 293:24]
  wire  inReady; // @[DivSqrtRecFN_small.scala 294:24]
  wire  entering; // @[DivSqrtRecFN_small.scala 295:28]
  wire  entering_normalCase; // @[DivSqrtRecFN_small.scala 296:40]
  wire  skipCycle2; // @[DivSqrtRecFN_small.scala 298:34]
  wire  _T_1; // @[DivSqrtRecFN_small.scala 300:18]
  wire  _cycleNum_T_1; // @[DivSqrtRecFN_small.scala 302:26]
  wire [1:0] _cycleNum_T_2; // @[DivSqrtRecFN_small.scala 302:16]
  wire [25:0] _cycleNum_T_4; // @[DivSqrtRecFN_small.scala 305:24]
  wire [26:0] _cycleNum_T_5; // @[DivSqrtRecFN_small.scala 304:20]
  wire [26:0] _cycleNum_T_6; // @[DivSqrtRecFN_small.scala 303:16]
  wire [26:0] _GEN_14; // @[DivSqrtRecFN_small.scala 302:59]
  wire [26:0] _cycleNum_T_7; // @[DivSqrtRecFN_small.scala 302:59]
  wire  _cycleNum_T_10; // @[DivSqrtRecFN_small.scala 310:28]
  wire [25:0] _cycleNum_T_12; // @[DivSqrtRecFN_small.scala 310:16]
  wire [26:0] _GEN_15; // @[DivSqrtRecFN_small.scala 309:15]
  wire [26:0] _cycleNum_T_13; // @[DivSqrtRecFN_small.scala 309:15]
  wire [1:0] _cycleNum_T_14; // @[DivSqrtRecFN_small.scala 311:16]
  wire [26:0] _GEN_16; // @[DivSqrtRecFN_small.scala 310:63]
  wire [26:0] _cycleNum_T_15; // @[DivSqrtRecFN_small.scala 310:63]
  wire [8:0] _sExp_Z_T; // @[DivSqrtRecFN_small.scala 329:29]
  wire [9:0] _sExp_Z_T_1; // @[DivSqrtRecFN_small.scala 329:34]
  wire  _T_3; // @[DivSqrtRecFN_small.scala 334:31]
  wire  _rem_T_1; // @[DivSqrtRecFN_small.scala 341:21]
  wire [25:0] _rem_T_2; // @[DivSqrtRecFN_small.scala 341:47]
  wire [25:0] _rem_T_3; // @[DivSqrtRecFN_small.scala 341:12]
  wire  _rem_T_4; // @[DivSqrtRecFN_small.scala 342:21]
  wire [1:0] rem_hi; // @[DivSqrtRecFN_small.scala 343:56]
  wire [24:0] rem_lo; // @[DivSqrtRecFN_small.scala 344:44]
  wire [26:0] _rem_T_8; // @[Cat.scala 30:58]
  wire [26:0] _rem_T_9; // @[DivSqrtRecFN_small.scala 342:12]
  wire [26:0] _GEN_17; // @[DivSqrtRecFN_small.scala 341:57]
  wire [26:0] _rem_T_10; // @[DivSqrtRecFN_small.scala 341:57]
  wire [26:0] _rem_T_12; // @[DivSqrtRecFN_small.scala 348:29]
  wire [26:0] _rem_T_13; // @[DivSqrtRecFN_small.scala 348:12]
  wire [26:0] rem; // @[DivSqrtRecFN_small.scala 347:11]
  wire [24:0] bitMask; // @[DivSqrtRecFN_small.scala 349:27]
  wire  _trialTerm_T_1; // @[DivSqrtRecFN_small.scala 351:21]
  wire [25:0] _trialTerm_T_2; // @[DivSqrtRecFN_small.scala 351:47]
  wire [25:0] _trialTerm_T_3; // @[DivSqrtRecFN_small.scala 351:12]
  wire  _trialTerm_T_4; // @[DivSqrtRecFN_small.scala 352:21]
  wire [24:0] _trialTerm_T_5; // @[DivSqrtRecFN_small.scala 352:12]
  wire [25:0] _GEN_18; // @[DivSqrtRecFN_small.scala 351:73]
  wire [25:0] _trialTerm_T_6; // @[DivSqrtRecFN_small.scala 351:73]
  wire [25:0] _trialTerm_T_8; // @[DivSqrtRecFN_small.scala 353:12]
  wire [25:0] _trialTerm_T_9; // @[DivSqrtRecFN_small.scala 352:73]
  wire  _trialTerm_T_12; // @[DivSqrtRecFN_small.scala 354:23]
  wire [23:0] _trialTerm_T_13; // @[Cat.scala 30:58]
  wire [24:0] _trialTerm_T_14; // @[DivSqrtRecFN_small.scala 354:56]
  wire [24:0] _trialTerm_T_15; // @[DivSqrtRecFN_small.scala 354:12]
  wire [25:0] _GEN_19; // @[DivSqrtRecFN_small.scala 353:73]
  wire [25:0] _trialTerm_T_16; // @[DivSqrtRecFN_small.scala 353:73]
  wire  _trialTerm_T_18; // @[DivSqrtRecFN_small.scala 355:23]
  wire [26:0] _trialTerm_T_19; // @[DivSqrtRecFN_small.scala 355:44]
  wire [26:0] _GEN_20; // @[DivSqrtRecFN_small.scala 355:48]
  wire [26:0] _trialTerm_T_20; // @[DivSqrtRecFN_small.scala 355:48]
  wire [26:0] _trialTerm_T_21; // @[DivSqrtRecFN_small.scala 355:12]
  wire [26:0] _GEN_21; // @[DivSqrtRecFN_small.scala 354:73]
  wire [26:0] trialTerm; // @[DivSqrtRecFN_small.scala 354:73]
  wire [27:0] _trialRem_T; // @[DivSqrtRecFN_small.scala 356:24]
  wire [27:0] _trialRem_T_1; // @[DivSqrtRecFN_small.scala 356:41]
  wire [27:0] trialRem; // @[DivSqrtRecFN_small.scala 356:29]
  wire  newBit; // @[DivSqrtRecFN_small.scala 357:23]
  wire  _T_5; // @[DivSqrtRecFN_small.scala 359:41]
  wire  _T_7; // @[DivSqrtRecFN_small.scala 359:31]
  wire [27:0] _rem_Z_T; // @[DivSqrtRecFN_small.scala 360:39]
  wire [27:0] _rem_Z_T_1; // @[DivSqrtRecFN_small.scala 360:21]
  wire [27:0] _GEN_10; // @[DivSqrtRecFN_small.scala 359:58]
  wire  _T_9; // @[DivSqrtRecFN_small.scala 362:45]
  wire  _T_10; // @[DivSqrtRecFN_small.scala 362:31]
  wire  _notZeroRem_Z_T; // @[DivSqrtRecFN_small.scala 363:35]
  wire [25:0] _sigX_Z_T_2; // @[DivSqrtRecFN_small.scala 365:47]
  wire [25:0] _sigX_Z_T_3; // @[DivSqrtRecFN_small.scala 365:16]
  wire  _sigX_Z_T_4; // @[DivSqrtRecFN_small.scala 366:25]
  wire [24:0] _sigX_Z_T_5; // @[DivSqrtRecFN_small.scala 366:16]
  wire [25:0] _GEN_22; // @[DivSqrtRecFN_small.scala 365:71]
  wire [25:0] _sigX_Z_T_6; // @[DivSqrtRecFN_small.scala 365:71]
  wire [23:0] _sigX_Z_T_8; // @[DivSqrtRecFN_small.scala 367:47]
  wire [23:0] _sigX_Z_T_9; // @[DivSqrtRecFN_small.scala 367:16]
  wire [25:0] _GEN_23; // @[DivSqrtRecFN_small.scala 366:71]
  wire [25:0] _sigX_Z_T_10; // @[DivSqrtRecFN_small.scala 366:71]
  wire [25:0] _GEN_24; // @[DivSqrtRecFN_small.scala 368:48]
  wire [25:0] _sigX_Z_T_12; // @[DivSqrtRecFN_small.scala 368:48]
  wire [25:0] _sigX_Z_T_13; // @[DivSqrtRecFN_small.scala 368:16]
  wire [25:0] _sigX_Z_T_14; // @[DivSqrtRecFN_small.scala 367:71]
  wire [26:0] _GEN_25; // @[DivSqrtRecFN_small.scala 385:35]
  reg [4:0] DivSqrtRawFN_small_state; // @[Register tracking DivSqrtRawFN_small state]
  reg [31:0] _RAND_13;
  reg  DivSqrtRawFN_small_cov [0:31]; // @[Coverage map for DivSqrtRawFN_small]
  reg [31:0] _RAND_14;
  wire  DivSqrtRawFN_small_cov_read_data; // @[Coverage map for DivSqrtRawFN_small]
  wire [4:0] DivSqrtRawFN_small_cov_read_addr; // @[Coverage map for DivSqrtRawFN_small]
  wire  DivSqrtRawFN_small_cov_write_data; // @[Coverage map for DivSqrtRawFN_small]
  wire [4:0] DivSqrtRawFN_small_cov_write_addr; // @[Coverage map for DivSqrtRawFN_small]
  wire  DivSqrtRawFN_small_cov_write_mask; // @[Coverage map for DivSqrtRawFN_small]
  wire  DivSqrtRawFN_small_cov_write_en; // @[Coverage map for DivSqrtRawFN_small]
  reg [29:0] DivSqrtRawFN_small_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_15;
  wire  mux_cond_0;
  wire  mux_cond_1;
  wire  mux_cond_2;
  wire  mux_cond_3;
  wire  sqrtOp_Z_shl;
  wire [4:0] sqrtOp_Z_pad;
  wire [1:0] mux_cond_0_shl;
  wire [4:0] mux_cond_0_pad;
  wire [2:0] mux_cond_1_shl;
  wire [4:0] mux_cond_1_pad;
  wire [3:0] mux_cond_2_shl;
  wire [4:0] mux_cond_2_pad;
  wire [4:0] mux_cond_3_shl;
  wire [4:0] mux_cond_3_pad;
  wire [4:0] DivSqrtRawFN_small_xor1;
  wire [4:0] DivSqrtRawFN_small_xor6;
  wire [4:0] DivSqrtRawFN_small_xor2;
  wire [4:0] DivSqrtRawFN_small_xor0;
  assign _notSigNaNIn_invalidExc_S_div_T = io_a_isZero & io_b_isZero; // @[DivSqrtRecFN_small.scala 251:24]
  assign _notSigNaNIn_invalidExc_S_div_T_1 = io_a_isInf & io_b_isInf; // @[DivSqrtRecFN_small.scala 251:59]
  assign notSigNaNIn_invalidExc_S_div = _notSigNaNIn_invalidExc_S_div_T | _notSigNaNIn_invalidExc_S_div_T_1; // @[DivSqrtRecFN_small.scala 251:42]
  assign _notSigNaNIn_invalidExc_S_sqrt_T_2 = ~io_a_isNaN & ~io_a_isZero; // @[DivSqrtRecFN_small.scala 253:24]
  assign notSigNaNIn_invalidExc_S_sqrt = _notSigNaNIn_invalidExc_S_sqrt_T_2 & io_a_sign; // @[DivSqrtRecFN_small.scala 253:43]
  assign _majorExc_S_T_2 = io_a_isNaN & ~io_a_sig[22]; // @[common.scala 81:46]
  assign _majorExc_S_T_3 = _majorExc_S_T_2 | notSigNaNIn_invalidExc_S_sqrt; // @[DivSqrtRecFN_small.scala 256:38]
  assign _majorExc_S_T_9 = io_b_isNaN & ~io_b_sig[22]; // @[common.scala 81:46]
  assign _majorExc_S_T_10 = _majorExc_S_T_2 | _majorExc_S_T_9; // @[DivSqrtRecFN_small.scala 257:38]
  assign _majorExc_S_T_11 = _majorExc_S_T_10 | notSigNaNIn_invalidExc_S_div; // @[DivSqrtRecFN_small.scala 257:66]
  assign _majorExc_S_T_14 = ~io_a_isNaN & ~io_a_isInf; // @[DivSqrtRecFN_small.scala 259:33]
  assign _majorExc_S_T_15 = _majorExc_S_T_14 & io_b_isZero; // @[DivSqrtRecFN_small.scala 259:51]
  assign _majorExc_S_T_16 = _majorExc_S_T_11 | _majorExc_S_T_15; // @[DivSqrtRecFN_small.scala 258:46]
  assign _isNaN_S_T = io_a_isNaN | notSigNaNIn_invalidExc_S_sqrt; // @[DivSqrtRecFN_small.scala 263:26]
  assign _isNaN_S_T_1 = io_a_isNaN | io_b_isNaN; // @[DivSqrtRecFN_small.scala 264:26]
  assign _isNaN_S_T_2 = _isNaN_S_T_1 | notSigNaNIn_invalidExc_S_div; // @[DivSqrtRecFN_small.scala 264:42]
  assign _isInf_S_T = io_a_isInf | io_b_isZero; // @[DivSqrtRecFN_small.scala 266:63]
  assign _isZero_S_T = io_a_isZero | io_b_isInf; // @[DivSqrtRecFN_small.scala 267:64]
  assign _sign_S_T_1 = ~io_sqrtOp & io_b_sign; // @[DivSqrtRecFN_small.scala 268:45]
  assign sign_S = io_a_sign ^ _sign_S_T_1; // @[DivSqrtRecFN_small.scala 268:30]
  assign _specialCaseA_S_T = io_a_isNaN | io_a_isInf; // @[DivSqrtRecFN_small.scala 270:39]
  assign specialCaseA_S = _specialCaseA_S_T | io_a_isZero; // @[DivSqrtRecFN_small.scala 270:55]
  assign _specialCaseB_S_T = io_b_isNaN | io_b_isInf; // @[DivSqrtRecFN_small.scala 271:39]
  assign specialCaseB_S = _specialCaseB_S_T | io_b_isZero; // @[DivSqrtRecFN_small.scala 271:55]
  assign normalCase_S_div = ~specialCaseA_S & ~specialCaseB_S; // @[DivSqrtRecFN_small.scala 272:45]
  assign normalCase_S_sqrt = ~specialCaseA_S & ~io_a_sign; // @[DivSqrtRecFN_small.scala 273:46]
  assign normalCase_S = io_sqrtOp ? normalCase_S_sqrt : normalCase_S_div; // @[DivSqrtRecFN_small.scala 274:27]
  assign sExpQuot_S_div_hi = io_b_sExp[8]; // @[DivSqrtRecFN_small.scala 278:28]
  assign sExpQuot_S_div_lo = ~io_b_sExp[7:0]; // @[DivSqrtRecFN_small.scala 278:40]
  assign _sExpQuot_S_div_T_2 = {sExpQuot_S_div_hi,sExpQuot_S_div_lo}; // @[DivSqrtRecFN_small.scala 278:71]
  assign _GEN_13 = {{1{_sExpQuot_S_div_T_2[8]}},_sExpQuot_S_div_T_2}; // @[DivSqrtRecFN_small.scala 277:21]
  assign sExpQuot_S_div = $signed(io_a_sExp) + $signed(_GEN_13); // @[DivSqrtRecFN_small.scala 277:21]
  assign _sSatExpQuot_S_div_T = 11'sh1c0 <= $signed(sExpQuot_S_div); // @[DivSqrtRecFN_small.scala 281:48]
  assign sSatExpQuot_S_div_hi = _sSatExpQuot_S_div_T ? 4'h6 : sExpQuot_S_div[9:6]; // @[DivSqrtRecFN_small.scala 281:16]
  assign sSatExpQuot_S_div_lo = sExpQuot_S_div[5:0]; // @[DivSqrtRecFN_small.scala 285:27]
  assign sSatExpQuot_S_div = {sSatExpQuot_S_div_hi,sSatExpQuot_S_div_lo}; // @[DivSqrtRecFN_small.scala 286:11]
  assign evenSqrt_S = io_sqrtOp & ~io_a_sExp[0]; // @[DivSqrtRecFN_small.scala 288:32]
  assign oddSqrt_S = io_sqrtOp & io_a_sExp[0]; // @[DivSqrtRecFN_small.scala 289:32]
  assign idle = cycleNum[0]; // @[DivSqrtRecFN_small.scala 293:24]
  assign inReady = idle | cycleNum[1]; // @[DivSqrtRecFN_small.scala 294:24]
  assign entering = inReady & io_inValid; // @[DivSqrtRecFN_small.scala 295:28]
  assign entering_normalCase = entering & normalCase_S; // @[DivSqrtRecFN_small.scala 296:40]
  assign skipCycle2 = cycleNum[3] & sigX_Z[25]; // @[DivSqrtRecFN_small.scala 298:34]
  assign _T_1 = ~idle | entering; // @[DivSqrtRecFN_small.scala 300:18]
  assign _cycleNum_T_1 = entering & ~normalCase_S; // @[DivSqrtRecFN_small.scala 302:26]
  assign _cycleNum_T_2 = _cycleNum_T_1 ? 2'h2 : 2'h0; // @[DivSqrtRecFN_small.scala 302:16]
  assign _cycleNum_T_4 = io_a_sExp[0] ? 26'h1000000 : 26'h2000000; // @[DivSqrtRecFN_small.scala 305:24]
  assign _cycleNum_T_5 = io_sqrtOp ? {{1'd0}, _cycleNum_T_4} : 27'h4000000; // @[DivSqrtRecFN_small.scala 304:20]
  assign _cycleNum_T_6 = entering_normalCase ? _cycleNum_T_5 : 27'h0; // @[DivSqrtRecFN_small.scala 303:16]
  assign _GEN_14 = {{25'd0}, _cycleNum_T_2}; // @[DivSqrtRecFN_small.scala 302:59]
  assign _cycleNum_T_7 = _GEN_14 | _cycleNum_T_6; // @[DivSqrtRecFN_small.scala 302:59]
  assign _cycleNum_T_10 = ~entering & ~skipCycle2; // @[DivSqrtRecFN_small.scala 310:28]
  assign _cycleNum_T_12 = _cycleNum_T_10 ? cycleNum[26:1] : 26'h0; // @[DivSqrtRecFN_small.scala 310:16]
  assign _GEN_15 = {{1'd0}, _cycleNum_T_12}; // @[DivSqrtRecFN_small.scala 309:15]
  assign _cycleNum_T_13 = _cycleNum_T_7 | _GEN_15; // @[DivSqrtRecFN_small.scala 309:15]
  assign _cycleNum_T_14 = skipCycle2 ? 2'h2 : 2'h0; // @[DivSqrtRecFN_small.scala 311:16]
  assign _GEN_16 = {{25'd0}, _cycleNum_T_14}; // @[DivSqrtRecFN_small.scala 310:63]
  assign _cycleNum_T_15 = _cycleNum_T_13 | _GEN_16; // @[DivSqrtRecFN_small.scala 310:63]
  assign _sExp_Z_T = io_a_sExp[9:1]; // @[DivSqrtRecFN_small.scala 329:29]
  assign _sExp_Z_T_1 = $signed(_sExp_Z_T) + 9'sh80; // @[DivSqrtRecFN_small.scala 329:34]
  assign _T_3 = entering_normalCase & ~io_sqrtOp; // @[DivSqrtRecFN_small.scala 334:31]
  assign _rem_T_1 = inReady & ~oddSqrt_S; // @[DivSqrtRecFN_small.scala 341:21]
  assign _rem_T_2 = {io_a_sig, 1'h0}; // @[DivSqrtRecFN_small.scala 341:47]
  assign _rem_T_3 = _rem_T_1 ? _rem_T_2 : 26'h0; // @[DivSqrtRecFN_small.scala 341:12]
  assign _rem_T_4 = inReady & oddSqrt_S; // @[DivSqrtRecFN_small.scala 342:21]
  assign rem_hi = io_a_sig[23:22] - 2'h1; // @[DivSqrtRecFN_small.scala 343:56]
  assign rem_lo = {io_a_sig[21:0], 3'h0}; // @[DivSqrtRecFN_small.scala 344:44]
  assign _rem_T_8 = {rem_hi,rem_lo}; // @[Cat.scala 30:58]
  assign _rem_T_9 = _rem_T_4 ? _rem_T_8 : 27'h0; // @[DivSqrtRecFN_small.scala 342:12]
  assign _GEN_17 = {{1'd0}, _rem_T_3}; // @[DivSqrtRecFN_small.scala 341:57]
  assign _rem_T_10 = _GEN_17 | _rem_T_9; // @[DivSqrtRecFN_small.scala 341:57]
  assign _rem_T_12 = {rem_Z, 1'h0}; // @[DivSqrtRecFN_small.scala 348:29]
  assign _rem_T_13 = inReady ? 27'h0 : _rem_T_12; // @[DivSqrtRecFN_small.scala 348:12]
  assign rem = _rem_T_10 | _rem_T_13; // @[DivSqrtRecFN_small.scala 347:11]
  assign bitMask = cycleNum[26:2]; // @[DivSqrtRecFN_small.scala 349:27]
  assign _trialTerm_T_1 = inReady & ~io_sqrtOp; // @[DivSqrtRecFN_small.scala 351:21]
  assign _trialTerm_T_2 = {io_b_sig, 1'h0}; // @[DivSqrtRecFN_small.scala 351:47]
  assign _trialTerm_T_3 = _trialTerm_T_1 ? _trialTerm_T_2 : 26'h0; // @[DivSqrtRecFN_small.scala 351:12]
  assign _trialTerm_T_4 = inReady & evenSqrt_S; // @[DivSqrtRecFN_small.scala 352:21]
  assign _trialTerm_T_5 = _trialTerm_T_4 ? 25'h1000000 : 25'h0; // @[DivSqrtRecFN_small.scala 352:12]
  assign _GEN_18 = {{1'd0}, _trialTerm_T_5}; // @[DivSqrtRecFN_small.scala 351:73]
  assign _trialTerm_T_6 = _trialTerm_T_3 | _GEN_18; // @[DivSqrtRecFN_small.scala 351:73]
  assign _trialTerm_T_8 = _rem_T_4 ? 26'h2800000 : 26'h0; // @[DivSqrtRecFN_small.scala 353:12]
  assign _trialTerm_T_9 = _trialTerm_T_6 | _trialTerm_T_8; // @[DivSqrtRecFN_small.scala 352:73]
  assign _trialTerm_T_12 = ~inReady & ~sqrtOp_Z; // @[DivSqrtRecFN_small.scala 354:23]
  assign _trialTerm_T_13 = {1'h1,fractB_Z}; // @[Cat.scala 30:58]
  assign _trialTerm_T_14 = {_trialTerm_T_13, 1'h0}; // @[DivSqrtRecFN_small.scala 354:56]
  assign _trialTerm_T_15 = _trialTerm_T_12 ? _trialTerm_T_14 : 25'h0; // @[DivSqrtRecFN_small.scala 354:12]
  assign _GEN_19 = {{1'd0}, _trialTerm_T_15}; // @[DivSqrtRecFN_small.scala 353:73]
  assign _trialTerm_T_16 = _trialTerm_T_9 | _GEN_19; // @[DivSqrtRecFN_small.scala 353:73]
  assign _trialTerm_T_18 = ~inReady & sqrtOp_Z; // @[DivSqrtRecFN_small.scala 355:23]
  assign _trialTerm_T_19 = {sigX_Z, 1'h0}; // @[DivSqrtRecFN_small.scala 355:44]
  assign _GEN_20 = {{2'd0}, bitMask}; // @[DivSqrtRecFN_small.scala 355:48]
  assign _trialTerm_T_20 = _trialTerm_T_19 | _GEN_20; // @[DivSqrtRecFN_small.scala 355:48]
  assign _trialTerm_T_21 = _trialTerm_T_18 ? _trialTerm_T_20 : 27'h0; // @[DivSqrtRecFN_small.scala 355:12]
  assign _GEN_21 = {{1'd0}, _trialTerm_T_16}; // @[DivSqrtRecFN_small.scala 354:73]
  assign trialTerm = _GEN_21 | _trialTerm_T_21; // @[DivSqrtRecFN_small.scala 354:73]
  assign _trialRem_T = {1'b0,$signed(rem)}; // @[DivSqrtRecFN_small.scala 356:24]
  assign _trialRem_T_1 = {1'b0,$signed(trialTerm)}; // @[DivSqrtRecFN_small.scala 356:41]
  assign trialRem = $signed(_trialRem_T) - $signed(_trialRem_T_1); // @[DivSqrtRecFN_small.scala 356:29]
  assign newBit = 28'sh0 <= $signed(trialRem); // @[DivSqrtRecFN_small.scala 357:23]
  assign _T_5 = idle | cycleNum[2]; // @[DivSqrtRecFN_small.scala 359:41]
  assign _T_7 = entering_normalCase | ~_T_5; // @[DivSqrtRecFN_small.scala 359:31]
  assign _rem_Z_T = $signed(_trialRem_T) - $signed(_trialRem_T_1); // @[DivSqrtRecFN_small.scala 360:39]
  assign _rem_Z_T_1 = newBit ? _rem_Z_T : {{1'd0}, rem}; // @[DivSqrtRecFN_small.scala 360:21]
  assign _GEN_10 = _T_7 ? _rem_Z_T_1 : {{2'd0}, rem_Z}; // @[DivSqrtRecFN_small.scala 359:58]
  assign _T_9 = ~inReady & newBit; // @[DivSqrtRecFN_small.scala 362:45]
  assign _T_10 = entering_normalCase | _T_9; // @[DivSqrtRecFN_small.scala 362:31]
  assign _notZeroRem_Z_T = $signed(trialRem) != 28'sh0; // @[DivSqrtRecFN_small.scala 363:35]
  assign _sigX_Z_T_2 = {newBit, 25'h0}; // @[DivSqrtRecFN_small.scala 365:47]
  assign _sigX_Z_T_3 = _trialTerm_T_1 ? _sigX_Z_T_2 : 26'h0; // @[DivSqrtRecFN_small.scala 365:16]
  assign _sigX_Z_T_4 = inReady & io_sqrtOp; // @[DivSqrtRecFN_small.scala 366:25]
  assign _sigX_Z_T_5 = _sigX_Z_T_4 ? 25'h1000000 : 25'h0; // @[DivSqrtRecFN_small.scala 366:16]
  assign _GEN_22 = {{1'd0}, _sigX_Z_T_5}; // @[DivSqrtRecFN_small.scala 365:71]
  assign _sigX_Z_T_6 = _sigX_Z_T_3 | _GEN_22; // @[DivSqrtRecFN_small.scala 365:71]
  assign _sigX_Z_T_8 = {newBit, 23'h0}; // @[DivSqrtRecFN_small.scala 367:47]
  assign _sigX_Z_T_9 = _rem_T_4 ? _sigX_Z_T_8 : 24'h0; // @[DivSqrtRecFN_small.scala 367:16]
  assign _GEN_23 = {{2'd0}, _sigX_Z_T_9}; // @[DivSqrtRecFN_small.scala 366:71]
  assign _sigX_Z_T_10 = _sigX_Z_T_6 | _GEN_23; // @[DivSqrtRecFN_small.scala 366:71]
  assign _GEN_24 = {{1'd0}, bitMask}; // @[DivSqrtRecFN_small.scala 368:48]
  assign _sigX_Z_T_12 = sigX_Z | _GEN_24; // @[DivSqrtRecFN_small.scala 368:48]
  assign _sigX_Z_T_13 = inReady ? 26'h0 : _sigX_Z_T_12; // @[DivSqrtRecFN_small.scala 368:16]
  assign _sigX_Z_T_14 = _sigX_Z_T_10 | _sigX_Z_T_13; // @[DivSqrtRecFN_small.scala 367:71]
  assign _GEN_25 = {{26'd0}, notZeroRem_Z}; // @[DivSqrtRecFN_small.scala 385:35]
  assign io_inReady = idle | cycleNum[1]; // @[DivSqrtRecFN_small.scala 314:16]
  assign io_rawOutValid_div = cycleNum[1] & ~sqrtOp_Z; // @[DivSqrtRecFN_small.scala 375:25]
  assign io_rawOutValid_sqrt = cycleNum[1] & sqrtOp_Z; // @[DivSqrtRecFN_small.scala 376:25]
  assign io_roundingModeOut = roundingMode_Z; // @[DivSqrtRecFN_small.scala 377:25]
  assign io_invalidExc = majorExc_Z & isNaN_Z; // @[DivSqrtRecFN_small.scala 378:22]
  assign io_infiniteExc = majorExc_Z & ~isNaN_Z; // @[DivSqrtRecFN_small.scala 379:22]
  assign io_rawOut_isNaN = isNaN_Z; // @[DivSqrtRecFN_small.scala 380:22]
  assign io_rawOut_isInf = isInf_Z; // @[DivSqrtRecFN_small.scala 381:22]
  assign io_rawOut_isZero = isZero_Z; // @[DivSqrtRecFN_small.scala 382:22]
  assign io_rawOut_sign = sign_Z; // @[DivSqrtRecFN_small.scala 383:22]
  assign io_rawOut_sExp = sExp_Z; // @[DivSqrtRecFN_small.scala 384:22]
  assign io_rawOut_sig = _trialTerm_T_19 | _GEN_25; // @[DivSqrtRecFN_small.scala 385:22]
  assign DivSqrtRawFN_small_cov_read_addr = DivSqrtRawFN_small_state;
  assign DivSqrtRawFN_small_cov_read_data = DivSqrtRawFN_small_cov[DivSqrtRawFN_small_cov_read_addr]; // @[Coverage map for DivSqrtRawFN_small]
  assign DivSqrtRawFN_small_cov_write_data = 1'h1;
  assign DivSqrtRawFN_small_cov_write_addr = DivSqrtRawFN_small_state;
  assign DivSqrtRawFN_small_cov_write_mask = 1'h1;
  assign DivSqrtRawFN_small_cov_write_en = 1'h1;
  assign mux_cond_0 = _T_10;
  assign mux_cond_1 = newBit;
  assign mux_cond_2 = skipCycle2;
  assign mux_cond_3 = _cycleNum_T_10;
  assign sqrtOp_Z_shl = sqrtOp_Z;
  assign sqrtOp_Z_pad = {4'h0,sqrtOp_Z_shl};
  assign mux_cond_0_shl = {mux_cond_0, 1'h0};
  assign mux_cond_0_pad = {3'h0,mux_cond_0_shl};
  assign mux_cond_1_shl = {mux_cond_1, 2'h0};
  assign mux_cond_1_pad = {2'h0,mux_cond_1_shl};
  assign mux_cond_2_shl = {mux_cond_2, 3'h0};
  assign mux_cond_2_pad = {1'h0,mux_cond_2_shl};
  assign mux_cond_3_shl = {mux_cond_3, 4'h0};
  assign mux_cond_3_pad = mux_cond_3_shl;
  assign DivSqrtRawFN_small_xor1 = sqrtOp_Z_pad ^ mux_cond_0_pad;
  assign DivSqrtRawFN_small_xor6 = mux_cond_2_pad ^ mux_cond_3_pad;
  assign DivSqrtRawFN_small_xor2 = mux_cond_1_pad ^ DivSqrtRawFN_small_xor6;
  assign DivSqrtRawFN_small_xor0 = DivSqrtRawFN_small_xor1 ^ DivSqrtRawFN_small_xor2;
  assign io_covSum = DivSqrtRawFN_small_covSum;
  assign metaAssert = 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycleNum = _RAND_0[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  sqrtOp_Z = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  majorExc_Z = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  isNaN_Z = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  isInf_Z = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  isZero_Z = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  sign_Z = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  sExp_Z = _RAND_7[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  fractB_Z = _RAND_8[22:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  roundingMode_Z = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  rem_Z = _RAND_10[25:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  notZeroRem_Z = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  sigX_Z = _RAND_12[25:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  DivSqrtRawFN_small_state = _RAND_13[4:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    DivSqrtRawFN_small_cov[initvar] = _RAND_14[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  DivSqrtRawFN_small_covSum = _RAND_15[29:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      cycleNum <= 27'h0;
    end else if (reset) begin
      cycleNum <= 27'h1;
    end else if (_T_1) begin
      cycleNum <= _cycleNum_T_15;
    end
    if (metaReset) begin
      sqrtOp_Z <= 1'h0;
    end else if (entering) begin
      sqrtOp_Z <= io_sqrtOp;
    end
    if (metaReset) begin
      majorExc_Z <= 1'h0;
    end else if (entering) begin
      if (io_sqrtOp) begin
        majorExc_Z <= _majorExc_S_T_3;
      end else begin
        majorExc_Z <= _majorExc_S_T_16;
      end
    end
    if (metaReset) begin
      isNaN_Z <= 1'h0;
    end else if (entering) begin
      if (io_sqrtOp) begin
        isNaN_Z <= _isNaN_S_T;
      end else begin
        isNaN_Z <= _isNaN_S_T_2;
      end
    end
    if (metaReset) begin
      isInf_Z <= 1'h0;
    end else if (entering) begin
      if (io_sqrtOp) begin
        isInf_Z <= io_a_isInf;
      end else begin
        isInf_Z <= _isInf_S_T;
      end
    end
    if (metaReset) begin
      isZero_Z <= 1'h0;
    end else if (entering) begin
      if (io_sqrtOp) begin
        isZero_Z <= io_a_isZero;
      end else begin
        isZero_Z <= _isZero_S_T;
      end
    end
    if (metaReset) begin
      sign_Z <= 1'h0;
    end else if (entering) begin
      sign_Z <= sign_S;
    end
    if (metaReset) begin
      sExp_Z <= 10'h0;
    end else if (entering_normalCase) begin
      if (io_sqrtOp) begin
        sExp_Z <= _sExp_Z_T_1;
      end else begin
        sExp_Z <= sSatExpQuot_S_div;
      end
    end
    if (metaReset) begin
      fractB_Z <= 23'h0;
    end else if (_T_3) begin
      fractB_Z <= io_b_sig[22:0];
    end
    if (metaReset) begin
      roundingMode_Z <= 3'h0;
    end else if (entering_normalCase) begin
      roundingMode_Z <= io_roundingMode;
    end
    if (metaReset) begin
      rem_Z <= 26'h0;
    end else begin
      rem_Z <= _GEN_10[25:0];
    end
    if (metaReset) begin
      notZeroRem_Z <= 1'h0;
    end else if (_T_10) begin
      notZeroRem_Z <= _notZeroRem_Z_T;
    end
    if (metaReset) begin
      sigX_Z <= 26'h0;
    end else if (_T_10) begin
      sigX_Z <= _sigX_Z_T_14;
    end
    DivSqrtRawFN_small_state <= DivSqrtRawFN_small_xor0;
    if (!(DivSqrtRawFN_small_cov_read_data)) begin
      DivSqrtRawFN_small_covSum <= DivSqrtRawFN_small_covSum + 1'h1;
    end
  end
  always @(posedge clock) begin
    if(DivSqrtRawFN_small_cov_write_en & DivSqrtRawFN_small_cov_write_mask) begin
      DivSqrtRawFN_small_cov[DivSqrtRawFN_small_cov_write_addr] <= DivSqrtRawFN_small_cov_write_data; // @[Coverage map for DivSqrtRawFN_small]
    end
  end
endmodule
module RoundAnyRawFNToRecFN_5(
  input         io_invalidExc,
  input         io_infiniteExc,
  input         io_in_isNaN,
  input         io_in_isInf,
  input         io_in_isZero,
  input         io_in_sign,
  input  [9:0]  io_in_sExp,
  input  [26:0] io_in_sig,
  input  [2:0]  io_roundingMode,
  input         io_detectTininess,
  output [32:0] io_out,
  output [4:0]  io_exceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  roundingMode_near_even; // @[RoundAnyRawFNToRecFN.scala 88:53]
  wire  roundingMode_min; // @[RoundAnyRawFNToRecFN.scala 90:53]
  wire  roundingMode_max; // @[RoundAnyRawFNToRecFN.scala 91:53]
  wire  roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 92:53]
  wire  roundingMode_odd; // @[RoundAnyRawFNToRecFN.scala 93:53]
  wire  _roundMagUp_T; // @[RoundAnyRawFNToRecFN.scala 96:27]
  wire  _roundMagUp_T_2; // @[RoundAnyRawFNToRecFN.scala 96:63]
  wire  roundMagUp; // @[RoundAnyRawFNToRecFN.scala 96:42]
  wire  doShiftSigDown1; // @[RoundAnyRawFNToRecFN.scala 118:61]
  wire  roundMask_msb; // @[primitives.scala 57:25]
  wire [7:0] roundMask_lsbs; // @[primitives.scala 58:26]
  wire  roundMask_msb_1; // @[primitives.scala 57:25]
  wire [6:0] roundMask_lsbs_1; // @[primitives.scala 58:26]
  wire  roundMask_msb_2; // @[primitives.scala 57:25]
  wire [5:0] roundMask_lsbs_2; // @[primitives.scala 58:26]
  wire [64:0] roundMask_shift; // @[primitives.scala 77:58]
  wire [15:0] _roundMask_T_7; // @[Bitwise.scala 103:31]
  wire [15:0] _roundMask_T_9; // @[Bitwise.scala 103:65]
  wire [15:0] _roundMask_T_11; // @[Bitwise.scala 103:75]
  wire [15:0] _roundMask_T_12; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_0; // @[Bitwise.scala 103:31]
  wire [15:0] _roundMask_T_17; // @[Bitwise.scala 103:31]
  wire [15:0] _roundMask_T_19; // @[Bitwise.scala 103:65]
  wire [15:0] _roundMask_T_21; // @[Bitwise.scala 103:75]
  wire [15:0] _roundMask_T_22; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_1; // @[Bitwise.scala 103:31]
  wire [15:0] _roundMask_T_27; // @[Bitwise.scala 103:31]
  wire [15:0] _roundMask_T_29; // @[Bitwise.scala 103:65]
  wire [15:0] _roundMask_T_31; // @[Bitwise.scala 103:75]
  wire [15:0] _roundMask_T_32; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_2; // @[Bitwise.scala 103:31]
  wire [15:0] _roundMask_T_37; // @[Bitwise.scala 103:31]
  wire [15:0] _roundMask_T_39; // @[Bitwise.scala 103:65]
  wire [15:0] _roundMask_T_41; // @[Bitwise.scala 103:75]
  wire [15:0] roundMask_hi; // @[Bitwise.scala 103:39]
  wire  roundMask_hi_1; // @[Bitwise.scala 109:18]
  wire  roundMask_lo; // @[Bitwise.scala 109:44]
  wire  roundMask_hi_3; // @[Bitwise.scala 109:18]
  wire  roundMask_lo_1; // @[Bitwise.scala 109:44]
  wire  roundMask_hi_5; // @[Bitwise.scala 109:18]
  wire  roundMask_lo_3; // @[Bitwise.scala 109:44]
  wire [21:0] _roundMask_T_47; // @[Cat.scala 30:58]
  wire [21:0] _roundMask_T_49; // @[primitives.scala 74:21]
  wire [21:0] roundMask_hi_6; // @[primitives.scala 74:17]
  wire [24:0] _roundMask_T_50; // @[Cat.scala 30:58]
  wire  roundMask_hi_7; // @[Bitwise.scala 109:18]
  wire  roundMask_lo_6; // @[Bitwise.scala 109:44]
  wire  roundMask_lo_7; // @[Bitwise.scala 109:44]
  wire [2:0] _roundMask_T_53; // @[Cat.scala 30:58]
  wire [2:0] _roundMask_T_54; // @[primitives.scala 61:24]
  wire [24:0] _roundMask_T_55; // @[primitives.scala 66:24]
  wire [24:0] _roundMask_T_56; // @[primitives.scala 61:24]
  wire [24:0] _GEN_3; // @[RoundAnyRawFNToRecFN.scala 157:23]
  wire [24:0] roundMask_hi_9; // @[RoundAnyRawFNToRecFN.scala 157:23]
  wire [26:0] roundMask; // @[Cat.scala 30:58]
  wire [25:0] shiftedRoundMask_lo; // @[RoundAnyRawFNToRecFN.scala 160:57]
  wire [26:0] shiftedRoundMask; // @[Cat.scala 30:58]
  wire [26:0] roundPosMask; // @[RoundAnyRawFNToRecFN.scala 161:46]
  wire [26:0] _roundPosBit_T; // @[RoundAnyRawFNToRecFN.scala 162:40]
  wire  roundPosBit; // @[RoundAnyRawFNToRecFN.scala 162:56]
  wire [26:0] _anyRoundExtra_T; // @[RoundAnyRawFNToRecFN.scala 163:42]
  wire  anyRoundExtra; // @[RoundAnyRawFNToRecFN.scala 163:62]
  wire  anyRound; // @[RoundAnyRawFNToRecFN.scala 164:36]
  wire  _roundIncr_T; // @[RoundAnyRawFNToRecFN.scala 167:38]
  wire  _roundIncr_T_1; // @[RoundAnyRawFNToRecFN.scala 167:67]
  wire  _roundIncr_T_2; // @[RoundAnyRawFNToRecFN.scala 169:29]
  wire  roundIncr; // @[RoundAnyRawFNToRecFN.scala 168:31]
  wire [26:0] _roundedSig_T; // @[RoundAnyRawFNToRecFN.scala 172:32]
  wire [25:0] _roundedSig_T_2; // @[RoundAnyRawFNToRecFN.scala 172:49]
  wire  _roundedSig_T_3; // @[RoundAnyRawFNToRecFN.scala 173:49]
  wire  _roundedSig_T_5; // @[RoundAnyRawFNToRecFN.scala 173:64]
  wire [25:0] _roundedSig_T_7; // @[RoundAnyRawFNToRecFN.scala 173:25]
  wire [25:0] _roundedSig_T_9; // @[RoundAnyRawFNToRecFN.scala 172:61]
  wire [26:0] _roundedSig_T_11; // @[RoundAnyRawFNToRecFN.scala 178:30]
  wire  _roundedSig_T_13; // @[RoundAnyRawFNToRecFN.scala 179:42]
  wire [25:0] _roundedSig_T_15; // @[RoundAnyRawFNToRecFN.scala 179:24]
  wire [25:0] _GEN_4; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [25:0] _roundedSig_T_16; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [25:0] roundedSig; // @[RoundAnyRawFNToRecFN.scala 171:16]
  wire [2:0] _sRoundedExp_T_1; // @[RoundAnyRawFNToRecFN.scala 183:69]
  wire [9:0] _GEN_5; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [10:0] sRoundedExp; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [8:0] common_expOut; // @[RoundAnyRawFNToRecFN.scala 185:37]
  wire [22:0] common_fractOut; // @[RoundAnyRawFNToRecFN.scala 187:16]
  wire [3:0] _common_overflow_T; // @[RoundAnyRawFNToRecFN.scala 194:30]
  wire  common_overflow; // @[RoundAnyRawFNToRecFN.scala 194:50]
  wire  common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 198:31]
  wire  unboundedRange_roundPosBit; // @[RoundAnyRawFNToRecFN.scala 201:16]
  wire  _unboundedRange_anyRound_T_1; // @[RoundAnyRawFNToRecFN.scala 203:30]
  wire  _unboundedRange_anyRound_T_3; // @[RoundAnyRawFNToRecFN.scala 203:70]
  wire  unboundedRange_anyRound; // @[RoundAnyRawFNToRecFN.scala 203:49]
  wire  _unboundedRange_roundIncr_T_1; // @[RoundAnyRawFNToRecFN.scala 205:67]
  wire  _unboundedRange_roundIncr_T_2; // @[RoundAnyRawFNToRecFN.scala 207:29]
  wire  unboundedRange_roundIncr; // @[RoundAnyRawFNToRecFN.scala 206:46]
  wire  roundCarry; // @[RoundAnyRawFNToRecFN.scala 209:16]
  wire [1:0] _common_underflow_T; // @[RoundAnyRawFNToRecFN.scala 218:48]
  wire  _common_underflow_T_1; // @[RoundAnyRawFNToRecFN.scala 218:62]
  wire  _common_underflow_T_2; // @[RoundAnyRawFNToRecFN.scala 218:32]
  wire  _common_underflow_T_5; // @[RoundAnyRawFNToRecFN.scala 219:30]
  wire  _common_underflow_T_6; // @[RoundAnyRawFNToRecFN.scala 218:74]
  wire  _common_underflow_T_10; // @[RoundAnyRawFNToRecFN.scala 221:39]
  wire  _common_underflow_T_12; // @[RoundAnyRawFNToRecFN.scala 220:77]
  wire  _common_underflow_T_13; // @[RoundAnyRawFNToRecFN.scala 224:38]
  wire  _common_underflow_T_14; // @[RoundAnyRawFNToRecFN.scala 225:45]
  wire  _common_underflow_T_15; // @[RoundAnyRawFNToRecFN.scala 225:60]
  wire  _common_underflow_T_17; // @[RoundAnyRawFNToRecFN.scala 219:76]
  wire  common_underflow; // @[RoundAnyRawFNToRecFN.scala 215:40]
  wire  common_inexact; // @[RoundAnyRawFNToRecFN.scala 228:49]
  wire  isNaNOut; // @[RoundAnyRawFNToRecFN.scala 233:34]
  wire  notNaN_isSpecialInfOut; // @[RoundAnyRawFNToRecFN.scala 234:49]
  wire  _commonCase_T_2; // @[RoundAnyRawFNToRecFN.scala 235:33]
  wire  commonCase; // @[RoundAnyRawFNToRecFN.scala 235:61]
  wire  overflow; // @[RoundAnyRawFNToRecFN.scala 236:32]
  wire  underflow; // @[RoundAnyRawFNToRecFN.scala 237:32]
  wire  _inexact_T; // @[RoundAnyRawFNToRecFN.scala 238:43]
  wire  inexact; // @[RoundAnyRawFNToRecFN.scala 238:28]
  wire  overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 241:60]
  wire  _pegMinNonzeroMagOut_T; // @[RoundAnyRawFNToRecFN.scala 243:20]
  wire  _pegMinNonzeroMagOut_T_1; // @[RoundAnyRawFNToRecFN.scala 243:60]
  wire  pegMinNonzeroMagOut; // @[RoundAnyRawFNToRecFN.scala 243:45]
  wire  pegMaxFiniteMagOut; // @[RoundAnyRawFNToRecFN.scala 244:39]
  wire  _notNaN_isInfOut_T; // @[RoundAnyRawFNToRecFN.scala 246:45]
  wire  notNaN_isInfOut; // @[RoundAnyRawFNToRecFN.scala 246:32]
  wire  signOut; // @[RoundAnyRawFNToRecFN.scala 248:22]
  wire  _expOut_T; // @[RoundAnyRawFNToRecFN.scala 251:32]
  wire [8:0] _expOut_T_1; // @[RoundAnyRawFNToRecFN.scala 251:18]
  wire [8:0] _expOut_T_3; // @[RoundAnyRawFNToRecFN.scala 250:24]
  wire [8:0] _expOut_T_5; // @[RoundAnyRawFNToRecFN.scala 255:18]
  wire [8:0] _expOut_T_7; // @[RoundAnyRawFNToRecFN.scala 254:17]
  wire [8:0] _expOut_T_8; // @[RoundAnyRawFNToRecFN.scala 259:18]
  wire [8:0] _expOut_T_10; // @[RoundAnyRawFNToRecFN.scala 258:17]
  wire [8:0] _expOut_T_11; // @[RoundAnyRawFNToRecFN.scala 263:18]
  wire [8:0] _expOut_T_13; // @[RoundAnyRawFNToRecFN.scala 262:17]
  wire [8:0] _expOut_T_14; // @[RoundAnyRawFNToRecFN.scala 267:16]
  wire [8:0] _expOut_T_15; // @[RoundAnyRawFNToRecFN.scala 266:18]
  wire [8:0] _expOut_T_16; // @[RoundAnyRawFNToRecFN.scala 271:16]
  wire [8:0] _expOut_T_17; // @[RoundAnyRawFNToRecFN.scala 270:15]
  wire [8:0] _expOut_T_18; // @[RoundAnyRawFNToRecFN.scala 275:16]
  wire [8:0] _expOut_T_19; // @[RoundAnyRawFNToRecFN.scala 274:15]
  wire [8:0] _expOut_T_20; // @[RoundAnyRawFNToRecFN.scala 276:16]
  wire [8:0] expOut; // @[RoundAnyRawFNToRecFN.scala 275:77]
  wire  _fractOut_T; // @[RoundAnyRawFNToRecFN.scala 278:22]
  wire  _fractOut_T_1; // @[RoundAnyRawFNToRecFN.scala 278:38]
  wire [22:0] _fractOut_T_2; // @[RoundAnyRawFNToRecFN.scala 279:16]
  wire [22:0] _fractOut_T_3; // @[RoundAnyRawFNToRecFN.scala 278:12]
  wire [22:0] _fractOut_T_5; // @[Bitwise.scala 72:12]
  wire [22:0] fractOut; // @[RoundAnyRawFNToRecFN.scala 281:11]
  wire [9:0] io_out_hi; // @[Cat.scala 30:58]
  wire [1:0] io_exceptionFlags_lo; // @[Cat.scala 30:58]
  wire [2:0] io_exceptionFlags_hi; // @[Cat.scala 30:58]
  wire [29:0] RoundAnyRawFNToRecFN_5_covSum;
  assign roundingMode_near_even = io_roundingMode == 3'h0; // @[RoundAnyRawFNToRecFN.scala 88:53]
  assign roundingMode_min = io_roundingMode == 3'h2; // @[RoundAnyRawFNToRecFN.scala 90:53]
  assign roundingMode_max = io_roundingMode == 3'h3; // @[RoundAnyRawFNToRecFN.scala 91:53]
  assign roundingMode_near_maxMag = io_roundingMode == 3'h4; // @[RoundAnyRawFNToRecFN.scala 92:53]
  assign roundingMode_odd = io_roundingMode == 3'h6; // @[RoundAnyRawFNToRecFN.scala 93:53]
  assign _roundMagUp_T = roundingMode_min & io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:27]
  assign _roundMagUp_T_2 = roundingMode_max & ~io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:63]
  assign roundMagUp = _roundMagUp_T | _roundMagUp_T_2; // @[RoundAnyRawFNToRecFN.scala 96:42]
  assign doShiftSigDown1 = io_in_sig[26]; // @[RoundAnyRawFNToRecFN.scala 118:61]
  assign roundMask_msb = ~io_in_sExp[8]; // @[primitives.scala 57:25]
  assign roundMask_lsbs = ~io_in_sExp[7:0]; // @[primitives.scala 58:26]
  assign roundMask_msb_1 = roundMask_lsbs[7]; // @[primitives.scala 57:25]
  assign roundMask_lsbs_1 = roundMask_lsbs[6:0]; // @[primitives.scala 58:26]
  assign roundMask_msb_2 = roundMask_lsbs_1[6]; // @[primitives.scala 57:25]
  assign roundMask_lsbs_2 = roundMask_lsbs_1[5:0]; // @[primitives.scala 58:26]
  assign roundMask_shift = -65'sh10000000000000000 >>> roundMask_lsbs_2; // @[primitives.scala 77:58]
  assign _roundMask_T_7 = {{8'd0}, roundMask_shift[57:50]}; // @[Bitwise.scala 103:31]
  assign _roundMask_T_9 = {roundMask_shift[49:42], 8'h0}; // @[Bitwise.scala 103:65]
  assign _roundMask_T_11 = _roundMask_T_9 & 16'hff00; // @[Bitwise.scala 103:75]
  assign _roundMask_T_12 = _roundMask_T_7 | _roundMask_T_11; // @[Bitwise.scala 103:39]
  assign _GEN_0 = {{4'd0}, _roundMask_T_12[15:4]}; // @[Bitwise.scala 103:31]
  assign _roundMask_T_17 = _GEN_0 & 16'hf0f; // @[Bitwise.scala 103:31]
  assign _roundMask_T_19 = {_roundMask_T_12[11:0], 4'h0}; // @[Bitwise.scala 103:65]
  assign _roundMask_T_21 = _roundMask_T_19 & 16'hf0f0; // @[Bitwise.scala 103:75]
  assign _roundMask_T_22 = _roundMask_T_17 | _roundMask_T_21; // @[Bitwise.scala 103:39]
  assign _GEN_1 = {{2'd0}, _roundMask_T_22[15:2]}; // @[Bitwise.scala 103:31]
  assign _roundMask_T_27 = _GEN_1 & 16'h3333; // @[Bitwise.scala 103:31]
  assign _roundMask_T_29 = {_roundMask_T_22[13:0], 2'h0}; // @[Bitwise.scala 103:65]
  assign _roundMask_T_31 = _roundMask_T_29 & 16'hcccc; // @[Bitwise.scala 103:75]
  assign _roundMask_T_32 = _roundMask_T_27 | _roundMask_T_31; // @[Bitwise.scala 103:39]
  assign _GEN_2 = {{1'd0}, _roundMask_T_32[15:1]}; // @[Bitwise.scala 103:31]
  assign _roundMask_T_37 = _GEN_2 & 16'h5555; // @[Bitwise.scala 103:31]
  assign _roundMask_T_39 = {_roundMask_T_32[14:0], 1'h0}; // @[Bitwise.scala 103:65]
  assign _roundMask_T_41 = _roundMask_T_39 & 16'haaaa; // @[Bitwise.scala 103:75]
  assign roundMask_hi = _roundMask_T_37 | _roundMask_T_41; // @[Bitwise.scala 103:39]
  assign roundMask_hi_1 = roundMask_shift[58]; // @[Bitwise.scala 109:18]
  assign roundMask_lo = roundMask_shift[59]; // @[Bitwise.scala 109:44]
  assign roundMask_hi_3 = roundMask_shift[60]; // @[Bitwise.scala 109:18]
  assign roundMask_lo_1 = roundMask_shift[61]; // @[Bitwise.scala 109:44]
  assign roundMask_hi_5 = roundMask_shift[62]; // @[Bitwise.scala 109:18]
  assign roundMask_lo_3 = roundMask_shift[63]; // @[Bitwise.scala 109:44]
  assign _roundMask_T_47 = {roundMask_hi,roundMask_hi_1,roundMask_lo,roundMask_hi_3,roundMask_lo_1,roundMask_hi_5,roundMask_lo_3}; // @[Cat.scala 30:58]
  assign _roundMask_T_49 = roundMask_msb_2 ? 22'h0 : ~_roundMask_T_47; // @[primitives.scala 74:21]
  assign roundMask_hi_6 = ~_roundMask_T_49; // @[primitives.scala 74:17]
  assign _roundMask_T_50 = {roundMask_hi_6,3'h7}; // @[Cat.scala 30:58]
  assign roundMask_hi_7 = roundMask_shift[0]; // @[Bitwise.scala 109:18]
  assign roundMask_lo_6 = roundMask_shift[1]; // @[Bitwise.scala 109:44]
  assign roundMask_lo_7 = roundMask_shift[2]; // @[Bitwise.scala 109:44]
  assign _roundMask_T_53 = {roundMask_hi_7,roundMask_lo_6,roundMask_lo_7}; // @[Cat.scala 30:58]
  assign _roundMask_T_54 = roundMask_msb_2 ? _roundMask_T_53 : 3'h0; // @[primitives.scala 61:24]
  assign _roundMask_T_55 = roundMask_msb_1 ? _roundMask_T_50 : {{22'd0}, _roundMask_T_54}; // @[primitives.scala 66:24]
  assign _roundMask_T_56 = roundMask_msb ? _roundMask_T_55 : 25'h0; // @[primitives.scala 61:24]
  assign _GEN_3 = {{24'd0}, doShiftSigDown1}; // @[RoundAnyRawFNToRecFN.scala 157:23]
  assign roundMask_hi_9 = _roundMask_T_56 | _GEN_3; // @[RoundAnyRawFNToRecFN.scala 157:23]
  assign roundMask = {roundMask_hi_9,2'h3}; // @[Cat.scala 30:58]
  assign shiftedRoundMask_lo = roundMask[26:1]; // @[RoundAnyRawFNToRecFN.scala 160:57]
  assign shiftedRoundMask = {1'h0,shiftedRoundMask_lo}; // @[Cat.scala 30:58]
  assign roundPosMask = ~shiftedRoundMask & roundMask; // @[RoundAnyRawFNToRecFN.scala 161:46]
  assign _roundPosBit_T = io_in_sig & roundPosMask; // @[RoundAnyRawFNToRecFN.scala 162:40]
  assign roundPosBit = |_roundPosBit_T; // @[RoundAnyRawFNToRecFN.scala 162:56]
  assign _anyRoundExtra_T = io_in_sig & shiftedRoundMask; // @[RoundAnyRawFNToRecFN.scala 163:42]
  assign anyRoundExtra = |_anyRoundExtra_T; // @[RoundAnyRawFNToRecFN.scala 163:62]
  assign anyRound = roundPosBit | anyRoundExtra; // @[RoundAnyRawFNToRecFN.scala 164:36]
  assign _roundIncr_T = roundingMode_near_even | roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 167:38]
  assign _roundIncr_T_1 = _roundIncr_T & roundPosBit; // @[RoundAnyRawFNToRecFN.scala 167:67]
  assign _roundIncr_T_2 = roundMagUp & anyRound; // @[RoundAnyRawFNToRecFN.scala 169:29]
  assign roundIncr = _roundIncr_T_1 | _roundIncr_T_2; // @[RoundAnyRawFNToRecFN.scala 168:31]
  assign _roundedSig_T = io_in_sig | roundMask; // @[RoundAnyRawFNToRecFN.scala 172:32]
  assign _roundedSig_T_2 = _roundedSig_T[26:2] + 25'h1; // @[RoundAnyRawFNToRecFN.scala 172:49]
  assign _roundedSig_T_3 = roundingMode_near_even & roundPosBit; // @[RoundAnyRawFNToRecFN.scala 173:49]
  assign _roundedSig_T_5 = _roundedSig_T_3 & ~anyRoundExtra; // @[RoundAnyRawFNToRecFN.scala 173:64]
  assign _roundedSig_T_7 = _roundedSig_T_5 ? shiftedRoundMask_lo : 26'h0; // @[RoundAnyRawFNToRecFN.scala 173:25]
  assign _roundedSig_T_9 = _roundedSig_T_2 & ~_roundedSig_T_7; // @[RoundAnyRawFNToRecFN.scala 172:61]
  assign _roundedSig_T_11 = io_in_sig & ~roundMask; // @[RoundAnyRawFNToRecFN.scala 178:30]
  assign _roundedSig_T_13 = roundingMode_odd & anyRound; // @[RoundAnyRawFNToRecFN.scala 179:42]
  assign _roundedSig_T_15 = _roundedSig_T_13 ? roundPosMask[26:1] : 26'h0; // @[RoundAnyRawFNToRecFN.scala 179:24]
  assign _GEN_4 = {{1'd0}, _roundedSig_T_11[26:2]}; // @[RoundAnyRawFNToRecFN.scala 178:47]
  assign _roundedSig_T_16 = _GEN_4 | _roundedSig_T_15; // @[RoundAnyRawFNToRecFN.scala 178:47]
  assign roundedSig = roundIncr ? _roundedSig_T_9 : _roundedSig_T_16; // @[RoundAnyRawFNToRecFN.scala 171:16]
  assign _sRoundedExp_T_1 = {1'b0,$signed(roundedSig[25:24])}; // @[RoundAnyRawFNToRecFN.scala 183:69]
  assign _GEN_5 = {{7{_sRoundedExp_T_1[2]}},_sRoundedExp_T_1}; // @[RoundAnyRawFNToRecFN.scala 183:40]
  assign sRoundedExp = $signed(io_in_sExp) + $signed(_GEN_5); // @[RoundAnyRawFNToRecFN.scala 183:40]
  assign common_expOut = sRoundedExp[8:0]; // @[RoundAnyRawFNToRecFN.scala 185:37]
  assign common_fractOut = doShiftSigDown1 ? roundedSig[23:1] : roundedSig[22:0]; // @[RoundAnyRawFNToRecFN.scala 187:16]
  assign _common_overflow_T = sRoundedExp[10:7]; // @[RoundAnyRawFNToRecFN.scala 194:30]
  assign common_overflow = $signed(_common_overflow_T) >= 4'sh3; // @[RoundAnyRawFNToRecFN.scala 194:50]
  assign common_totalUnderflow = $signed(sRoundedExp) < 11'sh6b; // @[RoundAnyRawFNToRecFN.scala 198:31]
  assign unboundedRange_roundPosBit = doShiftSigDown1 ? io_in_sig[2] : io_in_sig[1]; // @[RoundAnyRawFNToRecFN.scala 201:16]
  assign _unboundedRange_anyRound_T_1 = doShiftSigDown1 & io_in_sig[2]; // @[RoundAnyRawFNToRecFN.scala 203:30]
  assign _unboundedRange_anyRound_T_3 = |io_in_sig[1:0]; // @[RoundAnyRawFNToRecFN.scala 203:70]
  assign unboundedRange_anyRound = _unboundedRange_anyRound_T_1 | _unboundedRange_anyRound_T_3; // @[RoundAnyRawFNToRecFN.scala 203:49]
  assign _unboundedRange_roundIncr_T_1 = _roundIncr_T & unboundedRange_roundPosBit; // @[RoundAnyRawFNToRecFN.scala 205:67]
  assign _unboundedRange_roundIncr_T_2 = roundMagUp & unboundedRange_anyRound; // @[RoundAnyRawFNToRecFN.scala 207:29]
  assign unboundedRange_roundIncr = _unboundedRange_roundIncr_T_1 | _unboundedRange_roundIncr_T_2; // @[RoundAnyRawFNToRecFN.scala 206:46]
  assign roundCarry = doShiftSigDown1 ? roundedSig[25] : roundedSig[24]; // @[RoundAnyRawFNToRecFN.scala 209:16]
  assign _common_underflow_T = io_in_sExp[9:8]; // @[RoundAnyRawFNToRecFN.scala 218:48]
  assign _common_underflow_T_1 = $signed(_common_underflow_T) <= 2'sh0; // @[RoundAnyRawFNToRecFN.scala 218:62]
  assign _common_underflow_T_2 = anyRound & _common_underflow_T_1; // @[RoundAnyRawFNToRecFN.scala 218:32]
  assign _common_underflow_T_5 = doShiftSigDown1 ? roundMask[3] : roundMask[2]; // @[RoundAnyRawFNToRecFN.scala 219:30]
  assign _common_underflow_T_6 = _common_underflow_T_2 & _common_underflow_T_5; // @[RoundAnyRawFNToRecFN.scala 218:74]
  assign _common_underflow_T_10 = doShiftSigDown1 ? roundMask[4] : roundMask[3]; // @[RoundAnyRawFNToRecFN.scala 221:39]
  assign _common_underflow_T_12 = io_detectTininess & ~_common_underflow_T_10; // @[RoundAnyRawFNToRecFN.scala 220:77]
  assign _common_underflow_T_13 = _common_underflow_T_12 & roundCarry; // @[RoundAnyRawFNToRecFN.scala 224:38]
  assign _common_underflow_T_14 = _common_underflow_T_13 & roundPosBit; // @[RoundAnyRawFNToRecFN.scala 225:45]
  assign _common_underflow_T_15 = _common_underflow_T_14 & unboundedRange_roundIncr; // @[RoundAnyRawFNToRecFN.scala 225:60]
  assign _common_underflow_T_17 = _common_underflow_T_6 & ~_common_underflow_T_15; // @[RoundAnyRawFNToRecFN.scala 219:76]
  assign common_underflow = common_totalUnderflow | _common_underflow_T_17; // @[RoundAnyRawFNToRecFN.scala 215:40]
  assign common_inexact = common_totalUnderflow | anyRound; // @[RoundAnyRawFNToRecFN.scala 228:49]
  assign isNaNOut = io_invalidExc | io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 233:34]
  assign notNaN_isSpecialInfOut = io_infiniteExc | io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 234:49]
  assign _commonCase_T_2 = ~isNaNOut & ~notNaN_isSpecialInfOut; // @[RoundAnyRawFNToRecFN.scala 235:33]
  assign commonCase = _commonCase_T_2 & ~io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 235:61]
  assign overflow = commonCase & common_overflow; // @[RoundAnyRawFNToRecFN.scala 236:32]
  assign underflow = commonCase & common_underflow; // @[RoundAnyRawFNToRecFN.scala 237:32]
  assign _inexact_T = commonCase & common_inexact; // @[RoundAnyRawFNToRecFN.scala 238:43]
  assign inexact = overflow | _inexact_T; // @[RoundAnyRawFNToRecFN.scala 238:28]
  assign overflow_roundMagUp = _roundIncr_T | roundMagUp; // @[RoundAnyRawFNToRecFN.scala 241:60]
  assign _pegMinNonzeroMagOut_T = commonCase & common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 243:20]
  assign _pegMinNonzeroMagOut_T_1 = roundMagUp | roundingMode_odd; // @[RoundAnyRawFNToRecFN.scala 243:60]
  assign pegMinNonzeroMagOut = _pegMinNonzeroMagOut_T & _pegMinNonzeroMagOut_T_1; // @[RoundAnyRawFNToRecFN.scala 243:45]
  assign pegMaxFiniteMagOut = overflow & ~overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 244:39]
  assign _notNaN_isInfOut_T = overflow & overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 246:45]
  assign notNaN_isInfOut = notNaN_isSpecialInfOut | _notNaN_isInfOut_T; // @[RoundAnyRawFNToRecFN.scala 246:32]
  assign signOut = isNaNOut ? 1'h0 : io_in_sign; // @[RoundAnyRawFNToRecFN.scala 248:22]
  assign _expOut_T = io_in_isZero | common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 251:32]
  assign _expOut_T_1 = _expOut_T ? 9'h1c0 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 251:18]
  assign _expOut_T_3 = common_expOut & ~_expOut_T_1; // @[RoundAnyRawFNToRecFN.scala 250:24]
  assign _expOut_T_5 = pegMinNonzeroMagOut ? 9'h194 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 255:18]
  assign _expOut_T_7 = _expOut_T_3 & ~_expOut_T_5; // @[RoundAnyRawFNToRecFN.scala 254:17]
  assign _expOut_T_8 = pegMaxFiniteMagOut ? 9'h80 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 259:18]
  assign _expOut_T_10 = _expOut_T_7 & ~_expOut_T_8; // @[RoundAnyRawFNToRecFN.scala 258:17]
  assign _expOut_T_11 = notNaN_isInfOut ? 9'h40 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 263:18]
  assign _expOut_T_13 = _expOut_T_10 & ~_expOut_T_11; // @[RoundAnyRawFNToRecFN.scala 262:17]
  assign _expOut_T_14 = pegMinNonzeroMagOut ? 9'h6b : 9'h0; // @[RoundAnyRawFNToRecFN.scala 267:16]
  assign _expOut_T_15 = _expOut_T_13 | _expOut_T_14; // @[RoundAnyRawFNToRecFN.scala 266:18]
  assign _expOut_T_16 = pegMaxFiniteMagOut ? 9'h17f : 9'h0; // @[RoundAnyRawFNToRecFN.scala 271:16]
  assign _expOut_T_17 = _expOut_T_15 | _expOut_T_16; // @[RoundAnyRawFNToRecFN.scala 270:15]
  assign _expOut_T_18 = notNaN_isInfOut ? 9'h180 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 275:16]
  assign _expOut_T_19 = _expOut_T_17 | _expOut_T_18; // @[RoundAnyRawFNToRecFN.scala 274:15]
  assign _expOut_T_20 = isNaNOut ? 9'h1c0 : 9'h0; // @[RoundAnyRawFNToRecFN.scala 276:16]
  assign expOut = _expOut_T_19 | _expOut_T_20; // @[RoundAnyRawFNToRecFN.scala 275:77]
  assign _fractOut_T = isNaNOut | io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 278:22]
  assign _fractOut_T_1 = _fractOut_T | common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 278:38]
  assign _fractOut_T_2 = isNaNOut ? 23'h400000 : 23'h0; // @[RoundAnyRawFNToRecFN.scala 279:16]
  assign _fractOut_T_3 = _fractOut_T_1 ? _fractOut_T_2 : common_fractOut; // @[RoundAnyRawFNToRecFN.scala 278:12]
  assign _fractOut_T_5 = pegMaxFiniteMagOut ? 23'h7fffff : 23'h0; // @[Bitwise.scala 72:12]
  assign fractOut = _fractOut_T_3 | _fractOut_T_5; // @[RoundAnyRawFNToRecFN.scala 281:11]
  assign io_out_hi = {signOut,expOut}; // @[Cat.scala 30:58]
  assign io_exceptionFlags_lo = {underflow,inexact}; // @[Cat.scala 30:58]
  assign io_exceptionFlags_hi = {io_invalidExc,io_infiniteExc,overflow}; // @[Cat.scala 30:58]
  assign io_out = {io_out_hi,fractOut}; // @[RoundAnyRawFNToRecFN.scala 284:12]
  assign io_exceptionFlags = {io_exceptionFlags_hi,io_exceptionFlags_lo}; // @[RoundAnyRawFNToRecFN.scala 285:23]
  assign RoundAnyRawFNToRecFN_5_covSum = 30'h0;
  assign io_covSum = RoundAnyRawFNToRecFN_5_covSum;
  assign metaAssert = 1'h0;
endmodule
module DivSqrtRawFN_small_1(
  input         clock,
  input         reset,
  output        io_inReady,
  input         io_inValid,
  input         io_sqrtOp,
  input         io_a_isNaN,
  input         io_a_isInf,
  input         io_a_isZero,
  input         io_a_sign,
  input  [12:0] io_a_sExp,
  input  [53:0] io_a_sig,
  input         io_b_isNaN,
  input         io_b_isInf,
  input         io_b_isZero,
  input         io_b_sign,
  input  [12:0] io_b_sExp,
  input  [53:0] io_b_sig,
  input  [2:0]  io_roundingMode,
  output        io_rawOutValid_div,
  output        io_rawOutValid_sqrt,
  output [2:0]  io_roundingModeOut,
  output        io_invalidExc,
  output        io_infiniteExc,
  output        io_rawOut_isNaN,
  output        io_rawOut_isInf,
  output        io_rawOut_isZero,
  output        io_rawOut_sign,
  output [12:0] io_rawOut_sExp,
  output [55:0] io_rawOut_sig,
  output [29:0] io_covSum,
  output        metaAssert,
  input         metaReset
);
  reg [55:0] cycleNum; // @[DivSqrtRecFN_small.scala 223:33]
  reg [63:0] _RAND_0;
  reg  sqrtOp_Z; // @[DivSqrtRecFN_small.scala 225:29]
  reg [31:0] _RAND_1;
  reg  majorExc_Z; // @[DivSqrtRecFN_small.scala 226:29]
  reg [31:0] _RAND_2;
  reg  isNaN_Z; // @[DivSqrtRecFN_small.scala 228:29]
  reg [31:0] _RAND_3;
  reg  isInf_Z; // @[DivSqrtRecFN_small.scala 229:29]
  reg [31:0] _RAND_4;
  reg  isZero_Z; // @[DivSqrtRecFN_small.scala 230:29]
  reg [31:0] _RAND_5;
  reg  sign_Z; // @[DivSqrtRecFN_small.scala 231:29]
  reg [31:0] _RAND_6;
  reg [12:0] sExp_Z; // @[DivSqrtRecFN_small.scala 232:29]
  reg [31:0] _RAND_7;
  reg [51:0] fractB_Z; // @[DivSqrtRecFN_small.scala 233:29]
  reg [63:0] _RAND_8;
  reg [2:0] roundingMode_Z; // @[DivSqrtRecFN_small.scala 234:29]
  reg [31:0] _RAND_9;
  reg [54:0] rem_Z; // @[DivSqrtRecFN_small.scala 240:29]
  reg [63:0] _RAND_10;
  reg  notZeroRem_Z; // @[DivSqrtRecFN_small.scala 241:29]
  reg [31:0] _RAND_11;
  reg [54:0] sigX_Z; // @[DivSqrtRecFN_small.scala 242:29]
  reg [63:0] _RAND_12;
  wire  _notSigNaNIn_invalidExc_S_div_T; // @[DivSqrtRecFN_small.scala 251:24]
  wire  _notSigNaNIn_invalidExc_S_div_T_1; // @[DivSqrtRecFN_small.scala 251:59]
  wire  notSigNaNIn_invalidExc_S_div; // @[DivSqrtRecFN_small.scala 251:42]
  wire  _notSigNaNIn_invalidExc_S_sqrt_T_2; // @[DivSqrtRecFN_small.scala 253:24]
  wire  notSigNaNIn_invalidExc_S_sqrt; // @[DivSqrtRecFN_small.scala 253:43]
  wire  _majorExc_S_T_2; // @[common.scala 81:46]
  wire  _majorExc_S_T_3; // @[DivSqrtRecFN_small.scala 256:38]
  wire  _majorExc_S_T_9; // @[common.scala 81:46]
  wire  _majorExc_S_T_10; // @[DivSqrtRecFN_small.scala 257:38]
  wire  _majorExc_S_T_11; // @[DivSqrtRecFN_small.scala 257:66]
  wire  _majorExc_S_T_14; // @[DivSqrtRecFN_small.scala 259:33]
  wire  _majorExc_S_T_15; // @[DivSqrtRecFN_small.scala 259:51]
  wire  _majorExc_S_T_16; // @[DivSqrtRecFN_small.scala 258:46]
  wire  _isNaN_S_T; // @[DivSqrtRecFN_small.scala 263:26]
  wire  _isNaN_S_T_1; // @[DivSqrtRecFN_small.scala 264:26]
  wire  _isNaN_S_T_2; // @[DivSqrtRecFN_small.scala 264:42]
  wire  _isInf_S_T; // @[DivSqrtRecFN_small.scala 266:63]
  wire  _isZero_S_T; // @[DivSqrtRecFN_small.scala 267:64]
  wire  _sign_S_T_1; // @[DivSqrtRecFN_small.scala 268:45]
  wire  sign_S; // @[DivSqrtRecFN_small.scala 268:30]
  wire  _specialCaseA_S_T; // @[DivSqrtRecFN_small.scala 270:39]
  wire  specialCaseA_S; // @[DivSqrtRecFN_small.scala 270:55]
  wire  _specialCaseB_S_T; // @[DivSqrtRecFN_small.scala 271:39]
  wire  specialCaseB_S; // @[DivSqrtRecFN_small.scala 271:55]
  wire  normalCase_S_div; // @[DivSqrtRecFN_small.scala 272:45]
  wire  normalCase_S_sqrt; // @[DivSqrtRecFN_small.scala 273:46]
  wire  normalCase_S; // @[DivSqrtRecFN_small.scala 274:27]
  wire  sExpQuot_S_div_hi; // @[DivSqrtRecFN_small.scala 278:28]
  wire [10:0] sExpQuot_S_div_lo; // @[DivSqrtRecFN_small.scala 278:40]
  wire [11:0] _sExpQuot_S_div_T_2; // @[DivSqrtRecFN_small.scala 278:71]
  wire [12:0] _GEN_13; // @[DivSqrtRecFN_small.scala 277:21]
  wire [13:0] sExpQuot_S_div; // @[DivSqrtRecFN_small.scala 277:21]
  wire  _sSatExpQuot_S_div_T; // @[DivSqrtRecFN_small.scala 281:48]
  wire [3:0] sSatExpQuot_S_div_hi; // @[DivSqrtRecFN_small.scala 281:16]
  wire [8:0] sSatExpQuot_S_div_lo; // @[DivSqrtRecFN_small.scala 285:27]
  wire [12:0] sSatExpQuot_S_div; // @[DivSqrtRecFN_small.scala 286:11]
  wire  evenSqrt_S; // @[DivSqrtRecFN_small.scala 288:32]
  wire  oddSqrt_S; // @[DivSqrtRecFN_small.scala 289:32]
  wire  idle; // @[DivSqrtRecFN_small.scala 293:24]
  wire  inReady; // @[DivSqrtRecFN_small.scala 294:24]
  wire  entering; // @[DivSqrtRecFN_small.scala 295:28]
  wire  entering_normalCase; // @[DivSqrtRecFN_small.scala 296:40]
  wire  skipCycle2; // @[DivSqrtRecFN_small.scala 298:34]
  wire  _T_1; // @[DivSqrtRecFN_small.scala 300:18]
  wire  _cycleNum_T_1; // @[DivSqrtRecFN_small.scala 302:26]
  wire [1:0] _cycleNum_T_2; // @[DivSqrtRecFN_small.scala 302:16]
  wire [54:0] _cycleNum_T_4; // @[DivSqrtRecFN_small.scala 305:24]
  wire [55:0] _cycleNum_T_5; // @[DivSqrtRecFN_small.scala 304:20]
  wire [55:0] _cycleNum_T_6; // @[DivSqrtRecFN_small.scala 303:16]
  wire [55:0] _GEN_14; // @[DivSqrtRecFN_small.scala 302:59]
  wire [55:0] _cycleNum_T_7; // @[DivSqrtRecFN_small.scala 302:59]
  wire  _cycleNum_T_10; // @[DivSqrtRecFN_small.scala 310:28]
  wire [54:0] _cycleNum_T_12; // @[DivSqrtRecFN_small.scala 310:16]
  wire [55:0] _GEN_15; // @[DivSqrtRecFN_small.scala 309:15]
  wire [55:0] _cycleNum_T_13; // @[DivSqrtRecFN_small.scala 309:15]
  wire [1:0] _cycleNum_T_14; // @[DivSqrtRecFN_small.scala 311:16]
  wire [55:0] _GEN_16; // @[DivSqrtRecFN_small.scala 310:63]
  wire [55:0] _cycleNum_T_15; // @[DivSqrtRecFN_small.scala 310:63]
  wire [11:0] _sExp_Z_T; // @[DivSqrtRecFN_small.scala 329:29]
  wire [12:0] _sExp_Z_T_1; // @[DivSqrtRecFN_small.scala 329:34]
  wire  _T_3; // @[DivSqrtRecFN_small.scala 334:31]
  wire  _rem_T_1; // @[DivSqrtRecFN_small.scala 341:21]
  wire [54:0] _rem_T_2; // @[DivSqrtRecFN_small.scala 341:47]
  wire [54:0] _rem_T_3; // @[DivSqrtRecFN_small.scala 341:12]
  wire  _rem_T_4; // @[DivSqrtRecFN_small.scala 342:21]
  wire [1:0] rem_hi; // @[DivSqrtRecFN_small.scala 343:56]
  wire [53:0] rem_lo; // @[DivSqrtRecFN_small.scala 344:44]
  wire [55:0] _rem_T_8; // @[Cat.scala 30:58]
  wire [55:0] _rem_T_9; // @[DivSqrtRecFN_small.scala 342:12]
  wire [55:0] _GEN_17; // @[DivSqrtRecFN_small.scala 341:57]
  wire [55:0] _rem_T_10; // @[DivSqrtRecFN_small.scala 341:57]
  wire [55:0] _rem_T_12; // @[DivSqrtRecFN_small.scala 348:29]
  wire [55:0] _rem_T_13; // @[DivSqrtRecFN_small.scala 348:12]
  wire [55:0] rem; // @[DivSqrtRecFN_small.scala 347:11]
  wire [53:0] bitMask; // @[DivSqrtRecFN_small.scala 349:27]
  wire  _trialTerm_T_1; // @[DivSqrtRecFN_small.scala 351:21]
  wire [54:0] _trialTerm_T_2; // @[DivSqrtRecFN_small.scala 351:47]
  wire [54:0] _trialTerm_T_3; // @[DivSqrtRecFN_small.scala 351:12]
  wire  _trialTerm_T_4; // @[DivSqrtRecFN_small.scala 352:21]
  wire [53:0] _trialTerm_T_5; // @[DivSqrtRecFN_small.scala 352:12]
  wire [54:0] _GEN_18; // @[DivSqrtRecFN_small.scala 351:73]
  wire [54:0] _trialTerm_T_6; // @[DivSqrtRecFN_small.scala 351:73]
  wire [54:0] _trialTerm_T_8; // @[DivSqrtRecFN_small.scala 353:12]
  wire [54:0] _trialTerm_T_9; // @[DivSqrtRecFN_small.scala 352:73]
  wire  _trialTerm_T_12; // @[DivSqrtRecFN_small.scala 354:23]
  wire [52:0] _trialTerm_T_13; // @[Cat.scala 30:58]
  wire [53:0] _trialTerm_T_14; // @[DivSqrtRecFN_small.scala 354:56]
  wire [53:0] _trialTerm_T_15; // @[DivSqrtRecFN_small.scala 354:12]
  wire [54:0] _GEN_19; // @[DivSqrtRecFN_small.scala 353:73]
  wire [54:0] _trialTerm_T_16; // @[DivSqrtRecFN_small.scala 353:73]
  wire  _trialTerm_T_18; // @[DivSqrtRecFN_small.scala 355:23]
  wire [55:0] _trialTerm_T_19; // @[DivSqrtRecFN_small.scala 355:44]
  wire [55:0] _GEN_20; // @[DivSqrtRecFN_small.scala 355:48]
  wire [55:0] _trialTerm_T_20; // @[DivSqrtRecFN_small.scala 355:48]
  wire [55:0] _trialTerm_T_21; // @[DivSqrtRecFN_small.scala 355:12]
  wire [55:0] _GEN_21; // @[DivSqrtRecFN_small.scala 354:73]
  wire [55:0] trialTerm; // @[DivSqrtRecFN_small.scala 354:73]
  wire [56:0] _trialRem_T; // @[DivSqrtRecFN_small.scala 356:24]
  wire [56:0] _trialRem_T_1; // @[DivSqrtRecFN_small.scala 356:41]
  wire [56:0] trialRem; // @[DivSqrtRecFN_small.scala 356:29]
  wire  newBit; // @[DivSqrtRecFN_small.scala 357:23]
  wire  _T_5; // @[DivSqrtRecFN_small.scala 359:41]
  wire  _T_7; // @[DivSqrtRecFN_small.scala 359:31]
  wire [56:0] _rem_Z_T; // @[DivSqrtRecFN_small.scala 360:39]
  wire [56:0] _rem_Z_T_1; // @[DivSqrtRecFN_small.scala 360:21]
  wire [56:0] _GEN_10; // @[DivSqrtRecFN_small.scala 359:58]
  wire  _T_9; // @[DivSqrtRecFN_small.scala 362:45]
  wire  _T_10; // @[DivSqrtRecFN_small.scala 362:31]
  wire  _notZeroRem_Z_T; // @[DivSqrtRecFN_small.scala 363:35]
  wire [54:0] _sigX_Z_T_2; // @[DivSqrtRecFN_small.scala 365:47]
  wire [54:0] _sigX_Z_T_3; // @[DivSqrtRecFN_small.scala 365:16]
  wire  _sigX_Z_T_4; // @[DivSqrtRecFN_small.scala 366:25]
  wire [53:0] _sigX_Z_T_5; // @[DivSqrtRecFN_small.scala 366:16]
  wire [54:0] _GEN_22; // @[DivSqrtRecFN_small.scala 365:71]
  wire [54:0] _sigX_Z_T_6; // @[DivSqrtRecFN_small.scala 365:71]
  wire [52:0] _sigX_Z_T_8; // @[DivSqrtRecFN_small.scala 367:47]
  wire [52:0] _sigX_Z_T_9; // @[DivSqrtRecFN_small.scala 367:16]
  wire [54:0] _GEN_23; // @[DivSqrtRecFN_small.scala 366:71]
  wire [54:0] _sigX_Z_T_10; // @[DivSqrtRecFN_small.scala 366:71]
  wire [54:0] _GEN_24; // @[DivSqrtRecFN_small.scala 368:48]
  wire [54:0] _sigX_Z_T_12; // @[DivSqrtRecFN_small.scala 368:48]
  wire [54:0] _sigX_Z_T_13; // @[DivSqrtRecFN_small.scala 368:16]
  wire [54:0] _sigX_Z_T_14; // @[DivSqrtRecFN_small.scala 367:71]
  wire [55:0] _GEN_25; // @[DivSqrtRecFN_small.scala 385:35]
  reg [4:0] DivSqrtRawFN_small_1_state; // @[Register tracking DivSqrtRawFN_small_1 state]
  reg [31:0] _RAND_13;
  reg  DivSqrtRawFN_small_1_cov [0:31]; // @[Coverage map for DivSqrtRawFN_small_1]
  reg [31:0] _RAND_14;
  wire  DivSqrtRawFN_small_1_cov_read_data; // @[Coverage map for DivSqrtRawFN_small_1]
  wire [4:0] DivSqrtRawFN_small_1_cov_read_addr; // @[Coverage map for DivSqrtRawFN_small_1]
  wire  DivSqrtRawFN_small_1_cov_write_data; // @[Coverage map for DivSqrtRawFN_small_1]
  wire [4:0] DivSqrtRawFN_small_1_cov_write_addr; // @[Coverage map for DivSqrtRawFN_small_1]
  wire  DivSqrtRawFN_small_1_cov_write_mask; // @[Coverage map for DivSqrtRawFN_small_1]
  wire  DivSqrtRawFN_small_1_cov_write_en; // @[Coverage map for DivSqrtRawFN_small_1]
  reg [29:0] DivSqrtRawFN_small_1_covSum; // @[Sum of coverage map]
  reg [31:0] _RAND_15;
  wire  mux_cond_0;
  wire  mux_cond_1;
  wire  mux_cond_2;
  wire  mux_cond_3;
  wire  sqrtOp_Z_shl;
  wire [4:0] sqrtOp_Z_pad;
  wire [1:0] mux_cond_0_shl;
  wire [4:0] mux_cond_0_pad;
  wire [2:0] mux_cond_1_shl;
  wire [4:0] mux_cond_1_pad;
  wire [3:0] mux_cond_2_shl;
  wire [4:0] mux_cond_2_pad;
  wire [4:0] mux_cond_3_shl;
  wire [4:0] mux_cond_3_pad;
  wire [4:0] DivSqrtRawFN_small_1_xor1;
  wire [4:0] DivSqrtRawFN_small_1_xor6;
  wire [4:0] DivSqrtRawFN_small_1_xor2;
  wire [4:0] DivSqrtRawFN_small_1_xor0;
  assign _notSigNaNIn_invalidExc_S_div_T = io_a_isZero & io_b_isZero; // @[DivSqrtRecFN_small.scala 251:24]
  assign _notSigNaNIn_invalidExc_S_div_T_1 = io_a_isInf & io_b_isInf; // @[DivSqrtRecFN_small.scala 251:59]
  assign notSigNaNIn_invalidExc_S_div = _notSigNaNIn_invalidExc_S_div_T | _notSigNaNIn_invalidExc_S_div_T_1; // @[DivSqrtRecFN_small.scala 251:42]
  assign _notSigNaNIn_invalidExc_S_sqrt_T_2 = ~io_a_isNaN & ~io_a_isZero; // @[DivSqrtRecFN_small.scala 253:24]
  assign notSigNaNIn_invalidExc_S_sqrt = _notSigNaNIn_invalidExc_S_sqrt_T_2 & io_a_sign; // @[DivSqrtRecFN_small.scala 253:43]
  assign _majorExc_S_T_2 = io_a_isNaN & ~io_a_sig[51]; // @[common.scala 81:46]
  assign _majorExc_S_T_3 = _majorExc_S_T_2 | notSigNaNIn_invalidExc_S_sqrt; // @[DivSqrtRecFN_small.scala 256:38]
  assign _majorExc_S_T_9 = io_b_isNaN & ~io_b_sig[51]; // @[common.scala 81:46]
  assign _majorExc_S_T_10 = _majorExc_S_T_2 | _majorExc_S_T_9; // @[DivSqrtRecFN_small.scala 257:38]
  assign _majorExc_S_T_11 = _majorExc_S_T_10 | notSigNaNIn_invalidExc_S_div; // @[DivSqrtRecFN_small.scala 257:66]
  assign _majorExc_S_T_14 = ~io_a_isNaN & ~io_a_isInf; // @[DivSqrtRecFN_small.scala 259:33]
  assign _majorExc_S_T_15 = _majorExc_S_T_14 & io_b_isZero; // @[DivSqrtRecFN_small.scala 259:51]
  assign _majorExc_S_T_16 = _majorExc_S_T_11 | _majorExc_S_T_15; // @[DivSqrtRecFN_small.scala 258:46]
  assign _isNaN_S_T = io_a_isNaN | notSigNaNIn_invalidExc_S_sqrt; // @[DivSqrtRecFN_small.scala 263:26]
  assign _isNaN_S_T_1 = io_a_isNaN | io_b_isNaN; // @[DivSqrtRecFN_small.scala 264:26]
  assign _isNaN_S_T_2 = _isNaN_S_T_1 | notSigNaNIn_invalidExc_S_div; // @[DivSqrtRecFN_small.scala 264:42]
  assign _isInf_S_T = io_a_isInf | io_b_isZero; // @[DivSqrtRecFN_small.scala 266:63]
  assign _isZero_S_T = io_a_isZero | io_b_isInf; // @[DivSqrtRecFN_small.scala 267:64]
  assign _sign_S_T_1 = ~io_sqrtOp & io_b_sign; // @[DivSqrtRecFN_small.scala 268:45]
  assign sign_S = io_a_sign ^ _sign_S_T_1; // @[DivSqrtRecFN_small.scala 268:30]
  assign _specialCaseA_S_T = io_a_isNaN | io_a_isInf; // @[DivSqrtRecFN_small.scala 270:39]
  assign specialCaseA_S = _specialCaseA_S_T | io_a_isZero; // @[DivSqrtRecFN_small.scala 270:55]
  assign _specialCaseB_S_T = io_b_isNaN | io_b_isInf; // @[DivSqrtRecFN_small.scala 271:39]
  assign specialCaseB_S = _specialCaseB_S_T | io_b_isZero; // @[DivSqrtRecFN_small.scala 271:55]
  assign normalCase_S_div = ~specialCaseA_S & ~specialCaseB_S; // @[DivSqrtRecFN_small.scala 272:45]
  assign normalCase_S_sqrt = ~specialCaseA_S & ~io_a_sign; // @[DivSqrtRecFN_small.scala 273:46]
  assign normalCase_S = io_sqrtOp ? normalCase_S_sqrt : normalCase_S_div; // @[DivSqrtRecFN_small.scala 274:27]
  assign sExpQuot_S_div_hi = io_b_sExp[11]; // @[DivSqrtRecFN_small.scala 278:28]
  assign sExpQuot_S_div_lo = ~io_b_sExp[10:0]; // @[DivSqrtRecFN_small.scala 278:40]
  assign _sExpQuot_S_div_T_2 = {sExpQuot_S_div_hi,sExpQuot_S_div_lo}; // @[DivSqrtRecFN_small.scala 278:71]
  assign _GEN_13 = {{1{_sExpQuot_S_div_T_2[11]}},_sExpQuot_S_div_T_2}; // @[DivSqrtRecFN_small.scala 277:21]
  assign sExpQuot_S_div = $signed(io_a_sExp) + $signed(_GEN_13); // @[DivSqrtRecFN_small.scala 277:21]
  assign _sSatExpQuot_S_div_T = 14'she00 <= $signed(sExpQuot_S_div); // @[DivSqrtRecFN_small.scala 281:48]
  assign sSatExpQuot_S_div_hi = _sSatExpQuot_S_div_T ? 4'h6 : sExpQuot_S_div[12:9]; // @[DivSqrtRecFN_small.scala 281:16]
  assign sSatExpQuot_S_div_lo = sExpQuot_S_div[8:0]; // @[DivSqrtRecFN_small.scala 285:27]
  assign sSatExpQuot_S_div = {sSatExpQuot_S_div_hi,sSatExpQuot_S_div_lo}; // @[DivSqrtRecFN_small.scala 286:11]
  assign evenSqrt_S = io_sqrtOp & ~io_a_sExp[0]; // @[DivSqrtRecFN_small.scala 288:32]
  assign oddSqrt_S = io_sqrtOp & io_a_sExp[0]; // @[DivSqrtRecFN_small.scala 289:32]
  assign idle = cycleNum[0]; // @[DivSqrtRecFN_small.scala 293:24]
  assign inReady = idle | cycleNum[1]; // @[DivSqrtRecFN_small.scala 294:24]
  assign entering = inReady & io_inValid; // @[DivSqrtRecFN_small.scala 295:28]
  assign entering_normalCase = entering & normalCase_S; // @[DivSqrtRecFN_small.scala 296:40]
  assign skipCycle2 = cycleNum[3] & sigX_Z[54]; // @[DivSqrtRecFN_small.scala 298:34]
  assign _T_1 = ~idle | entering; // @[DivSqrtRecFN_small.scala 300:18]
  assign _cycleNum_T_1 = entering & ~normalCase_S; // @[DivSqrtRecFN_small.scala 302:26]
  assign _cycleNum_T_2 = _cycleNum_T_1 ? 2'h2 : 2'h0; // @[DivSqrtRecFN_small.scala 302:16]
  assign _cycleNum_T_4 = io_a_sExp[0] ? 55'h20000000000000 : 55'h40000000000000; // @[DivSqrtRecFN_small.scala 305:24]
  assign _cycleNum_T_5 = io_sqrtOp ? {{1'd0}, _cycleNum_T_4} : 56'h80000000000000; // @[DivSqrtRecFN_small.scala 304:20]
  assign _cycleNum_T_6 = entering_normalCase ? _cycleNum_T_5 : 56'h0; // @[DivSqrtRecFN_small.scala 303:16]
  assign _GEN_14 = {{54'd0}, _cycleNum_T_2}; // @[DivSqrtRecFN_small.scala 302:59]
  assign _cycleNum_T_7 = _GEN_14 | _cycleNum_T_6; // @[DivSqrtRecFN_small.scala 302:59]
  assign _cycleNum_T_10 = ~entering & ~skipCycle2; // @[DivSqrtRecFN_small.scala 310:28]
  assign _cycleNum_T_12 = _cycleNum_T_10 ? cycleNum[55:1] : 55'h0; // @[DivSqrtRecFN_small.scala 310:16]
  assign _GEN_15 = {{1'd0}, _cycleNum_T_12}; // @[DivSqrtRecFN_small.scala 309:15]
  assign _cycleNum_T_13 = _cycleNum_T_7 | _GEN_15; // @[DivSqrtRecFN_small.scala 309:15]
  assign _cycleNum_T_14 = skipCycle2 ? 2'h2 : 2'h0; // @[DivSqrtRecFN_small.scala 311:16]
  assign _GEN_16 = {{54'd0}, _cycleNum_T_14}; // @[DivSqrtRecFN_small.scala 310:63]
  assign _cycleNum_T_15 = _cycleNum_T_13 | _GEN_16; // @[DivSqrtRecFN_small.scala 310:63]
  assign _sExp_Z_T = io_a_sExp[12:1]; // @[DivSqrtRecFN_small.scala 329:29]
  assign _sExp_Z_T_1 = $signed(_sExp_Z_T) + 12'sh400; // @[DivSqrtRecFN_small.scala 329:34]
  assign _T_3 = entering_normalCase & ~io_sqrtOp; // @[DivSqrtRecFN_small.scala 334:31]
  assign _rem_T_1 = inReady & ~oddSqrt_S; // @[DivSqrtRecFN_small.scala 341:21]
  assign _rem_T_2 = {io_a_sig, 1'h0}; // @[DivSqrtRecFN_small.scala 341:47]
  assign _rem_T_3 = _rem_T_1 ? _rem_T_2 : 55'h0; // @[DivSqrtRecFN_small.scala 341:12]
  assign _rem_T_4 = inReady & oddSqrt_S; // @[DivSqrtRecFN_small.scala 342:21]
  assign rem_hi = io_a_sig[52:51] - 2'h1; // @[DivSqrtRecFN_small.scala 343:56]
  assign rem_lo = {io_a_sig[50:0], 3'h0}; // @[DivSqrtRecFN_small.scala 344:44]
  assign _rem_T_8 = {rem_hi,rem_lo}; // @[Cat.scala 30:58]
  assign _rem_T_9 = _rem_T_4 ? _rem_T_8 : 56'h0; // @[DivSqrtRecFN_small.scala 342:12]
  assign _GEN_17 = {{1'd0}, _rem_T_3}; // @[DivSqrtRecFN_small.scala 341:57]
  assign _rem_T_10 = _GEN_17 | _rem_T_9; // @[DivSqrtRecFN_small.scala 341:57]
  assign _rem_T_12 = {rem_Z, 1'h0}; // @[DivSqrtRecFN_small.scala 348:29]
  assign _rem_T_13 = inReady ? 56'h0 : _rem_T_12; // @[DivSqrtRecFN_small.scala 348:12]
  assign rem = _rem_T_10 | _rem_T_13; // @[DivSqrtRecFN_small.scala 347:11]
  assign bitMask = cycleNum[55:2]; // @[DivSqrtRecFN_small.scala 349:27]
  assign _trialTerm_T_1 = inReady & ~io_sqrtOp; // @[DivSqrtRecFN_small.scala 351:21]
  assign _trialTerm_T_2 = {io_b_sig, 1'h0}; // @[DivSqrtRecFN_small.scala 351:47]
  assign _trialTerm_T_3 = _trialTerm_T_1 ? _trialTerm_T_2 : 55'h0; // @[DivSqrtRecFN_small.scala 351:12]
  assign _trialTerm_T_4 = inReady & evenSqrt_S; // @[DivSqrtRecFN_small.scala 352:21]
  assign _trialTerm_T_5 = _trialTerm_T_4 ? 54'h20000000000000 : 54'h0; // @[DivSqrtRecFN_small.scala 352:12]
  assign _GEN_18 = {{1'd0}, _trialTerm_T_5}; // @[DivSqrtRecFN_small.scala 351:73]
  assign _trialTerm_T_6 = _trialTerm_T_3 | _GEN_18; // @[DivSqrtRecFN_small.scala 351:73]
  assign _trialTerm_T_8 = _rem_T_4 ? 55'h50000000000000 : 55'h0; // @[DivSqrtRecFN_small.scala 353:12]
  assign _trialTerm_T_9 = _trialTerm_T_6 | _trialTerm_T_8; // @[DivSqrtRecFN_small.scala 352:73]
  assign _trialTerm_T_12 = ~inReady & ~sqrtOp_Z; // @[DivSqrtRecFN_small.scala 354:23]
  assign _trialTerm_T_13 = {1'h1,fractB_Z}; // @[Cat.scala 30:58]
  assign _trialTerm_T_14 = {_trialTerm_T_13, 1'h0}; // @[DivSqrtRecFN_small.scala 354:56]
  assign _trialTerm_T_15 = _trialTerm_T_12 ? _trialTerm_T_14 : 54'h0; // @[DivSqrtRecFN_small.scala 354:12]
  assign _GEN_19 = {{1'd0}, _trialTerm_T_15}; // @[DivSqrtRecFN_small.scala 353:73]
  assign _trialTerm_T_16 = _trialTerm_T_9 | _GEN_19; // @[DivSqrtRecFN_small.scala 353:73]
  assign _trialTerm_T_18 = ~inReady & sqrtOp_Z; // @[DivSqrtRecFN_small.scala 355:23]
  assign _trialTerm_T_19 = {sigX_Z, 1'h0}; // @[DivSqrtRecFN_small.scala 355:44]
  assign _GEN_20 = {{2'd0}, bitMask}; // @[DivSqrtRecFN_small.scala 355:48]
  assign _trialTerm_T_20 = _trialTerm_T_19 | _GEN_20; // @[DivSqrtRecFN_small.scala 355:48]
  assign _trialTerm_T_21 = _trialTerm_T_18 ? _trialTerm_T_20 : 56'h0; // @[DivSqrtRecFN_small.scala 355:12]
  assign _GEN_21 = {{1'd0}, _trialTerm_T_16}; // @[DivSqrtRecFN_small.scala 354:73]
  assign trialTerm = _GEN_21 | _trialTerm_T_21; // @[DivSqrtRecFN_small.scala 354:73]
  assign _trialRem_T = {1'b0,$signed(rem)}; // @[DivSqrtRecFN_small.scala 356:24]
  assign _trialRem_T_1 = {1'b0,$signed(trialTerm)}; // @[DivSqrtRecFN_small.scala 356:41]
  assign trialRem = $signed(_trialRem_T) - $signed(_trialRem_T_1); // @[DivSqrtRecFN_small.scala 356:29]
  assign newBit = 57'sh0 <= $signed(trialRem); // @[DivSqrtRecFN_small.scala 357:23]
  assign _T_5 = idle | cycleNum[2]; // @[DivSqrtRecFN_small.scala 359:41]
  assign _T_7 = entering_normalCase | ~_T_5; // @[DivSqrtRecFN_small.scala 359:31]
  assign _rem_Z_T = $signed(_trialRem_T) - $signed(_trialRem_T_1); // @[DivSqrtRecFN_small.scala 360:39]
  assign _rem_Z_T_1 = newBit ? _rem_Z_T : {{1'd0}, rem}; // @[DivSqrtRecFN_small.scala 360:21]
  assign _GEN_10 = _T_7 ? _rem_Z_T_1 : {{2'd0}, rem_Z}; // @[DivSqrtRecFN_small.scala 359:58]
  assign _T_9 = ~inReady & newBit; // @[DivSqrtRecFN_small.scala 362:45]
  assign _T_10 = entering_normalCase | _T_9; // @[DivSqrtRecFN_small.scala 362:31]
  assign _notZeroRem_Z_T = $signed(trialRem) != 57'sh0; // @[DivSqrtRecFN_small.scala 363:35]
  assign _sigX_Z_T_2 = {newBit, 54'h0}; // @[DivSqrtRecFN_small.scala 365:47]
  assign _sigX_Z_T_3 = _trialTerm_T_1 ? _sigX_Z_T_2 : 55'h0; // @[DivSqrtRecFN_small.scala 365:16]
  assign _sigX_Z_T_4 = inReady & io_sqrtOp; // @[DivSqrtRecFN_small.scala 366:25]
  assign _sigX_Z_T_5 = _sigX_Z_T_4 ? 54'h20000000000000 : 54'h0; // @[DivSqrtRecFN_small.scala 366:16]
  assign _GEN_22 = {{1'd0}, _sigX_Z_T_5}; // @[DivSqrtRecFN_small.scala 365:71]
  assign _sigX_Z_T_6 = _sigX_Z_T_3 | _GEN_22; // @[DivSqrtRecFN_small.scala 365:71]
  assign _sigX_Z_T_8 = {newBit, 52'h0}; // @[DivSqrtRecFN_small.scala 367:47]
  assign _sigX_Z_T_9 = _rem_T_4 ? _sigX_Z_T_8 : 53'h0; // @[DivSqrtRecFN_small.scala 367:16]
  assign _GEN_23 = {{2'd0}, _sigX_Z_T_9}; // @[DivSqrtRecFN_small.scala 366:71]
  assign _sigX_Z_T_10 = _sigX_Z_T_6 | _GEN_23; // @[DivSqrtRecFN_small.scala 366:71]
  assign _GEN_24 = {{1'd0}, bitMask}; // @[DivSqrtRecFN_small.scala 368:48]
  assign _sigX_Z_T_12 = sigX_Z | _GEN_24; // @[DivSqrtRecFN_small.scala 368:48]
  assign _sigX_Z_T_13 = inReady ? 55'h0 : _sigX_Z_T_12; // @[DivSqrtRecFN_small.scala 368:16]
  assign _sigX_Z_T_14 = _sigX_Z_T_10 | _sigX_Z_T_13; // @[DivSqrtRecFN_small.scala 367:71]
  assign _GEN_25 = {{55'd0}, notZeroRem_Z}; // @[DivSqrtRecFN_small.scala 385:35]
  assign io_inReady = idle | cycleNum[1]; // @[DivSqrtRecFN_small.scala 314:16]
  assign io_rawOutValid_div = cycleNum[1] & ~sqrtOp_Z; // @[DivSqrtRecFN_small.scala 375:25]
  assign io_rawOutValid_sqrt = cycleNum[1] & sqrtOp_Z; // @[DivSqrtRecFN_small.scala 376:25]
  assign io_roundingModeOut = roundingMode_Z; // @[DivSqrtRecFN_small.scala 377:25]
  assign io_invalidExc = majorExc_Z & isNaN_Z; // @[DivSqrtRecFN_small.scala 378:22]
  assign io_infiniteExc = majorExc_Z & ~isNaN_Z; // @[DivSqrtRecFN_small.scala 379:22]
  assign io_rawOut_isNaN = isNaN_Z; // @[DivSqrtRecFN_small.scala 380:22]
  assign io_rawOut_isInf = isInf_Z; // @[DivSqrtRecFN_small.scala 381:22]
  assign io_rawOut_isZero = isZero_Z; // @[DivSqrtRecFN_small.scala 382:22]
  assign io_rawOut_sign = sign_Z; // @[DivSqrtRecFN_small.scala 383:22]
  assign io_rawOut_sExp = sExp_Z; // @[DivSqrtRecFN_small.scala 384:22]
  assign io_rawOut_sig = _trialTerm_T_19 | _GEN_25; // @[DivSqrtRecFN_small.scala 385:22]
  assign DivSqrtRawFN_small_1_cov_read_addr = DivSqrtRawFN_small_1_state;
  assign DivSqrtRawFN_small_1_cov_read_data = DivSqrtRawFN_small_1_cov[DivSqrtRawFN_small_1_cov_read_addr]; // @[Coverage map for DivSqrtRawFN_small_1]
  assign DivSqrtRawFN_small_1_cov_write_data = 1'h1;
  assign DivSqrtRawFN_small_1_cov_write_addr = DivSqrtRawFN_small_1_state;
  assign DivSqrtRawFN_small_1_cov_write_mask = 1'h1;
  assign DivSqrtRawFN_small_1_cov_write_en = 1'h1;
  assign mux_cond_0 = _T_10;
  assign mux_cond_1 = newBit;
  assign mux_cond_2 = skipCycle2;
  assign mux_cond_3 = _cycleNum_T_10;
  assign sqrtOp_Z_shl = sqrtOp_Z;
  assign sqrtOp_Z_pad = {4'h0,sqrtOp_Z_shl};
  assign mux_cond_0_shl = {mux_cond_0, 1'h0};
  assign mux_cond_0_pad = {3'h0,mux_cond_0_shl};
  assign mux_cond_1_shl = {mux_cond_1, 2'h0};
  assign mux_cond_1_pad = {2'h0,mux_cond_1_shl};
  assign mux_cond_2_shl = {mux_cond_2, 3'h0};
  assign mux_cond_2_pad = {1'h0,mux_cond_2_shl};
  assign mux_cond_3_shl = {mux_cond_3, 4'h0};
  assign mux_cond_3_pad = mux_cond_3_shl;
  assign DivSqrtRawFN_small_1_xor1 = sqrtOp_Z_pad ^ mux_cond_0_pad;
  assign DivSqrtRawFN_small_1_xor6 = mux_cond_2_pad ^ mux_cond_3_pad;
  assign DivSqrtRawFN_small_1_xor2 = mux_cond_1_pad ^ DivSqrtRawFN_small_1_xor6;
  assign DivSqrtRawFN_small_1_xor0 = DivSqrtRawFN_small_1_xor1 ^ DivSqrtRawFN_small_1_xor2;
  assign io_covSum = DivSqrtRawFN_small_1_covSum;
  assign metaAssert = 1'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  cycleNum = _RAND_0[55:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  sqrtOp_Z = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  majorExc_Z = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  isNaN_Z = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  isInf_Z = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  isZero_Z = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  sign_Z = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  sExp_Z = _RAND_7[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {2{`RANDOM}};
  fractB_Z = _RAND_8[51:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  roundingMode_Z = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {2{`RANDOM}};
  rem_Z = _RAND_10[54:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  notZeroRem_Z = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {2{`RANDOM}};
  sigX_Z = _RAND_12[54:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  DivSqrtRawFN_small_1_state = _RAND_13[4:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    DivSqrtRawFN_small_1_cov[initvar] = _RAND_14[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  DivSqrtRawFN_small_1_covSum = _RAND_15[29:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      cycleNum <= 56'h0;
    end else if (reset) begin
      cycleNum <= 56'h1;
    end else if (_T_1) begin
      cycleNum <= _cycleNum_T_15;
    end
    if (metaReset) begin
      sqrtOp_Z <= 1'h0;
    end else if (entering) begin
      sqrtOp_Z <= io_sqrtOp;
    end
    if (metaReset) begin
      majorExc_Z <= 1'h0;
    end else if (entering) begin
      if (io_sqrtOp) begin
        majorExc_Z <= _majorExc_S_T_3;
      end else begin
        majorExc_Z <= _majorExc_S_T_16;
      end
    end
    if (metaReset) begin
      isNaN_Z <= 1'h0;
    end else if (entering) begin
      if (io_sqrtOp) begin
        isNaN_Z <= _isNaN_S_T;
      end else begin
        isNaN_Z <= _isNaN_S_T_2;
      end
    end
    if (metaReset) begin
      isInf_Z <= 1'h0;
    end else if (entering) begin
      if (io_sqrtOp) begin
        isInf_Z <= io_a_isInf;
      end else begin
        isInf_Z <= _isInf_S_T;
      end
    end
    if (metaReset) begin
      isZero_Z <= 1'h0;
    end else if (entering) begin
      if (io_sqrtOp) begin
        isZero_Z <= io_a_isZero;
      end else begin
        isZero_Z <= _isZero_S_T;
      end
    end
    if (metaReset) begin
      sign_Z <= 1'h0;
    end else if (entering) begin
      sign_Z <= sign_S;
    end
    if (metaReset) begin
      sExp_Z <= 13'h0;
    end else if (entering_normalCase) begin
      if (io_sqrtOp) begin
        sExp_Z <= _sExp_Z_T_1;
      end else begin
        sExp_Z <= sSatExpQuot_S_div;
      end
    end
    if (metaReset) begin
      fractB_Z <= 52'h0;
    end else if (_T_3) begin
      fractB_Z <= io_b_sig[51:0];
    end
    if (metaReset) begin
      roundingMode_Z <= 3'h0;
    end else if (entering_normalCase) begin
      roundingMode_Z <= io_roundingMode;
    end
    if (metaReset) begin
      rem_Z <= 55'h0;
    end else begin
      rem_Z <= _GEN_10[54:0];
    end
    if (metaReset) begin
      notZeroRem_Z <= 1'h0;
    end else if (_T_10) begin
      notZeroRem_Z <= _notZeroRem_Z_T;
    end
    if (metaReset) begin
      sigX_Z <= 55'h0;
    end else if (_T_10) begin
      sigX_Z <= _sigX_Z_T_14;
    end
    DivSqrtRawFN_small_1_state <= DivSqrtRawFN_small_1_xor0;
    if (!(DivSqrtRawFN_small_1_cov_read_data)) begin
      DivSqrtRawFN_small_1_covSum <= DivSqrtRawFN_small_1_covSum + 1'h1;
    end
  end
  always @(posedge clock) begin
    if(DivSqrtRawFN_small_1_cov_write_en & DivSqrtRawFN_small_1_cov_write_mask) begin
      DivSqrtRawFN_small_1_cov[DivSqrtRawFN_small_1_cov_write_addr] <= DivSqrtRawFN_small_1_cov_write_data; // @[Coverage map for DivSqrtRawFN_small_1]
    end
  end
endmodule
module RoundAnyRawFNToRecFN_6(
  input         io_invalidExc,
  input         io_infiniteExc,
  input         io_in_isNaN,
  input         io_in_isInf,
  input         io_in_isZero,
  input         io_in_sign,
  input  [12:0] io_in_sExp,
  input  [55:0] io_in_sig,
  input  [2:0]  io_roundingMode,
  input         io_detectTininess,
  output [64:0] io_out,
  output [4:0]  io_exceptionFlags,
  output [29:0] io_covSum,
  output        metaAssert
);
  wire  roundingMode_near_even; // @[RoundAnyRawFNToRecFN.scala 88:53]
  wire  roundingMode_min; // @[RoundAnyRawFNToRecFN.scala 90:53]
  wire  roundingMode_max; // @[RoundAnyRawFNToRecFN.scala 91:53]
  wire  roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 92:53]
  wire  roundingMode_odd; // @[RoundAnyRawFNToRecFN.scala 93:53]
  wire  _roundMagUp_T; // @[RoundAnyRawFNToRecFN.scala 96:27]
  wire  _roundMagUp_T_2; // @[RoundAnyRawFNToRecFN.scala 96:63]
  wire  roundMagUp; // @[RoundAnyRawFNToRecFN.scala 96:42]
  wire  doShiftSigDown1; // @[RoundAnyRawFNToRecFN.scala 118:61]
  wire  roundMask_msb; // @[primitives.scala 57:25]
  wire [10:0] roundMask_lsbs; // @[primitives.scala 58:26]
  wire  roundMask_msb_1; // @[primitives.scala 57:25]
  wire [9:0] roundMask_lsbs_1; // @[primitives.scala 58:26]
  wire  roundMask_msb_2; // @[primitives.scala 57:25]
  wire [8:0] roundMask_lsbs_2; // @[primitives.scala 58:26]
  wire  roundMask_msb_3; // @[primitives.scala 57:25]
  wire [7:0] roundMask_lsbs_3; // @[primitives.scala 58:26]
  wire  roundMask_msb_4; // @[primitives.scala 57:25]
  wire [6:0] roundMask_lsbs_4; // @[primitives.scala 58:26]
  wire  roundMask_msb_5; // @[primitives.scala 57:25]
  wire [5:0] roundMask_lsbs_5; // @[primitives.scala 58:26]
  wire [64:0] roundMask_shift; // @[primitives.scala 77:58]
  wire [31:0] _roundMask_T_7; // @[Bitwise.scala 103:31]
  wire [31:0] _roundMask_T_9; // @[Bitwise.scala 103:65]
  wire [31:0] _roundMask_T_11; // @[Bitwise.scala 103:75]
  wire [31:0] _roundMask_T_12; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_0; // @[Bitwise.scala 103:31]
  wire [31:0] _roundMask_T_17; // @[Bitwise.scala 103:31]
  wire [31:0] _roundMask_T_19; // @[Bitwise.scala 103:65]
  wire [31:0] _roundMask_T_21; // @[Bitwise.scala 103:75]
  wire [31:0] _roundMask_T_22; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_1; // @[Bitwise.scala 103:31]
  wire [31:0] _roundMask_T_27; // @[Bitwise.scala 103:31]
  wire [31:0] _roundMask_T_29; // @[Bitwise.scala 103:65]
  wire [31:0] _roundMask_T_31; // @[Bitwise.scala 103:75]
  wire [31:0] _roundMask_T_32; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_2; // @[Bitwise.scala 103:31]
  wire [31:0] _roundMask_T_37; // @[Bitwise.scala 103:31]
  wire [31:0] _roundMask_T_39; // @[Bitwise.scala 103:65]
  wire [31:0] _roundMask_T_41; // @[Bitwise.scala 103:75]
  wire [31:0] _roundMask_T_42; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_3; // @[Bitwise.scala 103:31]
  wire [31:0] _roundMask_T_47; // @[Bitwise.scala 103:31]
  wire [31:0] _roundMask_T_49; // @[Bitwise.scala 103:65]
  wire [31:0] _roundMask_T_51; // @[Bitwise.scala 103:75]
  wire [31:0] roundMask_hi; // @[Bitwise.scala 103:39]
  wire [15:0] _roundMask_T_57; // @[Bitwise.scala 103:31]
  wire [15:0] _roundMask_T_59; // @[Bitwise.scala 103:65]
  wire [15:0] _roundMask_T_61; // @[Bitwise.scala 103:75]
  wire [15:0] _roundMask_T_62; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_4; // @[Bitwise.scala 103:31]
  wire [15:0] _roundMask_T_67; // @[Bitwise.scala 103:31]
  wire [15:0] _roundMask_T_69; // @[Bitwise.scala 103:65]
  wire [15:0] _roundMask_T_71; // @[Bitwise.scala 103:75]
  wire [15:0] _roundMask_T_72; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_5; // @[Bitwise.scala 103:31]
  wire [15:0] _roundMask_T_77; // @[Bitwise.scala 103:31]
  wire [15:0] _roundMask_T_79; // @[Bitwise.scala 103:65]
  wire [15:0] _roundMask_T_81; // @[Bitwise.scala 103:75]
  wire [15:0] _roundMask_T_82; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_6; // @[Bitwise.scala 103:31]
  wire [15:0] _roundMask_T_87; // @[Bitwise.scala 103:31]
  wire [15:0] _roundMask_T_89; // @[Bitwise.scala 103:65]
  wire [15:0] _roundMask_T_91; // @[Bitwise.scala 103:75]
  wire [15:0] roundMask_hi_1; // @[Bitwise.scala 103:39]
  wire  roundMask_hi_2; // @[Bitwise.scala 109:18]
  wire  roundMask_lo; // @[Bitwise.scala 109:44]
  wire  roundMask_lo_1; // @[Bitwise.scala 109:44]
  wire [50:0] _roundMask_T_94; // @[Cat.scala 30:58]
  wire [50:0] _roundMask_T_96; // @[primitives.scala 74:21]
  wire [50:0] _roundMask_T_99; // @[primitives.scala 74:21]
  wire [50:0] _roundMask_T_102; // @[primitives.scala 74:21]
  wire [50:0] _roundMask_T_105; // @[primitives.scala 74:21]
  wire [50:0] roundMask_hi_4; // @[primitives.scala 74:17]
  wire [53:0] _roundMask_T_106; // @[Cat.scala 30:58]
  wire  roundMask_hi_5; // @[Bitwise.scala 109:18]
  wire  roundMask_lo_4; // @[Bitwise.scala 109:44]
  wire  roundMask_lo_5; // @[Bitwise.scala 109:44]
  wire [2:0] _roundMask_T_109; // @[Cat.scala 30:58]
  wire [2:0] _roundMask_T_110; // @[primitives.scala 61:24]
  wire [2:0] _roundMask_T_111; // @[primitives.scala 61:24]
  wire [2:0] _roundMask_T_112; // @[primitives.scala 61:24]
  wire [2:0] _roundMask_T_113; // @[primitives.scala 61:24]
  wire [53:0] _roundMask_T_114; // @[primitives.scala 66:24]
  wire [53:0] _roundMask_T_115; // @[primitives.scala 61:24]
  wire [53:0] _GEN_7; // @[RoundAnyRawFNToRecFN.scala 157:23]
  wire [53:0] roundMask_hi_7; // @[RoundAnyRawFNToRecFN.scala 157:23]
  wire [55:0] roundMask; // @[Cat.scala 30:58]
  wire [54:0] shiftedRoundMask_lo; // @[RoundAnyRawFNToRecFN.scala 160:57]
  wire [55:0] shiftedRoundMask; // @[Cat.scala 30:58]
  wire [55:0] roundPosMask; // @[RoundAnyRawFNToRecFN.scala 161:46]
  wire [55:0] _roundPosBit_T; // @[RoundAnyRawFNToRecFN.scala 162:40]
  wire  roundPosBit; // @[RoundAnyRawFNToRecFN.scala 162:56]
  wire [55:0] _anyRoundExtra_T; // @[RoundAnyRawFNToRecFN.scala 163:42]
  wire  anyRoundExtra; // @[RoundAnyRawFNToRecFN.scala 163:62]
  wire  anyRound; // @[RoundAnyRawFNToRecFN.scala 164:36]
  wire  _roundIncr_T; // @[RoundAnyRawFNToRecFN.scala 167:38]
  wire  _roundIncr_T_1; // @[RoundAnyRawFNToRecFN.scala 167:67]
  wire  _roundIncr_T_2; // @[RoundAnyRawFNToRecFN.scala 169:29]
  wire  roundIncr; // @[RoundAnyRawFNToRecFN.scala 168:31]
  wire [55:0] _roundedSig_T; // @[RoundAnyRawFNToRecFN.scala 172:32]
  wire [54:0] _roundedSig_T_2; // @[RoundAnyRawFNToRecFN.scala 172:49]
  wire  _roundedSig_T_3; // @[RoundAnyRawFNToRecFN.scala 173:49]
  wire  _roundedSig_T_5; // @[RoundAnyRawFNToRecFN.scala 173:64]
  wire [54:0] _roundedSig_T_7; // @[RoundAnyRawFNToRecFN.scala 173:25]
  wire [54:0] _roundedSig_T_9; // @[RoundAnyRawFNToRecFN.scala 172:61]
  wire [55:0] _roundedSig_T_11; // @[RoundAnyRawFNToRecFN.scala 178:30]
  wire  _roundedSig_T_13; // @[RoundAnyRawFNToRecFN.scala 179:42]
  wire [54:0] _roundedSig_T_15; // @[RoundAnyRawFNToRecFN.scala 179:24]
  wire [54:0] _GEN_8; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [54:0] _roundedSig_T_16; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [54:0] roundedSig; // @[RoundAnyRawFNToRecFN.scala 171:16]
  wire [2:0] _sRoundedExp_T_1; // @[RoundAnyRawFNToRecFN.scala 183:69]
  wire [12:0] _GEN_9; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [13:0] sRoundedExp; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [11:0] common_expOut; // @[RoundAnyRawFNToRecFN.scala 185:37]
  wire [51:0] common_fractOut; // @[RoundAnyRawFNToRecFN.scala 187:16]
  wire [3:0] _common_overflow_T; // @[RoundAnyRawFNToRecFN.scala 194:30]
  wire  common_overflow; // @[RoundAnyRawFNToRecFN.scala 194:50]
  wire  common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 198:31]
  wire  unboundedRange_roundPosBit; // @[RoundAnyRawFNToRecFN.scala 201:16]
  wire  _unboundedRange_anyRound_T_1; // @[RoundAnyRawFNToRecFN.scala 203:30]
  wire  _unboundedRange_anyRound_T_3; // @[RoundAnyRawFNToRecFN.scala 203:70]
  wire  unboundedRange_anyRound; // @[RoundAnyRawFNToRecFN.scala 203:49]
  wire  _unboundedRange_roundIncr_T_1; // @[RoundAnyRawFNToRecFN.scala 205:67]
  wire  _unboundedRange_roundIncr_T_2; // @[RoundAnyRawFNToRecFN.scala 207:29]
  wire  unboundedRange_roundIncr; // @[RoundAnyRawFNToRecFN.scala 206:46]
  wire  roundCarry; // @[RoundAnyRawFNToRecFN.scala 209:16]
  wire [1:0] _common_underflow_T; // @[RoundAnyRawFNToRecFN.scala 218:48]
  wire  _common_underflow_T_1; // @[RoundAnyRawFNToRecFN.scala 218:62]
  wire  _common_underflow_T_2; // @[RoundAnyRawFNToRecFN.scala 218:32]
  wire  _common_underflow_T_5; // @[RoundAnyRawFNToRecFN.scala 219:30]
  wire  _common_underflow_T_6; // @[RoundAnyRawFNToRecFN.scala 218:74]
  wire  _common_underflow_T_10; // @[RoundAnyRawFNToRecFN.scala 221:39]
  wire  _common_underflow_T_12; // @[RoundAnyRawFNToRecFN.scala 220:77]
  wire  _common_underflow_T_13; // @[RoundAnyRawFNToRecFN.scala 224:38]
  wire  _common_underflow_T_14; // @[RoundAnyRawFNToRecFN.scala 225:45]
  wire  _common_underflow_T_15; // @[RoundAnyRawFNToRecFN.scala 225:60]
  wire  _common_underflow_T_17; // @[RoundAnyRawFNToRecFN.scala 219:76]
  wire  common_underflow; // @[RoundAnyRawFNToRecFN.scala 215:40]
  wire  common_inexact; // @[RoundAnyRawFNToRecFN.scala 228:49]
  wire  isNaNOut; // @[RoundAnyRawFNToRecFN.scala 233:34]
  wire  notNaN_isSpecialInfOut; // @[RoundAnyRawFNToRecFN.scala 234:49]
  wire  _commonCase_T_2; // @[RoundAnyRawFNToRecFN.scala 235:33]
  wire  commonCase; // @[RoundAnyRawFNToRecFN.scala 235:61]
  wire  overflow; // @[RoundAnyRawFNToRecFN.scala 236:32]
  wire  underflow; // @[RoundAnyRawFNToRecFN.scala 237:32]
  wire  _inexact_T; // @[RoundAnyRawFNToRecFN.scala 238:43]
  wire  inexact; // @[RoundAnyRawFNToRecFN.scala 238:28]
  wire  overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 241:60]
  wire  _pegMinNonzeroMagOut_T; // @[RoundAnyRawFNToRecFN.scala 243:20]
  wire  _pegMinNonzeroMagOut_T_1; // @[RoundAnyRawFNToRecFN.scala 243:60]
  wire  pegMinNonzeroMagOut; // @[RoundAnyRawFNToRecFN.scala 243:45]
  wire  pegMaxFiniteMagOut; // @[RoundAnyRawFNToRecFN.scala 244:39]
  wire  _notNaN_isInfOut_T; // @[RoundAnyRawFNToRecFN.scala 246:45]
  wire  notNaN_isInfOut; // @[RoundAnyRawFNToRecFN.scala 246:32]
  wire  signOut; // @[RoundAnyRawFNToRecFN.scala 248:22]
  wire  _expOut_T; // @[RoundAnyRawFNToRecFN.scala 251:32]
  wire [11:0] _expOut_T_1; // @[RoundAnyRawFNToRecFN.scala 251:18]
  wire [11:0] _expOut_T_3; // @[RoundAnyRawFNToRecFN.scala 250:24]
  wire [11:0] _expOut_T_5; // @[RoundAnyRawFNToRecFN.scala 255:18]
  wire [11:0] _expOut_T_7; // @[RoundAnyRawFNToRecFN.scala 254:17]
  wire [11:0] _expOut_T_8; // @[RoundAnyRawFNToRecFN.scala 259:18]
  wire [11:0] _expOut_T_10; // @[RoundAnyRawFNToRecFN.scala 258:17]
  wire [11:0] _expOut_T_11; // @[RoundAnyRawFNToRecFN.scala 263:18]
  wire [11:0] _expOut_T_13; // @[RoundAnyRawFNToRecFN.scala 262:17]
  wire [11:0] _expOut_T_14; // @[RoundAnyRawFNToRecFN.scala 267:16]
  wire [11:0] _expOut_T_15; // @[RoundAnyRawFNToRecFN.scala 266:18]
  wire [11:0] _expOut_T_16; // @[RoundAnyRawFNToRecFN.scala 271:16]
  wire [11:0] _expOut_T_17; // @[RoundAnyRawFNToRecFN.scala 270:15]
  wire [11:0] _expOut_T_18; // @[RoundAnyRawFNToRecFN.scala 275:16]
  wire [11:0] _expOut_T_19; // @[RoundAnyRawFNToRecFN.scala 274:15]
  wire [11:0] _expOut_T_20; // @[RoundAnyRawFNToRecFN.scala 276:16]
  wire [11:0] expOut; // @[RoundAnyRawFNToRecFN.scala 275:77]
  wire  _fractOut_T; // @[RoundAnyRawFNToRecFN.scala 278:22]
  wire  _fractOut_T_1; // @[RoundAnyRawFNToRecFN.scala 278:38]
  wire [51:0] _fractOut_T_2; // @[RoundAnyRawFNToRecFN.scala 279:16]
  wire [51:0] _fractOut_T_3; // @[RoundAnyRawFNToRecFN.scala 278:12]
  wire [51:0] _fractOut_T_5; // @[Bitwise.scala 72:12]
  wire [51:0] fractOut; // @[RoundAnyRawFNToRecFN.scala 281:11]
  wire [12:0] io_out_hi; // @[Cat.scala 30:58]
  wire [1:0] io_exceptionFlags_lo; // @[Cat.scala 30:58]
  wire [2:0] io_exceptionFlags_hi; // @[Cat.scala 30:58]
  wire [29:0] RoundAnyRawFNToRecFN_6_covSum;
  assign roundingMode_near_even = io_roundingMode == 3'h0; // @[RoundAnyRawFNToRecFN.scala 88:53]
  assign roundingMode_min = io_roundingMode == 3'h2; // @[RoundAnyRawFNToRecFN.scala 90:53]
  assign roundingMode_max = io_roundingMode == 3'h3; // @[RoundAnyRawFNToRecFN.scala 91:53]
  assign roundingMode_near_maxMag = io_roundingMode == 3'h4; // @[RoundAnyRawFNToRecFN.scala 92:53]
  assign roundingMode_odd = io_roundingMode == 3'h6; // @[RoundAnyRawFNToRecFN.scala 93:53]
  assign _roundMagUp_T = roundingMode_min & io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:27]
  assign _roundMagUp_T_2 = roundingMode_max & ~io_in_sign; // @[RoundAnyRawFNToRecFN.scala 96:63]
  assign roundMagUp = _roundMagUp_T | _roundMagUp_T_2; // @[RoundAnyRawFNToRecFN.scala 96:42]
  assign doShiftSigDown1 = io_in_sig[55]; // @[RoundAnyRawFNToRecFN.scala 118:61]
  assign roundMask_msb = ~io_in_sExp[11]; // @[primitives.scala 57:25]
  assign roundMask_lsbs = ~io_in_sExp[10:0]; // @[primitives.scala 58:26]
  assign roundMask_msb_1 = roundMask_lsbs[10]; // @[primitives.scala 57:25]
  assign roundMask_lsbs_1 = roundMask_lsbs[9:0]; // @[primitives.scala 58:26]
  assign roundMask_msb_2 = roundMask_lsbs_1[9]; // @[primitives.scala 57:25]
  assign roundMask_lsbs_2 = roundMask_lsbs_1[8:0]; // @[primitives.scala 58:26]
  assign roundMask_msb_3 = roundMask_lsbs_2[8]; // @[primitives.scala 57:25]
  assign roundMask_lsbs_3 = roundMask_lsbs_2[7:0]; // @[primitives.scala 58:26]
  assign roundMask_msb_4 = roundMask_lsbs_3[7]; // @[primitives.scala 57:25]
  assign roundMask_lsbs_4 = roundMask_lsbs_3[6:0]; // @[primitives.scala 58:26]
  assign roundMask_msb_5 = roundMask_lsbs_4[6]; // @[primitives.scala 57:25]
  assign roundMask_lsbs_5 = roundMask_lsbs_4[5:0]; // @[primitives.scala 58:26]
  assign roundMask_shift = -65'sh10000000000000000 >>> roundMask_lsbs_5; // @[primitives.scala 77:58]
  assign _roundMask_T_7 = {{16'd0}, roundMask_shift[44:29]}; // @[Bitwise.scala 103:31]
  assign _roundMask_T_9 = {roundMask_shift[28:13], 16'h0}; // @[Bitwise.scala 103:65]
  assign _roundMask_T_11 = _roundMask_T_9 & 32'hffff0000; // @[Bitwise.scala 103:75]
  assign _roundMask_T_12 = _roundMask_T_7 | _roundMask_T_11; // @[Bitwise.scala 103:39]
  assign _GEN_0 = {{8'd0}, _roundMask_T_12[31:8]}; // @[Bitwise.scala 103:31]
  assign _roundMask_T_17 = _GEN_0 & 32'hff00ff; // @[Bitwise.scala 103:31]
  assign _roundMask_T_19 = {_roundMask_T_12[23:0], 8'h0}; // @[Bitwise.scala 103:65]
  assign _roundMask_T_21 = _roundMask_T_19 & 32'hff00ff00; // @[Bitwise.scala 103:75]
  assign _roundMask_T_22 = _roundMask_T_17 | _roundMask_T_21; // @[Bitwise.scala 103:39]
  assign _GEN_1 = {{4'd0}, _roundMask_T_22[31:4]}; // @[Bitwise.scala 103:31]
  assign _roundMask_T_27 = _GEN_1 & 32'hf0f0f0f; // @[Bitwise.scala 103:31]
  assign _roundMask_T_29 = {_roundMask_T_22[27:0], 4'h0}; // @[Bitwise.scala 103:65]
  assign _roundMask_T_31 = _roundMask_T_29 & 32'hf0f0f0f0; // @[Bitwise.scala 103:75]
  assign _roundMask_T_32 = _roundMask_T_27 | _roundMask_T_31; // @[Bitwise.scala 103:39]
  assign _GEN_2 = {{2'd0}, _roundMask_T_32[31:2]}; // @[Bitwise.scala 103:31]
  assign _roundMask_T_37 = _GEN_2 & 32'h33333333; // @[Bitwise.scala 103:31]
  assign _roundMask_T_39 = {_roundMask_T_32[29:0], 2'h0}; // @[Bitwise.scala 103:65]
  assign _roundMask_T_41 = _roundMask_T_39 & 32'hcccccccc; // @[Bitwise.scala 103:75]
  assign _roundMask_T_42 = _roundMask_T_37 | _roundMask_T_41; // @[Bitwise.scala 103:39]
  assign _GEN_3 = {{1'd0}, _roundMask_T_42[31:1]}; // @[Bitwise.scala 103:31]
  assign _roundMask_T_47 = _GEN_3 & 32'h55555555; // @[Bitwise.scala 103:31]
  assign _roundMask_T_49 = {_roundMask_T_42[30:0], 1'h0}; // @[Bitwise.scala 103:65]
  assign _roundMask_T_51 = _roundMask_T_49 & 32'haaaaaaaa; // @[Bitwise.scala 103:75]
  assign roundMask_hi = _roundMask_T_47 | _roundMask_T_51; // @[Bitwise.scala 103:39]
  assign _roundMask_T_57 = {{8'd0}, roundMask_shift[60:53]}; // @[Bitwise.scala 103:31]
  assign _roundMask_T_59 = {roundMask_shift[52:45], 8'h0}; // @[Bitwise.scala 103:65]
  assign _roundMask_T_61 = _roundMask_T_59 & 16'hff00; // @[Bitwise.scala 103:75]
  assign _roundMask_T_62 = _roundMask_T_57 | _roundMask_T_61; // @[Bitwise.scala 103:39]
  assign _GEN_4 = {{4'd0}, _roundMask_T_62[15:4]}; // @[Bitwise.scala 103:31]
  assign _roundMask_T_67 = _GEN_4 & 16'hf0f; // @[Bitwise.scala 103:31]
  assign _roundMask_T_69 = {_roundMask_T_62[11:0], 4'h0}; // @[Bitwise.scala 103:65]
  assign _roundMask_T_71 = _roundMask_T_69 & 16'hf0f0; // @[Bitwise.scala 103:75]
  assign _roundMask_T_72 = _roundMask_T_67 | _roundMask_T_71; // @[Bitwise.scala 103:39]
  assign _GEN_5 = {{2'd0}, _roundMask_T_72[15:2]}; // @[Bitwise.scala 103:31]
  assign _roundMask_T_77 = _GEN_5 & 16'h3333; // @[Bitwise.scala 103:31]
  assign _roundMask_T_79 = {_roundMask_T_72[13:0], 2'h0}; // @[Bitwise.scala 103:65]
  assign _roundMask_T_81 = _roundMask_T_79 & 16'hcccc; // @[Bitwise.scala 103:75]
  assign _roundMask_T_82 = _roundMask_T_77 | _roundMask_T_81; // @[Bitwise.scala 103:39]
  assign _GEN_6 = {{1'd0}, _roundMask_T_82[15:1]}; // @[Bitwise.scala 103:31]
  assign _roundMask_T_87 = _GEN_6 & 16'h5555; // @[Bitwise.scala 103:31]
  assign _roundMask_T_89 = {_roundMask_T_82[14:0], 1'h0}; // @[Bitwise.scala 103:65]
  assign _roundMask_T_91 = _roundMask_T_89 & 16'haaaa; // @[Bitwise.scala 103:75]
  assign roundMask_hi_1 = _roundMask_T_87 | _roundMask_T_91; // @[Bitwise.scala 103:39]
  assign roundMask_hi_2 = roundMask_shift[61]; // @[Bitwise.scala 109:18]
  assign roundMask_lo = roundMask_shift[62]; // @[Bitwise.scala 109:44]
  assign roundMask_lo_1 = roundMask_shift[63]; // @[Bitwise.scala 109:44]
  assign _roundMask_T_94 = {roundMask_hi,roundMask_hi_1,roundMask_hi_2,roundMask_lo,roundMask_lo_1}; // @[Cat.scala 30:58]
  assign _roundMask_T_96 = roundMask_msb_5 ? 51'h0 : ~_roundMask_T_94; // @[primitives.scala 74:21]
  assign _roundMask_T_99 = roundMask_msb_4 ? 51'h0 : _roundMask_T_96[50:0]; // @[primitives.scala 74:21]
  assign _roundMask_T_102 = roundMask_msb_3 ? 51'h0 : _roundMask_T_99[50:0]; // @[primitives.scala 74:21]
  assign _roundMask_T_105 = roundMask_msb_2 ? 51'h0 : _roundMask_T_102[50:0]; // @[primitives.scala 74:21]
  assign roundMask_hi_4 = ~_roundMask_T_105; // @[primitives.scala 74:17]
  assign _roundMask_T_106 = {roundMask_hi_4,3'h7}; // @[Cat.scala 30:58]
  assign roundMask_hi_5 = roundMask_shift[0]; // @[Bitwise.scala 109:18]
  assign roundMask_lo_4 = roundMask_shift[1]; // @[Bitwise.scala 109:44]
  assign roundMask_lo_5 = roundMask_shift[2]; // @[Bitwise.scala 109:44]
  assign _roundMask_T_109 = {roundMask_hi_5,roundMask_lo_4,roundMask_lo_5}; // @[Cat.scala 30:58]
  assign _roundMask_T_110 = roundMask_msb_5 ? _roundMask_T_109 : 3'h0; // @[primitives.scala 61:24]
  assign _roundMask_T_111 = roundMask_msb_4 ? _roundMask_T_110 : 3'h0; // @[primitives.scala 61:24]
  assign _roundMask_T_112 = roundMask_msb_3 ? _roundMask_T_111 : 3'h0; // @[primitives.scala 61:24]
  assign _roundMask_T_113 = roundMask_msb_2 ? _roundMask_T_112 : 3'h0; // @[primitives.scala 61:24]
  assign _roundMask_T_114 = roundMask_msb_1 ? _roundMask_T_106 : {{51'd0}, _roundMask_T_113}; // @[primitives.scala 66:24]
  assign _roundMask_T_115 = roundMask_msb ? _roundMask_T_114 : 54'h0; // @[primitives.scala 61:24]
  assign _GEN_7 = {{53'd0}, doShiftSigDown1}; // @[RoundAnyRawFNToRecFN.scala 157:23]
  assign roundMask_hi_7 = _roundMask_T_115 | _GEN_7; // @[RoundAnyRawFNToRecFN.scala 157:23]
  assign roundMask = {roundMask_hi_7,2'h3}; // @[Cat.scala 30:58]
  assign shiftedRoundMask_lo = roundMask[55:1]; // @[RoundAnyRawFNToRecFN.scala 160:57]
  assign shiftedRoundMask = {1'h0,shiftedRoundMask_lo}; // @[Cat.scala 30:58]
  assign roundPosMask = ~shiftedRoundMask & roundMask; // @[RoundAnyRawFNToRecFN.scala 161:46]
  assign _roundPosBit_T = io_in_sig & roundPosMask; // @[RoundAnyRawFNToRecFN.scala 162:40]
  assign roundPosBit = |_roundPosBit_T; // @[RoundAnyRawFNToRecFN.scala 162:56]
  assign _anyRoundExtra_T = io_in_sig & shiftedRoundMask; // @[RoundAnyRawFNToRecFN.scala 163:42]
  assign anyRoundExtra = |_anyRoundExtra_T; // @[RoundAnyRawFNToRecFN.scala 163:62]
  assign anyRound = roundPosBit | anyRoundExtra; // @[RoundAnyRawFNToRecFN.scala 164:36]
  assign _roundIncr_T = roundingMode_near_even | roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 167:38]
  assign _roundIncr_T_1 = _roundIncr_T & roundPosBit; // @[RoundAnyRawFNToRecFN.scala 167:67]
  assign _roundIncr_T_2 = roundMagUp & anyRound; // @[RoundAnyRawFNToRecFN.scala 169:29]
  assign roundIncr = _roundIncr_T_1 | _roundIncr_T_2; // @[RoundAnyRawFNToRecFN.scala 168:31]
  assign _roundedSig_T = io_in_sig | roundMask; // @[RoundAnyRawFNToRecFN.scala 172:32]
  assign _roundedSig_T_2 = _roundedSig_T[55:2] + 54'h1; // @[RoundAnyRawFNToRecFN.scala 172:49]
  assign _roundedSig_T_3 = roundingMode_near_even & roundPosBit; // @[RoundAnyRawFNToRecFN.scala 173:49]
  assign _roundedSig_T_5 = _roundedSig_T_3 & ~anyRoundExtra; // @[RoundAnyRawFNToRecFN.scala 173:64]
  assign _roundedSig_T_7 = _roundedSig_T_5 ? shiftedRoundMask_lo : 55'h0; // @[RoundAnyRawFNToRecFN.scala 173:25]
  assign _roundedSig_T_9 = _roundedSig_T_2 & ~_roundedSig_T_7; // @[RoundAnyRawFNToRecFN.scala 172:61]
  assign _roundedSig_T_11 = io_in_sig & ~roundMask; // @[RoundAnyRawFNToRecFN.scala 178:30]
  assign _roundedSig_T_13 = roundingMode_odd & anyRound; // @[RoundAnyRawFNToRecFN.scala 179:42]
  assign _roundedSig_T_15 = _roundedSig_T_13 ? roundPosMask[55:1] : 55'h0; // @[RoundAnyRawFNToRecFN.scala 179:24]
  assign _GEN_8 = {{1'd0}, _roundedSig_T_11[55:2]}; // @[RoundAnyRawFNToRecFN.scala 178:47]
  assign _roundedSig_T_16 = _GEN_8 | _roundedSig_T_15; // @[RoundAnyRawFNToRecFN.scala 178:47]
  assign roundedSig = roundIncr ? _roundedSig_T_9 : _roundedSig_T_16; // @[RoundAnyRawFNToRecFN.scala 171:16]
  assign _sRoundedExp_T_1 = {1'b0,$signed(roundedSig[54:53])}; // @[RoundAnyRawFNToRecFN.scala 183:69]
  assign _GEN_9 = {{10{_sRoundedExp_T_1[2]}},_sRoundedExp_T_1}; // @[RoundAnyRawFNToRecFN.scala 183:40]
  assign sRoundedExp = $signed(io_in_sExp) + $signed(_GEN_9); // @[RoundAnyRawFNToRecFN.scala 183:40]
  assign common_expOut = sRoundedExp[11:0]; // @[RoundAnyRawFNToRecFN.scala 185:37]
  assign common_fractOut = doShiftSigDown1 ? roundedSig[52:1] : roundedSig[51:0]; // @[RoundAnyRawFNToRecFN.scala 187:16]
  assign _common_overflow_T = sRoundedExp[13:10]; // @[RoundAnyRawFNToRecFN.scala 194:30]
  assign common_overflow = $signed(_common_overflow_T) >= 4'sh3; // @[RoundAnyRawFNToRecFN.scala 194:50]
  assign common_totalUnderflow = $signed(sRoundedExp) < 14'sh3ce; // @[RoundAnyRawFNToRecFN.scala 198:31]
  assign unboundedRange_roundPosBit = doShiftSigDown1 ? io_in_sig[2] : io_in_sig[1]; // @[RoundAnyRawFNToRecFN.scala 201:16]
  assign _unboundedRange_anyRound_T_1 = doShiftSigDown1 & io_in_sig[2]; // @[RoundAnyRawFNToRecFN.scala 203:30]
  assign _unboundedRange_anyRound_T_3 = |io_in_sig[1:0]; // @[RoundAnyRawFNToRecFN.scala 203:70]
  assign unboundedRange_anyRound = _unboundedRange_anyRound_T_1 | _unboundedRange_anyRound_T_3; // @[RoundAnyRawFNToRecFN.scala 203:49]
  assign _unboundedRange_roundIncr_T_1 = _roundIncr_T & unboundedRange_roundPosBit; // @[RoundAnyRawFNToRecFN.scala 205:67]
  assign _unboundedRange_roundIncr_T_2 = roundMagUp & unboundedRange_anyRound; // @[RoundAnyRawFNToRecFN.scala 207:29]
  assign unboundedRange_roundIncr = _unboundedRange_roundIncr_T_1 | _unboundedRange_roundIncr_T_2; // @[RoundAnyRawFNToRecFN.scala 206:46]
  assign roundCarry = doShiftSigDown1 ? roundedSig[54] : roundedSig[53]; // @[RoundAnyRawFNToRecFN.scala 209:16]
  assign _common_underflow_T = io_in_sExp[12:11]; // @[RoundAnyRawFNToRecFN.scala 218:48]
  assign _common_underflow_T_1 = $signed(_common_underflow_T) <= 2'sh0; // @[RoundAnyRawFNToRecFN.scala 218:62]
  assign _common_underflow_T_2 = anyRound & _common_underflow_T_1; // @[RoundAnyRawFNToRecFN.scala 218:32]
  assign _common_underflow_T_5 = doShiftSigDown1 ? roundMask[3] : roundMask[2]; // @[RoundAnyRawFNToRecFN.scala 219:30]
  assign _common_underflow_T_6 = _common_underflow_T_2 & _common_underflow_T_5; // @[RoundAnyRawFNToRecFN.scala 218:74]
  assign _common_underflow_T_10 = doShiftSigDown1 ? roundMask[4] : roundMask[3]; // @[RoundAnyRawFNToRecFN.scala 221:39]
  assign _common_underflow_T_12 = io_detectTininess & ~_common_underflow_T_10; // @[RoundAnyRawFNToRecFN.scala 220:77]
  assign _common_underflow_T_13 = _common_underflow_T_12 & roundCarry; // @[RoundAnyRawFNToRecFN.scala 224:38]
  assign _common_underflow_T_14 = _common_underflow_T_13 & roundPosBit; // @[RoundAnyRawFNToRecFN.scala 225:45]
  assign _common_underflow_T_15 = _common_underflow_T_14 & unboundedRange_roundIncr; // @[RoundAnyRawFNToRecFN.scala 225:60]
  assign _common_underflow_T_17 = _common_underflow_T_6 & ~_common_underflow_T_15; // @[RoundAnyRawFNToRecFN.scala 219:76]
  assign common_underflow = common_totalUnderflow | _common_underflow_T_17; // @[RoundAnyRawFNToRecFN.scala 215:40]
  assign common_inexact = common_totalUnderflow | anyRound; // @[RoundAnyRawFNToRecFN.scala 228:49]
  assign isNaNOut = io_invalidExc | io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 233:34]
  assign notNaN_isSpecialInfOut = io_infiniteExc | io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 234:49]
  assign _commonCase_T_2 = ~isNaNOut & ~notNaN_isSpecialInfOut; // @[RoundAnyRawFNToRecFN.scala 235:33]
  assign commonCase = _commonCase_T_2 & ~io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 235:61]
  assign overflow = commonCase & common_overflow; // @[RoundAnyRawFNToRecFN.scala 236:32]
  assign underflow = commonCase & common_underflow; // @[RoundAnyRawFNToRecFN.scala 237:32]
  assign _inexact_T = commonCase & common_inexact; // @[RoundAnyRawFNToRecFN.scala 238:43]
  assign inexact = overflow | _inexact_T; // @[RoundAnyRawFNToRecFN.scala 238:28]
  assign overflow_roundMagUp = _roundIncr_T | roundMagUp; // @[RoundAnyRawFNToRecFN.scala 241:60]
  assign _pegMinNonzeroMagOut_T = commonCase & common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 243:20]
  assign _pegMinNonzeroMagOut_T_1 = roundMagUp | roundingMode_odd; // @[RoundAnyRawFNToRecFN.scala 243:60]
  assign pegMinNonzeroMagOut = _pegMinNonzeroMagOut_T & _pegMinNonzeroMagOut_T_1; // @[RoundAnyRawFNToRecFN.scala 243:45]
  assign pegMaxFiniteMagOut = overflow & ~overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 244:39]
  assign _notNaN_isInfOut_T = overflow & overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 246:45]
  assign notNaN_isInfOut = notNaN_isSpecialInfOut | _notNaN_isInfOut_T; // @[RoundAnyRawFNToRecFN.scala 246:32]
  assign signOut = isNaNOut ? 1'h0 : io_in_sign; // @[RoundAnyRawFNToRecFN.scala 248:22]
  assign _expOut_T = io_in_isZero | common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 251:32]
  assign _expOut_T_1 = _expOut_T ? 12'he00 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 251:18]
  assign _expOut_T_3 = common_expOut & ~_expOut_T_1; // @[RoundAnyRawFNToRecFN.scala 250:24]
  assign _expOut_T_5 = pegMinNonzeroMagOut ? 12'hc31 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 255:18]
  assign _expOut_T_7 = _expOut_T_3 & ~_expOut_T_5; // @[RoundAnyRawFNToRecFN.scala 254:17]
  assign _expOut_T_8 = pegMaxFiniteMagOut ? 12'h400 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 259:18]
  assign _expOut_T_10 = _expOut_T_7 & ~_expOut_T_8; // @[RoundAnyRawFNToRecFN.scala 258:17]
  assign _expOut_T_11 = notNaN_isInfOut ? 12'h200 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 263:18]
  assign _expOut_T_13 = _expOut_T_10 & ~_expOut_T_11; // @[RoundAnyRawFNToRecFN.scala 262:17]
  assign _expOut_T_14 = pegMinNonzeroMagOut ? 12'h3ce : 12'h0; // @[RoundAnyRawFNToRecFN.scala 267:16]
  assign _expOut_T_15 = _expOut_T_13 | _expOut_T_14; // @[RoundAnyRawFNToRecFN.scala 266:18]
  assign _expOut_T_16 = pegMaxFiniteMagOut ? 12'hbff : 12'h0; // @[RoundAnyRawFNToRecFN.scala 271:16]
  assign _expOut_T_17 = _expOut_T_15 | _expOut_T_16; // @[RoundAnyRawFNToRecFN.scala 270:15]
  assign _expOut_T_18 = notNaN_isInfOut ? 12'hc00 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 275:16]
  assign _expOut_T_19 = _expOut_T_17 | _expOut_T_18; // @[RoundAnyRawFNToRecFN.scala 274:15]
  assign _expOut_T_20 = isNaNOut ? 12'he00 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 276:16]
  assign expOut = _expOut_T_19 | _expOut_T_20; // @[RoundAnyRawFNToRecFN.scala 275:77]
  assign _fractOut_T = isNaNOut | io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 278:22]
  assign _fractOut_T_1 = _fractOut_T | common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 278:38]
  assign _fractOut_T_2 = isNaNOut ? 52'h8000000000000 : 52'h0; // @[RoundAnyRawFNToRecFN.scala 279:16]
  assign _fractOut_T_3 = _fractOut_T_1 ? _fractOut_T_2 : common_fractOut; // @[RoundAnyRawFNToRecFN.scala 278:12]
  assign _fractOut_T_5 = pegMaxFiniteMagOut ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 72:12]
  assign fractOut = _fractOut_T_3 | _fractOut_T_5; // @[RoundAnyRawFNToRecFN.scala 281:11]
  assign io_out_hi = {signOut,expOut}; // @[Cat.scala 30:58]
  assign io_exceptionFlags_lo = {underflow,inexact}; // @[Cat.scala 30:58]
  assign io_exceptionFlags_hi = {io_invalidExc,io_infiniteExc,overflow}; // @[Cat.scala 30:58]
  assign io_out = {io_out_hi,fractOut}; // @[RoundAnyRawFNToRecFN.scala 284:12]
  assign io_exceptionFlags = {io_exceptionFlags_hi,io_exceptionFlags_lo}; // @[RoundAnyRawFNToRecFN.scala 285:23]
  assign RoundAnyRawFNToRecFN_6_covSum = 30'h0;
  assign io_covSum = RoundAnyRawFNToRecFN_6_covSum;
  assign metaAssert = 1'h0;
endmodule
